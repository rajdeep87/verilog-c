module m6s18 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74;

output p0;

wire na832,na850,na862,na880,na902,na844,na896,a874,na1318,na1334,na1342,na1336,na1354,na1328,na1348,
na1366,na1384,na1402,na1430,na1448,na1466,na1484,na1502,na1520,na1538,na1556,na1574,na1586,na1598,na1622,
na1674,na1708,na1730,na1742,na1760,na1778,na1796,na1814,na1832,na1848,na1880,na1916,na1954,na1970,na1982,
na2000,na2044,na2056,na2074,na2092,na2108,na2126,na2138,na2160,na2176,na2188,na2204,na2216,na2232,na2250,
na1312,na2244,na2226,na2210,na2264,na2198,na2258,na2182,na2278,na2170,na2292,na2306,na2272,na2300,na2286,
na2154,na2132,na2120,na2102,na2324,na2346,na2086,na2340,na2364,na2318,na2358,na2068,na2050,na2388,na2400,
na2412,na2424,na2436,na2448,na2466,na2482,na2038,na2476,na2460,na2494,na2442,na2506,na2488,na2518,na2500,
na2530,na2512,na2542,na2524,na2554,na2536,na2570,na2548,na2582,na2564,na2594,na2576,na2606,na2588,na2618,
na2600,na2612,na2430,na2418,na2406,na2394,na2382,na1994,na1976,na2636,na1964,na2658,na2630,na2652,na2708,
na2738,na2764,na2784,na1948,na2778,na2796,na2758,na2790,na2732,na2702,na1910,na1874,na1842,na1826,na1808,
na1790,na1772,na1754,na1736,na2830,na2860,na2886,na2912,na2942,na2964,na2986,na3004,na3026,na1724,na3020,
na2998,na2980,na2958,na2936,na2906,na2880,na2854,na2824,na1702,na1668,na1616,na1592,na1580,na1568,na1550,
na1532,na1514,na1496,na1478,na1460,na1442,na1424,na1396,na1378,na1360,na856,na3044,na3062,na826,na3056,
a3038,na3450,na3466,na3470,na3460,na3482,na3500,na3518,na3536,na3554,na3572,na3590,na3608,na3626,na3644,
na3662,na3680,na3692,na3742,na3754,na3778,na3818,na3836,na3848,na3866,na3884,na3902,na3920,na3938,na3954,
na3992,na4026,na4050,na4066,na4072,na4090,na4130,na4142,na4160,na4176,na4194,na4206,na4228,na4244,na4250,
na4266,na4272,na4288,na4306,na3444,na4300,na4282,na4320,na4260,na4314,na4334,na4238,na4348,na4362,na4328,
na4356,na4342,na4222,na4200,na4188,na4170,na4380,na4402,na4154,na4396,na4420,na4374,na4414,na4136,na4426,
na4442,na4448,na4454,na4460,na4472,na4492,na4510,na4124,na4504,na4486,na4522,na4466,na4534,na4516,na4546,
na4528,na4558,na4540,na4570,na4552,na4582,na4564,na4594,na4576,na4606,na4588,na4618,na4600,na4630,na4612,
na4642,na4624,na4636,na4436,na4084,na4660,na4060,na4682,na4654,na4676,na4720,na4752,na4772,na4798,na4044,
na4792,na4766,na4746,na4804,na4714,na4020,na3986,na3948,na3932,na3914,na3896,na3878,na3860,na3842,na4838,
na4868,na4894,na4920,na4950,na4972,na4994,na5012,na5034,na3830,na5028,na5006,na4988,na4966,na4944,na4914,
na4888,na4862,na4832,na3812,na3772,na3748,na3736,na3686,na3674,na3656,na3638,na3620,na3602,na3584,na3566,
na3548,na3530,na3512,na3494,na3476,c1,a810,a812,a814,a816,a818,a820,a822,a824,a826,
a828,a830,a832,a834,a836,a838,a840,a842,a844,a846,a848,a850,a852,a854,a856,
a858,a860,a862,a864,a866,a868,a870,a872,a876,a878,a880,a882,a884,a886,a888,
a890,a892,a894,a896,a898,a900,a902,a904,a906,a908,a910,a912,a914,a916,a918,
a920,a922,a924,a926,a928,a930,a932,a934,a936,a938,a940,a942,a944,a946,a948,
a950,a952,a954,a956,a958,a960,a962,a964,a966,a968,a970,a972,a974,a976,a978,
a980,a982,a984,a986,a988,a990,a992,a994,a996,a998,a1000,a1002,a1004,a1006,a1008,
a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,a1038,
a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,a1062,a1064,a1066,a1068,
a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,a1092,a1094,a1096,a1098,
a1100,a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,a1124,a1126,a1128,
a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,a1154,a1156,a1158,
a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,a1178,a1180,a1182,a1184,a1186,a1188,
a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,a1218,
a1220,a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,a1248,
a1250,a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,a1268,a1270,a1272,a1274,a1276,a1278,
a1280,a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,
a1310,a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,a1334,a1336,a1338,
a1340,a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,a1368,
a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,a1388,a1390,a1392,a1394,a1396,a1398,
a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1426,a1428,
a1430,a1432,a1434,a1436,a1438,a1440,a1442,a1444,a1446,a1448,a1450,a1452,a1454,a1456,a1458,
a1460,a1462,a1464,a1466,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1482,a1484,a1486,a1488,
a1490,a1492,a1494,a1496,a1498,a1500,a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,a1518,
a1520,a1522,a1524,a1526,a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,a1548,
a1550,a1552,a1554,a1556,a1558,a1560,a1562,a1564,a1566,a1568,a1570,a1572,a1574,a1576,a1578,
a1580,a1582,a1584,a1586,a1588,a1590,a1592,a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,
a1610,a1612,a1614,a1616,a1618,a1620,a1622,a1624,a1626,a1628,a1630,a1632,a1634,a1636,a1638,
a1640,a1642,a1644,a1646,a1648,a1650,a1652,a1654,a1656,a1658,a1660,a1662,a1664,a1666,a1668,
a1670,a1672,a1674,a1676,a1678,a1680,a1682,a1684,a1686,a1688,a1690,a1692,a1694,a1696,a1698,
a1700,a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,
a1730,a1732,a1734,a1736,a1738,a1740,a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,a1758,
a1760,a1762,a1764,a1766,a1768,a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,
a1790,a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,
a1820,a1822,a1824,a1826,a1828,a1830,a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,a1848,
a1850,a1852,a1854,a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,
a1880,a1882,a1884,a1886,a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,
a1910,a1912,a1914,a1916,a1918,a1920,a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,a1938,
a1940,a1942,a1944,a1946,a1948,a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,
a1970,a1972,a1974,a1976,a1978,a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,a1998,
a2000,a2002,a2004,a2006,a2008,a2010,a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,
a2030,a2032,a2034,a2036,a2038,a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,a2058,
a2060,a2062,a2064,a2066,a2068,a2070,a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,
a2090,a2092,a2094,a2096,a2098,a2100,a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,
a2120,a2122,a2124,a2126,a2128,a2130,a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,
a2150,a2152,a2154,a2156,a2158,a2160,a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,a2178,
a2180,a2182,a2184,a2186,a2188,a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,a2208,
a2210,a2212,a2214,a2216,a2218,a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,a2238,
a2240,a2242,a2244,a2246,a2248,a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,a2268,
a2270,a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,a2298,
a2300,a2302,a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,a2328,
a2330,a2332,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,a2358,
a2360,a2362,a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,a2388,
a2390,a2392,a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,
a2420,a2422,a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,a2448,
a2450,a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,a2478,
a2480,a2482,a2484,a2486,a2488,a2490,a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,a2508,
a2510,a2512,a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,
a2540,a2542,a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,
a2570,a2572,a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,
a2600,a2602,a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,
a2630,a2632,a2634,a2636,a2638,a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,
a2660,a2662,a2664,a2666,a2668,a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,
a2690,a2692,a2694,a2696,a2698,a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,a2718,
a2720,a2722,a2724,a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,
a2750,a2752,a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,
a2780,a2782,a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,
a2810,a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,
a2840,a2842,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,
a2870,a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,
a2900,a2902,a2904,a2906,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,
a2930,a2932,a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,
a2960,a2962,a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,a2988,
a2990,a2992,a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,
a3020,a3022,a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3040,a3042,a3044,a3046,a3048,a3050,
a3052,a3054,a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,a3078,a3080,
a3082,a3084,a3086,a3088,a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,
a3112,a3114,a3116,a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,
a3142,a3144,a3146,a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,
a3172,a3174,a3176,a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3200,
a3202,a3204,a3206,a3208,a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,a3228,a3230,
a3232,a3234,a3236,a3238,a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,
a3262,a3264,a3266,a3268,a3270,a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,a3288,a3290,
a3292,a3294,a3296,a3298,a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,
a3322,a3324,a3326,a3328,a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,
a3352,a3354,a3356,a3358,a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,
a3382,a3384,a3386,a3388,a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,a3408,a3410,
a3412,a3414,a3416,a3418,a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,a3438,a3440,
a3442,a3444,a3446,a3448,a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,a3468,a3470,
a3472,a3474,a3476,a3478,a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,a3498,a3500,
a3502,a3504,a3506,a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,a3528,a3530,
a3532,a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,a3558,a3560,
a3562,a3564,a3566,a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,a3588,a3590,
a3592,a3594,a3596,a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,a3618,a3620,
a3622,a3624,a3626,a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3648,a3650,
a3652,a3654,a3656,a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,a3678,a3680,
a3682,a3684,a3686,a3688,a3690,a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,
a3712,a3714,a3716,a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,a3738,a3740,
a3742,a3744,a3746,a3748,a3750,a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,a3768,a3770,
a3772,a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,a3798,a3800,
a3802,a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,a3828,a3830,
a3832,a3834,a3836,a3838,a3840,a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,a3858,a3860,
a3862,a3864,a3866,a3868,a3870,a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,a3888,a3890,
a3892,a3894,a3896,a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,a3918,a3920,
a3922,a3924,a3926,a3928,a3930,a3932,a3934,a3936,a3938,a3940,a3942,a3944,a3946,a3948,a3950,
a3952,a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,a3978,a3980,
a3982,a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,a4008,a4010,
a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,a4038,a4040,
a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,a4068,a4070,
a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,a4096,a4098,a4100,
a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4124,a4126,a4128,a4130,
a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,a4152,a4154,a4156,a4158,a4160,
a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,a4184,a4186,a4188,a4190,
a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,a4214,a4216,a4218,a4220,
a4222,a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,a4244,a4246,a4248,a4250,
a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,a4274,a4276,a4278,a4280,
a4282,a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,a4306,a4308,a4310,
a4312,a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,a4334,a4336,a4338,a4340,
a4342,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,a4368,a4370,
a4372,a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,a4394,a4396,a4398,a4400,
a4402,a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,
a4432,a4434,a4436,a4438,a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,a4458,a4460,
a4462,a4464,a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4482,a4484,a4486,a4488,a4490,
a4492,a4494,a4496,a4498,a4500,a4502,a4504,a4506,a4508,a4510,a4512,a4514,a4516,a4518,a4520,
a4522,a4524,a4526,a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,
a4552,a4554,a4556,a4558,a4560,a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,a4578,a4580,
a4582,a4584,a4586,a4588,a4590,a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,
a4612,a4614,a4616,a4618,a4620,a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,
a4642,a4644,a4646,a4648,a4650,a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,
a4672,a4674,a4676,a4678,a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,a4696,a4698,a4700,
a4702,a4704,a4706,a4708,a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,a4726,a4728,a4730,
a4732,a4734,a4736,a4738,a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,a4756,a4758,a4760,
a4762,a4764,a4766,a4768,a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4784,a4786,a4788,a4790,
a4792,a4794,a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,a4818,a4820,
a4822,a4824,a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,a4844,a4846,a4848,a4850,
a4852,a4854,a4856,a4858,a4860,a4862,a4864,a4866,a4868,a4870,a4872,a4874,a4876,a4878,a4880,
a4882,a4884,a4886,a4888,a4890,a4892,a4894,a4896,a4898,a4900,a4902,a4904,a4906,a4908,a4910,
a4912,a4914,a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,a4938,a4940,
a4942,a4944,a4946,a4948,a4950,a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,a4968,a4970,
a4972,a4974,a4976,a4978,a4980,a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,a4998,a5000,
a5002,a5004,a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,a5028,a5030,
a5032,a5034,p0;

reg l76,l78,l80,l82,l84,l86,l88,l90,l92,l94,l96,l98,l100,l102,l104,
l106,l108,l110,l112,l114,l116,l118,l120,l122,l124,l126,l128,l130,l132,l134,
l136,l138,l140,l142,l144,l146,l148,l150,l152,l154,l156,l158,l160,l162,l164,
l166,l168,l170,l172,l174,l176,l178,l180,l182,l184,l186,l188,l190,l192,l194,
l196,l198,l200,l202,l204,l206,l208,l210,l212,l214,l216,l218,l220,l222,l224,
l226,l228,l230,l232,l234,l236,l238,l240,l242,l244,l246,l248,l250,l252,l254,
l256,l258,l260,l262,l264,l266,l268,l270,l272,l274,l276,l278,l280,l282,l284,
l286,l288,l290,l292,l294,l296,l298,l300,l302,l304,l306,l308,l310,l312,l314,
l316,l318,l320,l322,l324,l326,l328,l330,l332,l334,l336,l338,l340,l342,l344,
l346,l348,l350,l352,l354,l356,l358,l360,l362,l364,l366,l368,l370,l372,l374,
l376,l378,l380,l382,l384,l386,l388,l390,l392,l394,l396,l398,l400,l402,l404,
l406,l408,l410,l412,l414,l416,l418,l420,l422,l424,l426,l428,l430,l432,l434,
l436,l438,l440,l442,l444,l446,l448,l450,l452,l454,l456,l458,l460,l462,l464,
l466,l468,l470,l472,l474,l476,l478,l480,l482,l484,l486,l488,l490,l492,l494,
l496,l498,l500,l502,l504,l506,l508,l510,l512,l514,l516,l518,l520,l522,l524,
l526,l528,l530,l532,l534,l536,l538,l540,l542,l544,l546,l548,l550,l552,l554,
l556,l558,l560,l562,l564,l566,l568,l570,l572,l574,l576,l578,l580,l582,l584,
l586,l588,l590,l592,l594,l596,l598,l600,l602,l604,l606,l608,l610,l612,l614,
l616,l618,l620,l622,l624,l626,l628,l630,l632,l634,l636,l638,l640,l642,l644,
l646,l648,l650,l652,l654,l656,l658,l660,l662,l664,l666,l668,l670,l672,l674,
l676,l678,l680,l682,l684,l686,l688,l690,l692,l694,l696,l698,l700,l702,l704,
l706,l708,l710,l712,l714,l716,l718,l720,l722,l724,l726,l728,l730,l732,l734,
l736,l738,l740,l742,l744,l746,l748,l750,l752,l754,l756,l758,l760,l762,l764,
l766,l768,l770,l772,l774,l776,l778,l780,l782,l784,l786,l788,l790,l792,l794,
l796,l798,l800,l802,l804,l806,l808;

initial
begin
   l76 = 0;
   l78 = 0;
   l80 = 0;
   l82 = 0;
   l84 = 0;
   l86 = 0;
   l88 = 0;
   l90 = 0;
   l92 = 0;
   l94 = 0;
   l96 = 0;
   l98 = 0;
   l100 = 0;
   l102 = 0;
   l104 = 0;
   l106 = 0;
   l108 = 0;
   l110 = 0;
   l112 = 0;
   l114 = 0;
   l116 = 0;
   l118 = 0;
   l120 = 0;
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
   l392 = 0;
   l394 = 0;
   l396 = 0;
   l398 = 0;
   l400 = 0;
   l402 = 0;
   l404 = 0;
   l406 = 0;
   l408 = 0;
   l410 = 0;
   l412 = 0;
   l414 = 0;
   l416 = 0;
   l418 = 0;
   l420 = 0;
   l422 = 0;
   l424 = 0;
   l426 = 0;
   l428 = 0;
   l430 = 0;
   l432 = 0;
   l434 = 0;
   l436 = 0;
   l438 = 0;
   l440 = 0;
   l442 = 0;
   l444 = 0;
   l446 = 0;
   l448 = 0;
   l450 = 0;
   l452 = 0;
   l454 = 0;
   l456 = 0;
   l458 = 0;
   l460 = 0;
   l462 = 0;
   l464 = 0;
   l466 = 0;
   l468 = 0;
   l470 = 0;
   l472 = 0;
   l474 = 0;
   l476 = 0;
   l478 = 0;
   l480 = 0;
   l482 = 0;
   l484 = 0;
   l486 = 0;
   l488 = 0;
   l490 = 0;
   l492 = 0;
   l494 = 0;
   l496 = 0;
   l498 = 0;
   l500 = 0;
   l502 = 0;
   l504 = 0;
   l506 = 0;
   l508 = 0;
   l510 = 0;
   l512 = 0;
   l514 = 0;
   l516 = 0;
   l518 = 0;
   l520 = 0;
   l522 = 0;
   l524 = 0;
   l526 = 0;
   l528 = 0;
   l530 = 0;
   l532 = 0;
   l534 = 0;
   l536 = 0;
   l538 = 0;
   l540 = 0;
   l542 = 0;
   l544 = 0;
   l546 = 0;
   l548 = 0;
   l550 = 0;
   l552 = 0;
   l554 = 0;
   l556 = 0;
   l558 = 0;
   l560 = 0;
   l562 = 0;
   l564 = 0;
   l566 = 0;
   l568 = 0;
   l570 = 0;
   l572 = 0;
   l574 = 0;
   l576 = 0;
   l578 = 0;
   l580 = 0;
   l582 = 0;
   l584 = 0;
   l586 = 0;
   l588 = 0;
   l590 = 0;
   l592 = 0;
   l594 = 0;
   l596 = 0;
   l598 = 0;
   l600 = 0;
   l602 = 0;
   l604 = 0;
   l606 = 0;
   l608 = 0;
   l610 = 0;
   l612 = 0;
   l614 = 0;
   l616 = 0;
   l618 = 0;
   l620 = 0;
   l622 = 0;
   l624 = 0;
   l626 = 0;
   l628 = 0;
   l630 = 0;
   l632 = 0;
   l634 = 0;
   l636 = 0;
   l638 = 0;
   l640 = 0;
   l642 = 0;
   l644 = 0;
   l646 = 0;
   l648 = 0;
   l650 = 0;
   l652 = 0;
   l654 = 0;
   l656 = 0;
   l658 = 0;
   l660 = 0;
   l662 = 0;
   l664 = 0;
   l666 = 0;
   l668 = 0;
   l670 = 0;
   l672 = 0;
   l674 = 0;
   l676 = 0;
   l678 = 0;
   l680 = 0;
   l682 = 0;
   l684 = 0;
   l686 = 0;
   l688 = 0;
   l690 = 0;
   l692 = 0;
   l694 = 0;
   l696 = 0;
   l698 = 0;
   l700 = 0;
   l702 = 0;
   l704 = 0;
   l706 = 0;
   l708 = 0;
   l710 = 0;
   l712 = 0;
   l714 = 0;
   l716 = 0;
   l718 = 0;
   l720 = 0;
   l722 = 0;
   l724 = 0;
   l726 = 0;
   l728 = 0;
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
   l802 = 0;
   l804 = 0;
   l806 = 0;
   l808 = 0;
end

always @(posedge na832)
   l76 <= na832;

always @(posedge na850)
   l78 <= na850;

always @(posedge i2)
   l80 <= i2;

always @(posedge na862)
   l82 <= na862;

always @(posedge na880)
   l84 <= na880;

always @(posedge na902)
   l86 <= na902;

always @(posedge na844)
   l88 <= na844;

always @(posedge na896)
   l90 <= na896;

always @(posedge a874)
   l92 <= a874;

always @(posedge na1318)
   l94 <= na1318;

always @(posedge na1334)
   l96 <= na1334;

always @(posedge na1342)
   l98 <= na1342;

always @(posedge na1336)
   l100 <= na1336;

always @(posedge na1354)
   l102 <= na1354;

always @(posedge na1328)
   l104 <= na1328;

always @(posedge na1348)
   l106 <= na1348;

always @(posedge na1366)
   l108 <= na1366;

always @(posedge na1384)
   l110 <= na1384;

always @(posedge na1402)
   l112 <= na1402;

always @(posedge na1430)
   l114 <= na1430;

always @(posedge na1448)
   l116 <= na1448;

always @(posedge na1466)
   l118 <= na1466;

always @(posedge na1484)
   l120 <= na1484;

always @(posedge na1502)
   l122 <= na1502;

always @(posedge na1520)
   l124 <= na1520;

always @(posedge na1538)
   l126 <= na1538;

always @(posedge na1556)
   l128 <= na1556;

always @(posedge na1574)
   l130 <= na1574;

always @(posedge na1586)
   l132 <= na1586;

always @(posedge na1598)
   l134 <= na1598;

always @(posedge na1622)
   l136 <= na1622;

always @(posedge na1674)
   l138 <= na1674;

always @(posedge na1708)
   l140 <= na1708;

always @(posedge na1730)
   l142 <= na1730;

always @(posedge na1742)
   l144 <= na1742;

always @(posedge na1760)
   l146 <= na1760;

always @(posedge na1778)
   l148 <= na1778;

always @(posedge na1796)
   l150 <= na1796;

always @(posedge na1814)
   l152 <= na1814;

always @(posedge na1832)
   l154 <= na1832;

always @(posedge na1848)
   l156 <= na1848;

always @(posedge na1880)
   l158 <= na1880;

always @(posedge na1916)
   l160 <= na1916;

always @(posedge na1954)
   l162 <= na1954;

always @(posedge na1970)
   l164 <= na1970;

always @(posedge na1982)
   l166 <= na1982;

always @(posedge na2000)
   l168 <= na2000;

always @(posedge na2044)
   l170 <= na2044;

always @(posedge na2056)
   l172 <= na2056;

always @(posedge na2074)
   l174 <= na2074;

always @(posedge na2092)
   l176 <= na2092;

always @(posedge na2108)
   l178 <= na2108;

always @(posedge na2126)
   l180 <= na2126;

always @(posedge na2138)
   l182 <= na2138;

always @(posedge na2160)
   l184 <= na2160;

always @(posedge na2176)
   l186 <= na2176;

always @(posedge na2188)
   l188 <= na2188;

always @(posedge na2204)
   l190 <= na2204;

always @(posedge na2216)
   l192 <= na2216;

always @(posedge na2232)
   l194 <= na2232;

always @(posedge na2250)
   l196 <= na2250;

always @(posedge na1312)
   l198 <= na1312;

always @(posedge na2244)
   l200 <= na2244;

always @(posedge na2226)
   l202 <= na2226;

always @(posedge na2210)
   l204 <= na2210;

always @(posedge na2264)
   l206 <= na2264;

always @(posedge na2198)
   l208 <= na2198;

always @(posedge na2258)
   l210 <= na2258;

always @(posedge na2182)
   l212 <= na2182;

always @(posedge na2278)
   l214 <= na2278;

always @(posedge na2170)
   l216 <= na2170;

always @(posedge na2292)
   l218 <= na2292;

always @(posedge na2306)
   l220 <= na2306;

always @(posedge na2272)
   l222 <= na2272;

always @(posedge na2300)
   l224 <= na2300;

always @(posedge na2286)
   l226 <= na2286;

always @(posedge na2154)
   l228 <= na2154;

always @(posedge na2132)
   l230 <= na2132;

always @(posedge na2120)
   l232 <= na2120;

always @(posedge na2102)
   l234 <= na2102;

always @(posedge na2324)
   l236 <= na2324;

always @(posedge na2346)
   l238 <= na2346;

always @(posedge na2086)
   l240 <= na2086;

always @(posedge na2340)
   l242 <= na2340;

always @(posedge na2364)
   l244 <= na2364;

always @(posedge na2318)
   l246 <= na2318;

always @(posedge na2358)
   l248 <= na2358;

always @(posedge na2068)
   l250 <= na2068;

always @(posedge na2050)
   l252 <= na2050;

always @(posedge na2388)
   l254 <= na2388;

always @(posedge na2400)
   l256 <= na2400;

always @(posedge na2412)
   l258 <= na2412;

always @(posedge na2424)
   l260 <= na2424;

always @(posedge na2436)
   l262 <= na2436;

always @(posedge na2448)
   l264 <= na2448;

always @(posedge na2466)
   l266 <= na2466;

always @(posedge na2482)
   l268 <= na2482;

always @(posedge na2038)
   l270 <= na2038;

always @(posedge na2476)
   l272 <= na2476;

always @(posedge na2460)
   l274 <= na2460;

always @(posedge na2494)
   l276 <= na2494;

always @(posedge na2442)
   l278 <= na2442;

always @(posedge na2506)
   l280 <= na2506;

always @(posedge na2488)
   l282 <= na2488;

always @(posedge na2518)
   l284 <= na2518;

always @(posedge na2500)
   l286 <= na2500;

always @(posedge na2530)
   l288 <= na2530;

always @(posedge na2512)
   l290 <= na2512;

always @(posedge na2542)
   l292 <= na2542;

always @(posedge na2524)
   l294 <= na2524;

always @(posedge na2554)
   l296 <= na2554;

always @(posedge na2536)
   l298 <= na2536;

always @(posedge na2570)
   l300 <= na2570;

always @(posedge na2548)
   l302 <= na2548;

always @(posedge na2582)
   l304 <= na2582;

always @(posedge na2564)
   l306 <= na2564;

always @(posedge na2594)
   l308 <= na2594;

always @(posedge na2576)
   l310 <= na2576;

always @(posedge na2606)
   l312 <= na2606;

always @(posedge na2588)
   l314 <= na2588;

always @(posedge na2618)
   l316 <= na2618;

always @(posedge na2600)
   l318 <= na2600;

always @(posedge na2612)
   l320 <= na2612;

always @(posedge na2430)
   l322 <= na2430;

always @(posedge na2418)
   l324 <= na2418;

always @(posedge na2406)
   l326 <= na2406;

always @(posedge na2394)
   l328 <= na2394;

always @(posedge na2382)
   l330 <= na2382;

always @(posedge na1994)
   l332 <= na1994;

always @(posedge na1976)
   l334 <= na1976;

always @(posedge na2636)
   l336 <= na2636;

always @(posedge na1964)
   l338 <= na1964;

always @(posedge na2658)
   l340 <= na2658;

always @(posedge na2630)
   l342 <= na2630;

always @(posedge na2652)
   l344 <= na2652;

always @(posedge na2708)
   l346 <= na2708;

always @(posedge na2738)
   l348 <= na2738;

always @(posedge na2764)
   l350 <= na2764;

always @(posedge na2784)
   l352 <= na2784;

always @(posedge na1948)
   l354 <= na1948;

always @(posedge na2778)
   l356 <= na2778;

always @(posedge na2796)
   l358 <= na2796;

always @(posedge na2758)
   l360 <= na2758;

always @(posedge na2790)
   l362 <= na2790;

always @(posedge na2732)
   l364 <= na2732;

always @(posedge na2702)
   l366 <= na2702;

always @(posedge na1910)
   l368 <= na1910;

always @(posedge na1874)
   l370 <= na1874;

always @(posedge na1842)
   l372 <= na1842;

always @(posedge na1826)
   l374 <= na1826;

always @(posedge na1808)
   l376 <= na1808;

always @(posedge na1790)
   l378 <= na1790;

always @(posedge na1772)
   l380 <= na1772;

always @(posedge na1754)
   l382 <= na1754;

always @(posedge na1736)
   l384 <= na1736;

always @(posedge na2830)
   l386 <= na2830;

always @(posedge na2860)
   l388 <= na2860;

always @(posedge na2886)
   l390 <= na2886;

always @(posedge na2912)
   l392 <= na2912;

always @(posedge na2942)
   l394 <= na2942;

always @(posedge na2964)
   l396 <= na2964;

always @(posedge na2986)
   l398 <= na2986;

always @(posedge na3004)
   l400 <= na3004;

always @(posedge na3026)
   l402 <= na3026;

always @(posedge na1724)
   l404 <= na1724;

always @(posedge na3020)
   l406 <= na3020;

always @(posedge na2998)
   l408 <= na2998;

always @(posedge na2980)
   l410 <= na2980;

always @(posedge na2958)
   l412 <= na2958;

always @(posedge na2936)
   l414 <= na2936;

always @(posedge na2906)
   l416 <= na2906;

always @(posedge na2880)
   l418 <= na2880;

always @(posedge na2854)
   l420 <= na2854;

always @(posedge na2824)
   l422 <= na2824;

always @(posedge na1702)
   l424 <= na1702;

always @(posedge na1668)
   l426 <= na1668;

always @(posedge na1616)
   l428 <= na1616;

always @(posedge na1592)
   l430 <= na1592;

always @(posedge na1580)
   l432 <= na1580;

always @(posedge na1568)
   l434 <= na1568;

always @(posedge na1550)
   l436 <= na1550;

always @(posedge na1532)
   l438 <= na1532;

always @(posedge na1514)
   l440 <= na1514;

always @(posedge na1496)
   l442 <= na1496;

always @(posedge na1478)
   l444 <= na1478;

always @(posedge na1460)
   l446 <= na1460;

always @(posedge na1442)
   l448 <= na1442;

always @(posedge na1424)
   l450 <= na1424;

always @(posedge na1396)
   l452 <= na1396;

always @(posedge na1378)
   l454 <= na1378;

always @(posedge na1360)
   l456 <= na1360;

always @(posedge na856)
   l458 <= na856;

always @(posedge na3044)
   l460 <= na3044;

always @(posedge na3062)
   l462 <= na3062;

always @(posedge na826)
   l464 <= na826;

always @(posedge na3056)
   l466 <= na3056;

always @(posedge a3038)
   l468 <= a3038;

always @(posedge na3450)
   l470 <= na3450;

always @(posedge na3466)
   l472 <= na3466;

always @(posedge na3470)
   l474 <= na3470;

always @(posedge na3460)
   l476 <= na3460;

always @(posedge na3482)
   l478 <= na3482;

always @(posedge na3500)
   l480 <= na3500;

always @(posedge na3518)
   l482 <= na3518;

always @(posedge na3536)
   l484 <= na3536;

always @(posedge na3554)
   l486 <= na3554;

always @(posedge na3572)
   l488 <= na3572;

always @(posedge na3590)
   l490 <= na3590;

always @(posedge na3608)
   l492 <= na3608;

always @(posedge na3626)
   l494 <= na3626;

always @(posedge na3644)
   l496 <= na3644;

always @(posedge na3662)
   l498 <= na3662;

always @(posedge na3680)
   l500 <= na3680;

always @(posedge na3692)
   l502 <= na3692;

always @(posedge na3742)
   l504 <= na3742;

always @(posedge na3754)
   l506 <= na3754;

always @(posedge na3778)
   l508 <= na3778;

always @(posedge na3818)
   l510 <= na3818;

always @(posedge na3836)
   l512 <= na3836;

always @(posedge na3848)
   l514 <= na3848;

always @(posedge na3866)
   l516 <= na3866;

always @(posedge na3884)
   l518 <= na3884;

always @(posedge na3902)
   l520 <= na3902;

always @(posedge na3920)
   l522 <= na3920;

always @(posedge na3938)
   l524 <= na3938;

always @(posedge na3954)
   l526 <= na3954;

always @(posedge na3992)
   l528 <= na3992;

always @(posedge na4026)
   l530 <= na4026;

always @(posedge na4050)
   l532 <= na4050;

always @(posedge na4066)
   l534 <= na4066;

always @(posedge na4072)
   l536 <= na4072;

always @(posedge na4090)
   l538 <= na4090;

always @(posedge na4130)
   l540 <= na4130;

always @(posedge na4142)
   l542 <= na4142;

always @(posedge na4160)
   l544 <= na4160;

always @(posedge na4176)
   l546 <= na4176;

always @(posedge na4194)
   l548 <= na4194;

always @(posedge na4206)
   l550 <= na4206;

always @(posedge na4228)
   l552 <= na4228;

always @(posedge na4244)
   l554 <= na4244;

always @(posedge na4250)
   l556 <= na4250;

always @(posedge na4266)
   l558 <= na4266;

always @(posedge na4272)
   l560 <= na4272;

always @(posedge na4288)
   l562 <= na4288;

always @(posedge na4306)
   l564 <= na4306;

always @(posedge na3444)
   l566 <= na3444;

always @(posedge na4300)
   l568 <= na4300;

always @(posedge na4282)
   l570 <= na4282;

always @(posedge na4320)
   l572 <= na4320;

always @(posedge na4260)
   l574 <= na4260;

always @(posedge na4314)
   l576 <= na4314;

always @(posedge na4334)
   l578 <= na4334;

always @(posedge na4238)
   l580 <= na4238;

always @(posedge na4348)
   l582 <= na4348;

always @(posedge na4362)
   l584 <= na4362;

always @(posedge na4328)
   l586 <= na4328;

always @(posedge na4356)
   l588 <= na4356;

always @(posedge na4342)
   l590 <= na4342;

always @(posedge na4222)
   l592 <= na4222;

always @(posedge na4200)
   l594 <= na4200;

always @(posedge na4188)
   l596 <= na4188;

always @(posedge na4170)
   l598 <= na4170;

always @(posedge na4380)
   l600 <= na4380;

always @(posedge na4402)
   l602 <= na4402;

always @(posedge na4154)
   l604 <= na4154;

always @(posedge na4396)
   l606 <= na4396;

always @(posedge na4420)
   l608 <= na4420;

always @(posedge na4374)
   l610 <= na4374;

always @(posedge na4414)
   l612 <= na4414;

always @(posedge na4136)
   l614 <= na4136;

always @(posedge na4426)
   l616 <= na4426;

always @(posedge na4442)
   l618 <= na4442;

always @(posedge na4448)
   l620 <= na4448;

always @(posedge na4454)
   l622 <= na4454;

always @(posedge na4460)
   l624 <= na4460;

always @(posedge na4472)
   l626 <= na4472;

always @(posedge na4492)
   l628 <= na4492;

always @(posedge na4510)
   l630 <= na4510;

always @(posedge na4124)
   l632 <= na4124;

always @(posedge na4504)
   l634 <= na4504;

always @(posedge na4486)
   l636 <= na4486;

always @(posedge na4522)
   l638 <= na4522;

always @(posedge na4466)
   l640 <= na4466;

always @(posedge na4534)
   l642 <= na4534;

always @(posedge na4516)
   l644 <= na4516;

always @(posedge na4546)
   l646 <= na4546;

always @(posedge na4528)
   l648 <= na4528;

always @(posedge na4558)
   l650 <= na4558;

always @(posedge na4540)
   l652 <= na4540;

always @(posedge na4570)
   l654 <= na4570;

always @(posedge na4552)
   l656 <= na4552;

always @(posedge na4582)
   l658 <= na4582;

always @(posedge na4564)
   l660 <= na4564;

always @(posedge na4594)
   l662 <= na4594;

always @(posedge na4576)
   l664 <= na4576;

always @(posedge na4606)
   l666 <= na4606;

always @(posedge na4588)
   l668 <= na4588;

always @(posedge na4618)
   l670 <= na4618;

always @(posedge na4600)
   l672 <= na4600;

always @(posedge na4630)
   l674 <= na4630;

always @(posedge na4612)
   l676 <= na4612;

always @(posedge na4642)
   l678 <= na4642;

always @(posedge na4624)
   l680 <= na4624;

always @(posedge na4636)
   l682 <= na4636;

always @(posedge na4436)
   l684 <= na4436;

always @(posedge na4084)
   l686 <= na4084;

always @(posedge na4660)
   l688 <= na4660;

always @(posedge na4060)
   l690 <= na4060;

always @(posedge na4682)
   l692 <= na4682;

always @(posedge na4654)
   l694 <= na4654;

always @(posedge na4676)
   l696 <= na4676;

always @(posedge na4720)
   l698 <= na4720;

always @(posedge na4752)
   l700 <= na4752;

always @(posedge na4772)
   l702 <= na4772;

always @(posedge na4798)
   l704 <= na4798;

always @(posedge na4044)
   l706 <= na4044;

always @(posedge na4792)
   l708 <= na4792;

always @(posedge na4766)
   l710 <= na4766;

always @(posedge na4746)
   l712 <= na4746;

always @(posedge na4804)
   l714 <= na4804;

always @(posedge na4714)
   l716 <= na4714;

always @(posedge na4020)
   l718 <= na4020;

always @(posedge na3986)
   l720 <= na3986;

always @(posedge na3948)
   l722 <= na3948;

always @(posedge na3932)
   l724 <= na3932;

always @(posedge na3914)
   l726 <= na3914;

always @(posedge na3896)
   l728 <= na3896;

always @(posedge na3878)
   l730 <= na3878;

always @(posedge na3860)
   l732 <= na3860;

always @(posedge na3842)
   l734 <= na3842;

always @(posedge na4838)
   l736 <= na4838;

always @(posedge na4868)
   l738 <= na4868;

always @(posedge na4894)
   l740 <= na4894;

always @(posedge na4920)
   l742 <= na4920;

always @(posedge na4950)
   l744 <= na4950;

always @(posedge na4972)
   l746 <= na4972;

always @(posedge na4994)
   l748 <= na4994;

always @(posedge na5012)
   l750 <= na5012;

always @(posedge na5034)
   l752 <= na5034;

always @(posedge na3830)
   l754 <= na3830;

always @(posedge na5028)
   l756 <= na5028;

always @(posedge na5006)
   l758 <= na5006;

always @(posedge na4988)
   l760 <= na4988;

always @(posedge na4966)
   l762 <= na4966;

always @(posedge na4944)
   l764 <= na4944;

always @(posedge na4914)
   l766 <= na4914;

always @(posedge na4888)
   l768 <= na4888;

always @(posedge na4862)
   l770 <= na4862;

always @(posedge na4832)
   l772 <= na4832;

always @(posedge na3812)
   l774 <= na3812;

always @(posedge na3772)
   l776 <= na3772;

always @(posedge na3748)
   l778 <= na3748;

always @(posedge na3736)
   l780 <= na3736;

always @(posedge na3686)
   l782 <= na3686;

always @(posedge na3674)
   l784 <= na3674;

always @(posedge na3656)
   l786 <= na3656;

always @(posedge na3638)
   l788 <= na3638;

always @(posedge na3620)
   l790 <= na3620;

always @(posedge na3602)
   l792 <= na3602;

always @(posedge na3584)
   l794 <= na3584;

always @(posedge na3566)
   l796 <= na3566;

always @(posedge na3548)
   l798 <= na3548;

always @(posedge na3530)
   l800 <= na3530;

always @(posedge na3512)
   l802 <= na3512;

always @(posedge na3494)
   l804 <= na3494;

always @(posedge na3476)
   l806 <= na3476;

always @(posedge c1)
   l808 <= c1;


assign na832 = ~a832;
assign na850 = ~a850;
assign na862 = ~a862;
assign na880 = ~a880;
assign na902 = ~a902;
assign na844 = ~a844;
assign na896 = ~a896;
assign a874 = ~a872 & ~a864;
assign na1318 = ~a1318;
assign na1334 = ~a1334;
assign na1342 = ~a1342;
assign na1336 = ~a1336;
assign na1354 = ~a1354;
assign na1328 = ~a1328;
assign na1348 = ~a1348;
assign na1366 = ~a1366;
assign na1384 = ~a1384;
assign na1402 = ~a1402;
assign na1430 = ~a1430;
assign na1448 = ~a1448;
assign na1466 = ~a1466;
assign na1484 = ~a1484;
assign na1502 = ~a1502;
assign na1520 = ~a1520;
assign na1538 = ~a1538;
assign na1556 = ~a1556;
assign na1574 = ~a1574;
assign na1586 = ~a1586;
assign na1598 = ~a1598;
assign na1622 = ~a1622;
assign na1674 = ~a1674;
assign na1708 = ~a1708;
assign na1730 = ~a1730;
assign na1742 = ~a1742;
assign na1760 = ~a1760;
assign na1778 = ~a1778;
assign na1796 = ~a1796;
assign na1814 = ~a1814;
assign na1832 = ~a1832;
assign na1848 = ~a1848;
assign na1880 = ~a1880;
assign na1916 = ~a1916;
assign na1954 = ~a1954;
assign na1970 = ~a1970;
assign na1982 = ~a1982;
assign na2000 = ~a2000;
assign na2044 = ~a2044;
assign na2056 = ~a2056;
assign na2074 = ~a2074;
assign na2092 = ~a2092;
assign na2108 = ~a2108;
assign na2126 = ~a2126;
assign na2138 = ~a2138;
assign na2160 = ~a2160;
assign na2176 = ~a2176;
assign na2188 = ~a2188;
assign na2204 = ~a2204;
assign na2216 = ~a2216;
assign na2232 = ~a2232;
assign na2250 = ~a2250;
assign na1312 = ~a1312;
assign na2244 = ~a2244;
assign na2226 = ~a2226;
assign na2210 = ~a2210;
assign na2264 = ~a2264;
assign na2198 = ~a2198;
assign na2258 = ~a2258;
assign na2182 = ~a2182;
assign na2278 = ~a2278;
assign na2170 = ~a2170;
assign na2292 = ~a2292;
assign na2306 = ~a2306;
assign na2272 = ~a2272;
assign na2300 = ~a2300;
assign na2286 = ~a2286;
assign na2154 = ~a2154;
assign na2132 = ~a2132;
assign na2120 = ~a2120;
assign na2102 = ~a2102;
assign na2324 = ~a2324;
assign na2346 = ~a2346;
assign na2086 = ~a2086;
assign na2340 = ~a2340;
assign na2364 = ~a2364;
assign na2318 = ~a2318;
assign na2358 = ~a2358;
assign na2068 = ~a2068;
assign na2050 = ~a2050;
assign na2388 = ~a2388;
assign na2400 = ~a2400;
assign na2412 = ~a2412;
assign na2424 = ~a2424;
assign na2436 = ~a2436;
assign na2448 = ~a2448;
assign na2466 = ~a2466;
assign na2482 = ~a2482;
assign na2038 = ~a2038;
assign na2476 = ~a2476;
assign na2460 = ~a2460;
assign na2494 = ~a2494;
assign na2442 = ~a2442;
assign na2506 = ~a2506;
assign na2488 = ~a2488;
assign na2518 = ~a2518;
assign na2500 = ~a2500;
assign na2530 = ~a2530;
assign na2512 = ~a2512;
assign na2542 = ~a2542;
assign na2524 = ~a2524;
assign na2554 = ~a2554;
assign na2536 = ~a2536;
assign na2570 = ~a2570;
assign na2548 = ~a2548;
assign na2582 = ~a2582;
assign na2564 = ~a2564;
assign na2594 = ~a2594;
assign na2576 = ~a2576;
assign na2606 = ~a2606;
assign na2588 = ~a2588;
assign na2618 = ~a2618;
assign na2600 = ~a2600;
assign na2612 = ~a2612;
assign na2430 = ~a2430;
assign na2418 = ~a2418;
assign na2406 = ~a2406;
assign na2394 = ~a2394;
assign na2382 = ~a2382;
assign na1994 = ~a1994;
assign na1976 = ~a1976;
assign na2636 = ~a2636;
assign na1964 = ~a1964;
assign na2658 = ~a2658;
assign na2630 = ~a2630;
assign na2652 = ~a2652;
assign na2708 = ~a2708;
assign na2738 = ~a2738;
assign na2764 = ~a2764;
assign na2784 = ~a2784;
assign na1948 = ~a1948;
assign na2778 = ~a2778;
assign na2796 = ~a2796;
assign na2758 = ~a2758;
assign na2790 = ~a2790;
assign na2732 = ~a2732;
assign na2702 = ~a2702;
assign na1910 = ~a1910;
assign na1874 = ~a1874;
assign na1842 = ~a1842;
assign na1826 = ~a1826;
assign na1808 = ~a1808;
assign na1790 = ~a1790;
assign na1772 = ~a1772;
assign na1754 = ~a1754;
assign na1736 = ~a1736;
assign na2830 = ~a2830;
assign na2860 = ~a2860;
assign na2886 = ~a2886;
assign na2912 = ~a2912;
assign na2942 = ~a2942;
assign na2964 = ~a2964;
assign na2986 = ~a2986;
assign na3004 = ~a3004;
assign na3026 = ~a3026;
assign na1724 = ~a1724;
assign na3020 = ~a3020;
assign na2998 = ~a2998;
assign na2980 = ~a2980;
assign na2958 = ~a2958;
assign na2936 = ~a2936;
assign na2906 = ~a2906;
assign na2880 = ~a2880;
assign na2854 = ~a2854;
assign na2824 = ~a2824;
assign na1702 = ~a1702;
assign na1668 = ~a1668;
assign na1616 = ~a1616;
assign na1592 = ~a1592;
assign na1580 = ~a1580;
assign na1568 = ~a1568;
assign na1550 = ~a1550;
assign na1532 = ~a1532;
assign na1514 = ~a1514;
assign na1496 = ~a1496;
assign na1478 = ~a1478;
assign na1460 = ~a1460;
assign na1442 = ~a1442;
assign na1424 = ~a1424;
assign na1396 = ~a1396;
assign na1378 = ~a1378;
assign na1360 = ~a1360;
assign na856 = ~a856;
assign na3044 = ~a3044;
assign na3062 = ~a3062;
assign na826 = ~a826;
assign na3056 = ~a3056;
assign a3038 = ~a3036 & ~a3028;
assign na3450 = ~a3450;
assign na3466 = ~a3466;
assign na3470 = ~a3470;
assign na3460 = ~a3460;
assign na3482 = ~a3482;
assign na3500 = ~a3500;
assign na3518 = ~a3518;
assign na3536 = ~a3536;
assign na3554 = ~a3554;
assign na3572 = ~a3572;
assign na3590 = ~a3590;
assign na3608 = ~a3608;
assign na3626 = ~a3626;
assign na3644 = ~a3644;
assign na3662 = ~a3662;
assign na3680 = ~a3680;
assign na3692 = ~a3692;
assign na3742 = ~a3742;
assign na3754 = ~a3754;
assign na3778 = ~a3778;
assign na3818 = ~a3818;
assign na3836 = ~a3836;
assign na3848 = ~a3848;
assign na3866 = ~a3866;
assign na3884 = ~a3884;
assign na3902 = ~a3902;
assign na3920 = ~a3920;
assign na3938 = ~a3938;
assign na3954 = ~a3954;
assign na3992 = ~a3992;
assign na4026 = ~a4026;
assign na4050 = ~a4050;
assign na4066 = ~a4066;
assign na4072 = ~a4072;
assign na4090 = ~a4090;
assign na4130 = ~a4130;
assign na4142 = ~a4142;
assign na4160 = ~a4160;
assign na4176 = ~a4176;
assign na4194 = ~a4194;
assign na4206 = ~a4206;
assign na4228 = ~a4228;
assign na4244 = ~a4244;
assign na4250 = ~a4250;
assign na4266 = ~a4266;
assign na4272 = ~a4272;
assign na4288 = ~a4288;
assign na4306 = ~a4306;
assign na3444 = ~a3444;
assign na4300 = ~a4300;
assign na4282 = ~a4282;
assign na4320 = ~a4320;
assign na4260 = ~a4260;
assign na4314 = ~a4314;
assign na4334 = ~a4334;
assign na4238 = ~a4238;
assign na4348 = ~a4348;
assign na4362 = ~a4362;
assign na4328 = ~a4328;
assign na4356 = ~a4356;
assign na4342 = ~a4342;
assign na4222 = ~a4222;
assign na4200 = ~a4200;
assign na4188 = ~a4188;
assign na4170 = ~a4170;
assign na4380 = ~a4380;
assign na4402 = ~a4402;
assign na4154 = ~a4154;
assign na4396 = ~a4396;
assign na4420 = ~a4420;
assign na4374 = ~a4374;
assign na4414 = ~a4414;
assign na4136 = ~a4136;
assign na4426 = ~a4426;
assign na4442 = ~a4442;
assign na4448 = ~a4448;
assign na4454 = ~a4454;
assign na4460 = ~a4460;
assign na4472 = ~a4472;
assign na4492 = ~a4492;
assign na4510 = ~a4510;
assign na4124 = ~a4124;
assign na4504 = ~a4504;
assign na4486 = ~a4486;
assign na4522 = ~a4522;
assign na4466 = ~a4466;
assign na4534 = ~a4534;
assign na4516 = ~a4516;
assign na4546 = ~a4546;
assign na4528 = ~a4528;
assign na4558 = ~a4558;
assign na4540 = ~a4540;
assign na4570 = ~a4570;
assign na4552 = ~a4552;
assign na4582 = ~a4582;
assign na4564 = ~a4564;
assign na4594 = ~a4594;
assign na4576 = ~a4576;
assign na4606 = ~a4606;
assign na4588 = ~a4588;
assign na4618 = ~a4618;
assign na4600 = ~a4600;
assign na4630 = ~a4630;
assign na4612 = ~a4612;
assign na4642 = ~a4642;
assign na4624 = ~a4624;
assign na4636 = ~a4636;
assign na4436 = ~a4436;
assign na4084 = ~a4084;
assign na4660 = ~a4660;
assign na4060 = ~a4060;
assign na4682 = ~a4682;
assign na4654 = ~a4654;
assign na4676 = ~a4676;
assign na4720 = ~a4720;
assign na4752 = ~a4752;
assign na4772 = ~a4772;
assign na4798 = ~a4798;
assign na4044 = ~a4044;
assign na4792 = ~a4792;
assign na4766 = ~a4766;
assign na4746 = ~a4746;
assign na4804 = ~a4804;
assign na4714 = ~a4714;
assign na4020 = ~a4020;
assign na3986 = ~a3986;
assign na3948 = ~a3948;
assign na3932 = ~a3932;
assign na3914 = ~a3914;
assign na3896 = ~a3896;
assign na3878 = ~a3878;
assign na3860 = ~a3860;
assign na3842 = ~a3842;
assign na4838 = ~a4838;
assign na4868 = ~a4868;
assign na4894 = ~a4894;
assign na4920 = ~a4920;
assign na4950 = ~a4950;
assign na4972 = ~a4972;
assign na4994 = ~a4994;
assign na5012 = ~a5012;
assign na5034 = ~a5034;
assign na3830 = ~a3830;
assign na5028 = ~a5028;
assign na5006 = ~a5006;
assign na4988 = ~a4988;
assign na4966 = ~a4966;
assign na4944 = ~a4944;
assign na4914 = ~a4914;
assign na4888 = ~a4888;
assign na4862 = ~a4862;
assign na4832 = ~a4832;
assign na3812 = ~a3812;
assign na3772 = ~a3772;
assign na3748 = ~a3748;
assign na3736 = ~a3736;
assign na3686 = ~a3686;
assign na3674 = ~a3674;
assign na3656 = ~a3656;
assign na3638 = ~a3638;
assign na3620 = ~a3620;
assign na3602 = ~a3602;
assign na3584 = ~a3584;
assign na3566 = ~a3566;
assign na3548 = ~a3548;
assign na3530 = ~a3530;
assign na3512 = ~a3512;
assign na3494 = ~a3494;
assign na3476 = ~a3476;
assign c1 = 1;
assign a810 = l78 & ~l76;
assign a812 = ~l78 & l76;
assign a814 = ~a812 & ~a810;
assign a816 = l460 & ~l82;
assign a818 = a816 & l80;
assign a820 = ~a818 & i2;
assign a822 = l462 & l80;
assign a824 = l464 & ~l80;
assign a826 = ~a824 & ~a822;
assign a828 = ~a826 & a820;
assign a830 = ~a820 & l76;
assign a832 = ~a830 & ~a828;
assign a834 = l84 & ~l82;
assign a836 = a834 & l80;
assign a838 = ~a836 & i2;
assign a840 = l86 & l80;
assign a842 = l88 & ~l80;
assign a844 = ~a842 & ~a840;
assign a846 = ~a844 & a838;
assign a848 = ~a838 & l78;
assign a850 = ~a848 & ~a846;
assign a852 = l80 & i74;
assign a854 = l458 & ~l80;
assign a856 = ~a854 & ~a852;
assign a858 = ~a856 & i2;
assign a860 = l82 & ~i2;
assign a862 = ~a860 & ~a858;
assign a864 = ~l92 & ~l80;
assign a866 = l96 & l94;
assign a868 = ~a866 & l80;
assign a870 = ~a834 & l98;
assign a872 = a870 & a868;
assign a876 = a874 & a838;
assign a878 = ~a838 & l84;
assign a880 = ~a878 & ~a876;
assign a882 = l80 & i4;
assign a884 = ~a882 & i2;
assign a886 = a834 & i6;
assign a888 = ~a834 & l86;
assign a890 = ~a888 & ~a886;
assign a892 = ~a890 & l80;
assign a894 = l90 & ~l80;
assign a896 = ~a894 & ~a892;
assign a898 = ~a896 & a884;
assign a900 = ~a884 & l86;
assign a902 = ~a900 & ~a898;
assign a904 = ~l112 & ~l110;
assign a906 = ~l118 & ~l116;
assign a908 = a906 & l114;
assign a910 = a908 & a904;
assign a912 = a906 & ~l114;
assign a914 = a904 & l120;
assign a916 = a914 & a912;
assign a918 = a912 & ~l120;
assign a920 = a918 & ~l110;
assign a922 = ~a920 & ~a916;
assign a924 = a922 & ~a910;
assign a926 = ~l124 & l122;
assign a928 = l128 & l126;
assign a930 = ~a928 & a926;
assign a932 = a930 & ~a924;
assign a934 = l124 & l122;
assign a936 = l118 & l116;
assign a938 = l120 & l114;
assign a940 = l112 & l110;
assign a942 = a940 & a938;
assign a944 = a942 & a936;
assign a946 = a944 & ~a934;
assign a948 = l130 & ~l126;
assign a950 = l124 & ~l122;
assign a952 = a950 & a948;
assign a954 = a952 & a910;
assign a956 = a954 & ~l128;
assign a958 = ~a956 & ~a946;
assign a960 = a958 & ~a932;
assign a962 = ~l144 & ~l142;
assign a964 = a962 & ~l140;
assign a966 = ~a964 & ~l138;
assign a968 = a918 & l110;
assign a970 = a968 & ~l112;
assign a972 = ~l152 & ~l150;
assign a974 = a972 & l148;
assign a976 = a974 & ~l146;
assign a978 = l154 & l146;
assign a980 = a972 & ~l148;
assign a982 = a980 & a978;
assign a984 = ~a982 & ~a976;
assign a986 = ~a984 & a970;
assign a988 = ~l154 & l146;
assign a990 = ~l152 & l150;
assign a992 = a990 & ~l148;
assign a994 = ~a992 & ~a974;
assign a996 = ~a994 & a988;
assign a998 = a996 & ~a924;
assign a1000 = ~a998 & ~a986;
assign a1002 = a1000 & a966;
assign a1004 = ~a970 & a924;
assign a1006 = ~a1004 & a926;
assign a1008 = a1006 & a1002;
assign a1010 = a1008 & l136;
assign a1012 = a952 & ~l128;
assign a1014 = ~a1012 & ~l122;
assign a1016 = ~a1014 & a970;
assign a1018 = ~a1016 & a924;
assign a1020 = a1018 & l102;
assign a1022 = l134 & ~l94;
assign a1024 = l156 & i8;
assign a1026 = ~a1024 & ~a1022;
assign a1028 = a1026 & ~a1020;
assign a1030 = a1028 & ~a1010;
assign a1032 = a1030 & ~l134;
assign a1034 = ~a944 & l102;
assign a1036 = ~a1034 & ~l96;
assign a1038 = ~a1036 & l142;
assign a1040 = a1038 & ~a1032;
assign a1042 = a1040 & l132;
assign a1044 = l160 & l158;
assign a1046 = a1044 & a1042;
assign a1048 = l162 & l160;
assign a1050 = a1048 & a1042;
assign a1052 = ~a1050 & ~a1046;
assign a1054 = ~a1052 & ~a960;
assign a1056 = l108 & ~l94;
assign a1058 = a1056 & ~a1054;
assign a1060 = l166 & l164;
assign a1062 = a928 & a926;
assign a1064 = ~a1062 & ~a934;
assign a1066 = a1064 & ~a952;
assign a1068 = ~a1066 & ~a922;
assign a1070 = a944 & a934;
assign a1072 = ~a1064 & a910;
assign a1074 = ~a1072 & ~a1070;
assign a1076 = a1074 & ~a1068;
assign a1078 = l118 & ~l110;
assign a1080 = a1078 & ~l116;
assign a1082 = a1080 & l112;
assign a1084 = a1078 & l116;
assign a1086 = a1084 & ~l114;
assign a1088 = ~l168 & ~l120;
assign a1090 = ~a1088 & l112;
assign a1092 = a1090 & a1086;
assign a1094 = ~a1092 & ~a1082;
assign a1096 = a938 & l112;
assign a1098 = a1096 & a1084;
assign a1100 = ~l124 & ~l122;
assign a1102 = ~l130 & l126;
assign a1104 = a1102 & a1100;
assign a1106 = a1104 & l120;
assign a1108 = a940 & a906;
assign a1110 = a1108 & l114;
assign a1112 = a1110 & ~a1106;
assign a1114 = ~a1112 & ~a968;
assign a1116 = a1114 & ~a1098;
assign a1118 = a1116 & a1094;
assign a1120 = a1108 & a938;
assign a1122 = a1082 & ~a938;
assign a1124 = ~a1122 & ~a1120;
assign a1126 = ~a1124 & a1104;
assign a1128 = a1086 & ~l112;
assign a1130 = a938 & ~l112;
assign a1132 = a1130 & a1080;
assign a1134 = ~a1132 & ~a1128;
assign a1136 = a1134 & ~a1126;
assign a1138 = a1136 & a1118;
assign a1140 = a1138 & a1076;
assign a1142 = a1140 & l102;
assign a1144 = ~a1142 & ~a1060;
assign a1146 = a1144 & ~a1058;
assign a1148 = a1146 & ~l108;
assign a1150 = l170 & l80;
assign a1152 = a1150 & a1040;
assign a1154 = a1152 & ~a1148;
assign a1156 = ~l130 & ~l126;
assign a1158 = a1156 & a934;
assign a1160 = a916 & ~l174;
assign a1162 = a1160 & a1158;
assign a1164 = ~a1104 & a1082;
assign a1166 = ~a1164 & a1116;
assign a1168 = a1166 & ~a1162;
assign a1170 = l128 & l122;
assign a1172 = a1170 & ~a1168;
assign a1174 = a926 & l130;
assign a1176 = ~a944 & a924;
assign a1178 = ~a1176 & ~l126;
assign a1180 = a1178 & a1174;
assign a1182 = a1174 & l126;
assign a1184 = a948 & a934;
assign a1186 = ~a1184 & ~a1182;
assign a1188 = ~a1186 & ~a924;
assign a1190 = a1188 & l128;
assign a1192 = ~a1190 & ~a1180;
assign a1194 = a1192 & ~a1172;
assign a1196 = ~a1194 & l158;
assign a1198 = a926 & ~l126;
assign a1200 = a1198 & l130;
assign a1202 = ~a1200 & ~a1126;
assign a1204 = ~a1202 & ~l158;
assign a1206 = ~a1204 & ~a1196;
assign a1208 = a990 & l148;
assign a1210 = a1206 & l154;
assign a1212 = ~a1210 & ~l146;
assign a1214 = ~a1212 & ~a978;
assign a1216 = a1214 & a1208;
assign a1218 = a966 & l176;
assign a1220 = a1218 & ~a1216;
assign a1222 = a1220 & ~a1206;
assign a1224 = ~a1046 & ~l94;
assign a1226 = a1224 & l172;
assign a1228 = l178 & i10;
assign a1230 = a934 & l180;
assign a1232 = ~a1230 & ~a926;
assign a1234 = ~a1232 & a1102;
assign a1236 = ~a1234 & ~a1158;
assign a1238 = a1236 & ~a1198;
assign a1240 = ~a1128 & a1094;
assign a1242 = ~a1240 & ~a1238;
assign a1244 = ~a1242 & ~a1126;
assign a1246 = a1244 & l102;
assign a1248 = ~a1246 & ~a1228;
assign a1250 = a1248 & ~a1226;
assign a1252 = a1250 & ~a1222;
assign a1254 = a1252 & ~l172;
assign a1256 = a1010 & l184;
assign a1258 = l182 & ~l94;
assign a1260 = l188 & l186;
assign a1262 = ~a1260 & ~a1258;
assign a1264 = a1242 & ~a1200;
assign a1266 = ~a1264 & a1020;
assign a1268 = ~a1266 & a1262;
assign a1270 = a1268 & ~a1256;
assign a1272 = a1270 & ~l182;
assign a1274 = ~a1206 & a1172;
assign a1276 = ~a1274 & a1046;
assign a1278 = ~a1276 & ~a1050;
assign a1280 = l132 & ~l94;
assign a1282 = a1280 & a1278;
assign a1284 = l192 & l190;
assign a1286 = ~l196 & ~l86;
assign a1288 = a1286 & l194;
assign a1290 = ~a1288 & ~a1284;
assign a1292 = ~a1128 & ~a1092;
assign a1294 = a1292 & a1168;
assign a1296 = a1294 & l102;
assign a1298 = ~a1296 & a1290;
assign a1300 = a1298 & ~a1282;
assign a1302 = a1300 & ~l132;
assign a1304 = ~a1302 & ~a1272;
assign a1306 = a1304 & ~a1254;
assign a1308 = a1306 & a1154;
assign a1310 = l198 & ~l80;
assign a1312 = ~a1310 & ~a1308;
assign a1314 = ~a1312 & a838;
assign a1316 = ~a838 & l94;
assign a1318 = ~a1316 & ~a1314;
assign a1320 = l96 & ~l94;
assign a1322 = ~a1320 & ~l102;
assign a1324 = ~a1322 & l80;
assign a1326 = l104 & ~l80;
assign a1328 = ~a1326 & ~a1324;
assign a1330 = ~a1328 & a838;
assign a1332 = ~a838 & l96;
assign a1334 = ~a1332 & ~a1330;
assign a1336 = ~l100 & ~l80;
assign a1338 = ~a1336 & a838;
assign a1340 = ~a838 & l98;
assign a1342 = ~a1340 & ~a1338;
assign a1344 = l82 & l80;
assign a1346 = l106 & ~l80;
assign a1348 = ~a1346 & ~a1344;
assign a1350 = ~a1348 & a838;
assign a1352 = ~a838 & l102;
assign a1354 = ~a1352 & ~a1350;
assign a1356 = ~a1146 & l80;
assign a1358 = l456 & ~l80;
assign a1360 = ~a1358 & ~a1356;
assign a1362 = ~a1360 & a838;
assign a1364 = ~a838 & l108;
assign a1366 = ~a1364 & ~a1362;
assign a1368 = a834 & i72;
assign a1370 = ~a834 & l110;
assign a1372 = ~a1370 & ~a1368;
assign a1374 = ~a1372 & l80;
assign a1376 = l454 & ~l80;
assign a1378 = ~a1376 & ~a1374;
assign a1380 = ~a1378 & a884;
assign a1382 = ~a884 & l110;
assign a1384 = ~a1382 & ~a1380;
assign a1386 = a834 & i70;
assign a1388 = ~a834 & l112;
assign a1390 = ~a1388 & ~a1386;
assign a1392 = ~a1390 & l80;
assign a1394 = l452 & ~l80;
assign a1396 = ~a1394 & ~a1392;
assign a1398 = ~a1396 & a884;
assign a1400 = ~a884 & l112;
assign a1402 = ~a1400 & ~a1398;
assign a1404 = i72 & i70;
assign a1406 = a1404 & i66;
assign a1408 = a1406 & i64;
assign a1410 = a1408 & i62;
assign a1412 = ~a1410 & i68;
assign a1414 = a1412 & a834;
assign a1416 = ~a834 & l114;
assign a1418 = ~a1416 & ~a1414;
assign a1420 = ~a1418 & l80;
assign a1422 = l450 & ~l80;
assign a1424 = ~a1422 & ~a1420;
assign a1426 = ~a1424 & a884;
assign a1428 = ~a884 & l114;
assign a1430 = ~a1428 & ~a1426;
assign a1432 = a834 & i66;
assign a1434 = ~a834 & l116;
assign a1436 = ~a1434 & ~a1432;
assign a1438 = ~a1436 & l80;
assign a1440 = l448 & ~l80;
assign a1442 = ~a1440 & ~a1438;
assign a1444 = ~a1442 & a884;
assign a1446 = ~a884 & l116;
assign a1448 = ~a1446 & ~a1444;
assign a1450 = a834 & i64;
assign a1452 = ~a834 & l118;
assign a1454 = ~a1452 & ~a1450;
assign a1456 = ~a1454 & l80;
assign a1458 = l446 & ~l80;
assign a1460 = ~a1458 & ~a1456;
assign a1462 = ~a1460 & a884;
assign a1464 = ~a884 & l118;
assign a1466 = ~a1464 & ~a1462;
assign a1468 = a834 & i62;
assign a1470 = ~a834 & l120;
assign a1472 = ~a1470 & ~a1468;
assign a1474 = ~a1472 & l80;
assign a1476 = l444 & ~l80;
assign a1478 = ~a1476 & ~a1474;
assign a1480 = ~a1478 & a884;
assign a1482 = ~a884 & l120;
assign a1484 = ~a1482 & ~a1480;
assign a1486 = a834 & i60;
assign a1488 = ~a834 & l122;
assign a1490 = ~a1488 & ~a1486;
assign a1492 = ~a1490 & l80;
assign a1494 = l442 & ~l80;
assign a1496 = ~a1494 & ~a1492;
assign a1498 = ~a1496 & a884;
assign a1500 = ~a884 & l122;
assign a1502 = ~a1500 & ~a1498;
assign a1504 = a834 & i58;
assign a1506 = ~a834 & l124;
assign a1508 = ~a1506 & ~a1504;
assign a1510 = ~a1508 & l80;
assign a1512 = l440 & ~l80;
assign a1514 = ~a1512 & ~a1510;
assign a1516 = ~a1514 & a884;
assign a1518 = ~a884 & l124;
assign a1520 = ~a1518 & ~a1516;
assign a1522 = a834 & i56;
assign a1524 = ~a834 & l126;
assign a1526 = ~a1524 & ~a1522;
assign a1528 = ~a1526 & l80;
assign a1530 = l438 & ~l80;
assign a1532 = ~a1530 & ~a1528;
assign a1534 = ~a1532 & a884;
assign a1536 = ~a884 & l126;
assign a1538 = ~a1536 & ~a1534;
assign a1540 = a834 & i54;
assign a1542 = ~a834 & l128;
assign a1544 = ~a1542 & ~a1540;
assign a1546 = ~a1544 & l80;
assign a1548 = l436 & ~l80;
assign a1550 = ~a1548 & ~a1546;
assign a1552 = ~a1550 & a884;
assign a1554 = ~a884 & l128;
assign a1556 = ~a1554 & ~a1552;
assign a1558 = a834 & i52;
assign a1560 = ~a834 & l130;
assign a1562 = ~a1560 & ~a1558;
assign a1564 = ~a1562 & l80;
assign a1566 = l434 & ~l80;
assign a1568 = ~a1566 & ~a1564;
assign a1570 = ~a1568 & a884;
assign a1572 = ~a884 & l130;
assign a1574 = ~a1572 & ~a1570;
assign a1576 = ~a1300 & l80;
assign a1578 = l432 & ~l80;
assign a1580 = ~a1578 & ~a1576;
assign a1582 = ~a1580 & a838;
assign a1584 = ~a838 & l132;
assign a1586 = ~a1584 & ~a1582;
assign a1588 = ~a1030 & l80;
assign a1590 = l430 & ~l80;
assign a1592 = ~a1590 & ~a1588;
assign a1594 = ~a1592 & a838;
assign a1596 = ~a838 & l134;
assign a1598 = ~a1596 & ~a1594;
assign a1600 = ~a1018 & l102;
assign a1602 = ~a1000 & a966;
assign a1604 = ~a1602 & a1006;
assign a1606 = a1604 & l136;
assign a1608 = a1606 & ~a1008;
assign a1610 = ~a1608 & ~a1600;
assign a1612 = ~a1610 & l80;
assign a1614 = l428 & ~l80;
assign a1616 = ~a1614 & ~a1612;
assign a1618 = ~a1616 & a838;
assign a1620 = ~a838 & l136;
assign a1622 = ~a1620 & ~a1618;
assign a1624 = a1216 & a966;
assign a1626 = a1624 & l176;
assign a1628 = a1626 & l144;
assign a1630 = l138 & i40;
assign a1632 = ~l236 & ~l218;
assign a1634 = a1632 & ~l244;
assign a1636 = a1634 & ~l178;
assign a1638 = ~a1636 & ~l176;
assign a1640 = ~a1638 & a1630;
assign a1642 = ~a1640 & l138;
assign a1644 = l124 & l112;
assign a1646 = ~a1644 & a968;
assign a1648 = ~a1646 & ~a1112;
assign a1650 = ~a1648 & l122;
assign a1652 = ~a1650 & a924;
assign a1654 = a1652 & a1244;
assign a1656 = ~a1654 & l102;
assign a1658 = ~a1656 & ~a1642;
assign a1660 = a1658 & ~a1046;
assign a1662 = a1660 & ~a1628;
assign a1664 = ~a1662 & l80;
assign a1666 = l426 & ~l80;
assign a1668 = ~a1666 & ~a1664;
assign a1670 = ~a1668 & a838;
assign a1672 = ~a838 & l138;
assign a1674 = ~a1672 & ~a1670;
assign a1676 = ~a1626 & l144;
assign a1678 = ~l388 & ~l386;
assign a1680 = ~l392 & ~l390;
assign a1682 = a1680 & a1678;
assign a1684 = ~l396 & ~l394;
assign a1686 = ~l400 & ~l398;
assign a1688 = a1686 & ~l402;
assign a1690 = a1688 & a1684;
assign a1692 = a1690 & a1682;
assign a1694 = ~a1692 & l140;
assign a1696 = ~a1694 & ~a1676;
assign a1698 = ~a1696 & l80;
assign a1700 = l424 & ~l80;
assign a1702 = ~a1700 & ~a1698;
assign a1704 = ~a1702 & a838;
assign a1706 = ~a838 & l140;
assign a1708 = ~a1706 & ~a1704;
assign a1710 = a1224 & l142;
assign a1712 = a1692 & l140;
assign a1714 = a1654 & l102;
assign a1716 = ~a1714 & ~a1712;
assign a1718 = a1716 & ~a1710;
assign a1720 = ~a1718 & l80;
assign a1722 = l404 & ~l80;
assign a1724 = ~a1722 & ~a1720;
assign a1726 = ~a1724 & a838;
assign a1728 = ~a838 & l142;
assign a1730 = ~a1728 & ~a1726;
assign a1732 = a1640 & l80;
assign a1734 = l384 & ~l80;
assign a1736 = ~a1734 & ~a1732;
assign a1738 = ~a1736 & a838;
assign a1740 = ~a838 & l144;
assign a1742 = ~a1740 & ~a1738;
assign a1744 = a1640 & i50;
assign a1746 = ~a1640 & l146;
assign a1748 = ~a1746 & ~a1744;
assign a1750 = ~a1748 & l80;
assign a1752 = l382 & ~l80;
assign a1754 = ~a1752 & ~a1750;
assign a1756 = ~a1754 & a838;
assign a1758 = ~a838 & l146;
assign a1760 = ~a1758 & ~a1756;
assign a1762 = a1640 & i48;
assign a1764 = ~a1640 & l148;
assign a1766 = ~a1764 & ~a1762;
assign a1768 = ~a1766 & l80;
assign a1770 = l380 & ~l80;
assign a1772 = ~a1770 & ~a1768;
assign a1774 = ~a1772 & a838;
assign a1776 = ~a838 & l148;
assign a1778 = ~a1776 & ~a1774;
assign a1780 = a1640 & i46;
assign a1782 = ~a1640 & l150;
assign a1784 = ~a1782 & ~a1780;
assign a1786 = ~a1784 & l80;
assign a1788 = l378 & ~l80;
assign a1790 = ~a1788 & ~a1786;
assign a1792 = ~a1790 & a838;
assign a1794 = ~a838 & l150;
assign a1796 = ~a1794 & ~a1792;
assign a1798 = a1640 & i44;
assign a1800 = ~a1640 & l152;
assign a1802 = ~a1800 & ~a1798;
assign a1804 = ~a1802 & l80;
assign a1806 = l376 & ~l80;
assign a1808 = ~a1806 & ~a1804;
assign a1810 = ~a1808 & a838;
assign a1812 = ~a838 & l152;
assign a1814 = ~a1812 & ~a1810;
assign a1816 = a1640 & i42;
assign a1818 = ~a1640 & l154;
assign a1820 = ~a1818 & ~a1816;
assign a1822 = ~a1820 & l80;
assign a1824 = l374 & ~l80;
assign a1826 = ~a1824 & ~a1822;
assign a1828 = ~a1826 & a838;
assign a1830 = ~a838 & l154;
assign a1832 = ~a1830 & ~a1828;
assign a1834 = l156 & ~i8;
assign a1836 = ~a1834 & ~l220;
assign a1838 = ~a1836 & l80;
assign a1840 = l372 & ~l80;
assign a1842 = ~a1840 & ~a1838;
assign a1844 = ~a1842 & a838;
assign a1846 = ~a838 & l156;
assign a1848 = ~a1846 & ~a1844;
assign a1850 = l350 & l346;
assign a1852 = ~l348 & ~l346;
assign a1854 = ~a1852 & ~l352;
assign a1856 = a1854 & ~a1850;
assign a1858 = a1856 & ~a1018;
assign a1860 = ~a1238 & a944;
assign a1862 = ~a1860 & l264;
assign a1864 = a1862 & ~a1858;
assign a1866 = ~l264 & ~l158;
assign a1868 = ~a1866 & a868;
assign a1870 = a1868 & ~a1864;
assign a1872 = l370 & ~l80;
assign a1874 = ~a1872 & ~a1870;
assign a1876 = ~a1874 & a838;
assign a1878 = ~a838 & l158;
assign a1880 = ~a1878 & ~a1876;
assign a1882 = ~a1244 & l258;
assign a1884 = ~l262 & ~l258;
assign a1886 = a1884 & ~l260;
assign a1888 = a1176 & ~a1016;
assign a1890 = ~a1888 & ~a1886;
assign a1892 = ~a1890 & ~a1882;
assign a1894 = l266 & l264;
assign a1896 = a1894 & ~a1892;
assign a1898 = ~l162 & ~l158;
assign a1900 = ~a1898 & l160;
assign a1902 = a1900 & ~a1042;
assign a1904 = ~a1902 & ~a1896;
assign a1906 = ~a1904 & l80;
assign a1908 = l368 & ~l80;
assign a1910 = ~a1908 & ~a1906;
assign a1912 = ~a1910 & a838;
assign a1914 = ~a838 & l160;
assign a1916 = ~a1914 & ~a1912;
assign a1918 = l352 & ~l350;
assign a1920 = a1918 & a1852;
assign a1922 = ~l352 & l348;
assign a1924 = a1922 & a1850;
assign a1926 = ~a1924 & ~a1920;
assign a1928 = ~a1926 & ~a1018;
assign a1930 = a1186 & ~a950;
assign a1932 = ~a1930 & a944;
assign a1934 = ~a954 & l264;
assign a1936 = a1934 & ~a1932;
assign a1938 = a1936 & ~a1928;
assign a1940 = ~l264 & ~l162;
assign a1942 = ~a1940 & a868;
assign a1944 = a1942 & ~a1938;
assign a1946 = l354 & ~l80;
assign a1948 = ~a1946 & ~a1944;
assign a1950 = ~a1948 & a838;
assign a1952 = ~a838 & l162;
assign a1954 = ~a1952 & ~a1950;
assign a1956 = ~l166 & l164;
assign a1958 = ~a1956 & ~l336;
assign a1960 = ~a1958 & l80;
assign a1962 = l338 & ~l80;
assign a1964 = ~a1962 & ~a1960;
assign a1966 = ~a1964 & a838;
assign a1968 = ~a838 & l164;
assign a1970 = ~a1968 & ~a1966;
assign a1972 = l80 & i36;
assign a1974 = l334 & ~l80;
assign a1976 = ~a1974 & ~a1972;
assign a1978 = ~a1976 & a838;
assign a1980 = ~a838 & l166;
assign a1982 = ~a1980 & ~a1978;
assign a1984 = a834 & i34;
assign a1986 = ~a834 & l168;
assign a1988 = ~a1986 & ~a1984;
assign a1990 = ~a1988 & l80;
assign a1992 = l332 & ~l80;
assign a1994 = ~a1992 & ~a1990;
assign a1996 = ~a1994 & a884;
assign a1998 = ~a884 & l168;
assign a2000 = ~a1998 & ~a1996;
assign a2002 = a1010 & l254;
assign a2004 = ~a1264 & a1018;
assign a2006 = a2004 & ~a944;
assign a2008 = ~a2006 & l256;
assign a2010 = ~a2008 & l102;
assign a2012 = ~a2010 & ~a2002;
assign a2014 = a1894 & a1892;
assign a2016 = ~l178 & ~l172;
assign a2018 = ~a2016 & l132;
assign a2020 = a2018 & l268;
assign a2022 = l170 & ~l94;
assign a2024 = a1898 & l160;
assign a2026 = ~a2024 & ~a2022;
assign a2028 = a2026 & ~a2020;
assign a2030 = a2028 & ~a2014;
assign a2032 = a2030 & a2012;
assign a2034 = ~a2032 & l80;
assign a2036 = l270 & ~l80;
assign a2038 = ~a2036 & ~a2034;
assign a2040 = ~a2038 & a838;
assign a2042 = ~a838 & l170;
assign a2044 = ~a2042 & ~a2040;
assign a2046 = ~a1252 & l80;
assign a2048 = l252 & ~l80;
assign a2050 = ~a2048 & ~a2046;
assign a2052 = ~a2050 & a838;
assign a2054 = ~a838 & l172;
assign a2056 = ~a2054 & ~a2052;
assign a2058 = l82 & i24;
assign a2060 = l174 & ~l82;
assign a2062 = ~a2060 & ~a2058;
assign a2064 = ~a2062 & l80;
assign a2066 = l250 & ~l80;
assign a2068 = ~a2066 & ~a2064;
assign a2070 = ~a2068 & a838;
assign a2072 = ~a838 & l174;
assign a2074 = ~a2072 & ~a2070;
assign a2076 = ~l238 & l236;
assign a2078 = ~a966 & l176;
assign a2080 = ~a2078 & ~a2076;
assign a2082 = ~a2080 & l80;
assign a2084 = l240 & ~l80;
assign a2086 = ~a2084 & ~a2082;
assign a2088 = ~a2086 & a838;
assign a2090 = ~a838 & l176;
assign a2092 = ~a2090 & ~a2088;
assign a2094 = l178 & ~i10;
assign a2096 = ~a2094 & ~l218;
assign a2098 = ~a2096 & l80;
assign a2100 = l234 & ~l80;
assign a2102 = ~a2100 & ~a2098;
assign a2104 = ~a2102 & a838;
assign a2106 = ~a838 & l178;
assign a2108 = ~a2106 & ~a2104;
assign a2110 = a834 & i18;
assign a2112 = ~a834 & l180;
assign a2114 = ~a2112 & ~a2110;
assign a2116 = ~a2114 & l80;
assign a2118 = l232 & ~l80;
assign a2120 = ~a2118 & ~a2116;
assign a2122 = ~a2120 & a884;
assign a2124 = ~a884 & l180;
assign a2126 = ~a2124 & ~a2122;
assign a2128 = ~a1270 & l80;
assign a2130 = l230 & ~l80;
assign a2132 = ~a2130 & ~a2128;
assign a2134 = ~a2132 & a838;
assign a2136 = ~a838 & l182;
assign a2138 = ~a2136 & ~a2134;
assign a2140 = ~a2004 & l82;
assign a2142 = ~l220 & ~l218;
assign a2144 = a2142 & l184;
assign a2146 = a2144 & ~a1010;
assign a2148 = ~a2146 & ~a2140;
assign a2150 = ~a2148 & l80;
assign a2152 = l228 & ~l80;
assign a2154 = ~a2152 & ~a2150;
assign a2156 = ~a2154 & a838;
assign a2158 = ~a838 & l184;
assign a2160 = ~a2158 & ~a2156;
assign a2162 = ~l188 & l186;
assign a2164 = ~a2162 & ~l214;
assign a2166 = ~a2164 & l80;
assign a2168 = l216 & ~l80;
assign a2170 = ~a2168 & ~a2166;
assign a2172 = ~a2170 & a838;
assign a2174 = ~a838 & l186;
assign a2176 = ~a2174 & ~a2172;
assign a2178 = l80 & i16;
assign a2180 = l212 & ~l80;
assign a2182 = ~a2180 & ~a2178;
assign a2184 = ~a2182 & a838;
assign a2186 = ~a838 & l188;
assign a2188 = ~a2186 & ~a2184;
assign a2190 = ~l192 & l190;
assign a2192 = ~a2190 & ~l206;
assign a2194 = ~a2192 & l80;
assign a2196 = l208 & ~l80;
assign a2198 = ~a2196 & ~a2194;
assign a2200 = ~a2198 & a838;
assign a2202 = ~a838 & l190;
assign a2204 = ~a2202 & ~a2200;
assign a2206 = l80 & i14;
assign a2208 = l204 & ~l80;
assign a2210 = ~a2208 & ~a2206;
assign a2212 = ~a2210 & a838;
assign a2214 = ~a838 & l192;
assign a2216 = ~a2214 & ~a2212;
assign a2218 = ~a1294 & l102;
assign a2220 = ~a2218 & a1278;
assign a2222 = ~a2220 & l80;
assign a2224 = l202 & ~l80;
assign a2226 = ~a2224 & ~a2222;
assign a2228 = ~a2226 & a838;
assign a2230 = ~a838 & l194;
assign a2232 = ~a2230 & ~a2228;
assign a2234 = a834 & i12;
assign a2236 = ~a834 & l196;
assign a2238 = ~a2236 & ~a2234;
assign a2240 = ~a2238 & l80;
assign a2242 = l200 & ~l80;
assign a2244 = ~a2242 & ~a2240;
assign a2246 = ~a2244 & a884;
assign a2248 = ~a884 & l196;
assign a2250 = ~a2248 & ~a2246;
assign a2252 = l194 & l80;
assign a2254 = a2252 & ~a1286;
assign a2256 = l210 & ~l80;
assign a2258 = ~a2256 & ~a2254;
assign a2260 = ~a2258 & a838;
assign a2262 = ~a838 & l206;
assign a2264 = ~a2262 & ~a2260;
assign a2266 = l184 & l80;
assign a2268 = a2266 & ~a2142;
assign a2270 = l222 & ~l80;
assign a2272 = ~a2270 & ~a2268;
assign a2274 = ~a2272 & a838;
assign a2276 = ~a838 & l214;
assign a2278 = ~a2276 & ~a2274;
assign a2280 = a1206 & l80;
assign a2282 = a2280 & a1220;
assign a2284 = l226 & ~l80;
assign a2286 = ~a2284 & ~a2282;
assign a2288 = ~a2286 & a838;
assign a2290 = ~a838 & l218;
assign a2292 = ~a2290 & ~a2288;
assign a2294 = l136 & l80;
assign a2296 = a2294 & ~a1604;
assign a2298 = l224 & ~l80;
assign a2300 = ~a2298 & ~a2296;
assign a2302 = ~a2300 & a838;
assign a2304 = ~a838 & l220;
assign a2306 = ~a2304 & ~a2302;
assign a2308 = l238 & l236;
assign a2310 = ~a2308 & ~l244;
assign a2312 = a2310 & ~a1626;
assign a2314 = ~a2312 & l80;
assign a2316 = l246 & ~l80;
assign a2318 = ~a2316 & ~a2314;
assign a2320 = ~a2318 & a838;
assign a2322 = ~a838 & l236;
assign a2324 = ~a2322 & ~a2320;
assign a2326 = a1624 & i20;
assign a2328 = ~a2326 & ~l238;
assign a2330 = ~a1624 & i22;
assign a2332 = ~l84 & l80;
assign a2334 = a2332 & ~a2330;
assign a2336 = a2334 & ~a2328;
assign a2338 = l242 & ~l80;
assign a2340 = ~a2338 & ~a2336;
assign a2342 = ~a2340 & a838;
assign a2344 = ~a838 & l238;
assign a2346 = ~a2344 & ~a2342;
assign a2348 = a1046 & l172;
assign a2350 = ~a1244 & l102;
assign a2352 = ~a2350 & ~a2348;
assign a2354 = ~a2352 & l80;
assign a2356 = l248 & ~l80;
assign a2358 = ~a2356 & ~a2354;
assign a2360 = ~a2358 & a838;
assign a2362 = ~a838 & l244;
assign a2364 = ~a2362 & ~a2360;
assign a2366 = a2008 & l102;
assign a2368 = ~a1272 & ~a1010;
assign a2370 = ~a2368 & ~a944;
assign a2372 = ~a1010 & l254;
assign a2374 = a2372 & a2370;
assign a2376 = ~a2374 & ~a2366;
assign a2378 = ~a2376 & l80;
assign a2380 = l330 & ~l80;
assign a2382 = ~a2380 & ~a2378;
assign a2384 = ~a2382 & a838;
assign a2386 = ~a838 & l254;
assign a2388 = ~a2386 & ~a2384;
assign a2390 = l80 & i32;
assign a2392 = l328 & ~l80;
assign a2394 = ~a2392 & ~a2390;
assign a2396 = ~a2394 & a838;
assign a2398 = ~a838 & l256;
assign a2400 = ~a2398 & ~a2396;
assign a2402 = l80 & i30;
assign a2404 = l326 & ~l80;
assign a2406 = ~a2404 & ~a2402;
assign a2408 = ~a2406 & a838;
assign a2410 = ~a838 & l258;
assign a2412 = ~a2410 & ~a2408;
assign a2414 = l80 & i28;
assign a2416 = l324 & ~l80;
assign a2418 = ~a2416 & ~a2414;
assign a2420 = ~a2418 & a838;
assign a2422 = ~a838 & l260;
assign a2424 = ~a2422 & ~a2420;
assign a2426 = l80 & i26;
assign a2428 = l322 & ~l80;
assign a2430 = ~a2428 & ~a2426;
assign a2432 = ~a2430 & a838;
assign a2434 = ~a838 & l262;
assign a2436 = ~a2434 & ~a2432;
assign a2438 = l276 & l80;
assign a2440 = l278 & ~l80;
assign a2442 = ~a2440 & ~a2438;
assign a2444 = ~a2442 & a838;
assign a2446 = ~a838 & l264;
assign a2448 = ~a2446 & ~a2444;
assign a2450 = ~a2370 & l254;
assign a2452 = l266 & ~l264;
assign a2454 = ~a2452 & ~a2450;
assign a2456 = ~a2454 & l80;
assign a2458 = l274 & ~l80;
assign a2460 = ~a2458 & ~a2456;
assign a2462 = ~a2460 & a838;
assign a2464 = ~a838 & l266;
assign a2466 = ~a2464 & ~a2462;
assign a2468 = ~a2018 & l268;
assign a2470 = ~a2468 & a1052;
assign a2472 = ~a2470 & l80;
assign a2474 = l272 & ~l80;
assign a2476 = ~a2474 & ~a2472;
assign a2478 = ~a2476 & a838;
assign a2480 = ~a838 & l268;
assign a2482 = ~a2480 & ~a2478;
assign a2484 = l280 & l80;
assign a2486 = l282 & ~l80;
assign a2488 = ~a2486 & ~a2484;
assign a2490 = ~a2488 & a838;
assign a2492 = ~a838 & l276;
assign a2494 = ~a2492 & ~a2490;
assign a2496 = l284 & l80;
assign a2498 = l286 & ~l80;
assign a2500 = ~a2498 & ~a2496;
assign a2502 = ~a2500 & a838;
assign a2504 = ~a838 & l280;
assign a2506 = ~a2504 & ~a2502;
assign a2508 = l288 & l80;
assign a2510 = l290 & ~l80;
assign a2512 = ~a2510 & ~a2508;
assign a2514 = ~a2512 & a838;
assign a2516 = ~a838 & l284;
assign a2518 = ~a2516 & ~a2514;
assign a2520 = l292 & l80;
assign a2522 = l294 & ~l80;
assign a2524 = ~a2522 & ~a2520;
assign a2526 = ~a2524 & a838;
assign a2528 = ~a838 & l288;
assign a2530 = ~a2528 & ~a2526;
assign a2532 = l296 & l80;
assign a2534 = l298 & ~l80;
assign a2536 = ~a2534 & ~a2532;
assign a2538 = ~a2536 & a838;
assign a2540 = ~a838 & l292;
assign a2542 = ~a2540 & ~a2538;
assign a2544 = l300 & l80;
assign a2546 = l302 & ~l80;
assign a2548 = ~a2546 & ~a2544;
assign a2550 = ~a2548 & a838;
assign a2552 = ~a838 & l296;
assign a2554 = ~a2552 & ~a2550;
assign a2556 = a944 & l102;
assign a2558 = ~a2556 & ~l304;
assign a2560 = ~a2558 & l80;
assign a2562 = l306 & ~l80;
assign a2564 = ~a2562 & ~a2560;
assign a2566 = ~a2564 & a838;
assign a2568 = ~a838 & l300;
assign a2570 = ~a2568 & ~a2566;
assign a2572 = l308 & l80;
assign a2574 = l310 & ~l80;
assign a2576 = ~a2574 & ~a2572;
assign a2578 = ~a2576 & a838;
assign a2580 = ~a838 & l304;
assign a2582 = ~a2580 & ~a2578;
assign a2584 = l312 & l80;
assign a2586 = l314 & ~l80;
assign a2588 = ~a2586 & ~a2584;
assign a2590 = ~a2588 & a838;
assign a2592 = ~a838 & l308;
assign a2594 = ~a2592 & ~a2590;
assign a2596 = l316 & l80;
assign a2598 = l318 & ~l80;
assign a2600 = ~a2598 & ~a2596;
assign a2602 = ~a2600 & a838;
assign a2604 = ~a838 & l312;
assign a2606 = ~a2604 & ~a2602;
assign a2608 = a2450 & l80;
assign a2610 = l320 & ~l80;
assign a2612 = ~a2610 & ~a2608;
assign a2614 = ~a2612 & a838;
assign a2616 = ~a838 & l316;
assign a2618 = ~a2616 & ~a2614;
assign a2620 = ~l268 & ~l170;
assign a2622 = ~a2620 & a1304;
assign a2624 = l340 & l80;
assign a2626 = a2624 & a2622;
assign a2628 = l342 & ~l80;
assign a2630 = ~a2628 & ~a2626;
assign a2632 = ~a2630 & a838;
assign a2634 = ~a838 & l336;
assign a2636 = ~a2634 & ~a2632;
assign a2638 = ~a2622 & l340;
assign a2640 = a1054 & l108;
assign a2642 = ~a1140 & l102;
assign a2644 = ~a2642 & ~a2640;
assign a2646 = a2644 & ~a2638;
assign a2648 = ~a2646 & l80;
assign a2650 = l344 & ~l80;
assign a2652 = ~a2650 & ~a2648;
assign a2654 = ~a2652 & a838;
assign a2656 = ~a838 & l340;
assign a2658 = ~a2656 & ~a2654;
assign a2660 = ~a1896 & l102;
assign a2662 = ~a1100 & ~l128;
assign a2664 = a2662 & ~a1168;
assign a2666 = ~a2664 & ~a1172;
assign a2668 = ~a1186 & a944;
assign a2670 = a1188 & ~l128;
assign a2672 = ~a2670 & ~a2668;
assign a2674 = ~a1236 & a944;
assign a2676 = ~a1160 & a1158;
assign a2678 = ~a2676 & ~a1234;
assign a2680 = ~a2678 & ~a924;
assign a2682 = a2680 & ~l128;
assign a2684 = ~a2682 & ~a2674;
assign a2686 = a2684 & a2672;
assign a2688 = a2686 & a2666;
assign a2690 = ~a2688 & a2660;
assign a2692 = ~a1896 & ~l102;
assign a2694 = a2692 & l346;
assign a2696 = ~a2694 & ~a2690;
assign a2698 = ~a2696 & l80;
assign a2700 = l366 & ~l80;
assign a2702 = ~a2700 & ~a2698;
assign a2704 = ~a2702 & a838;
assign a2706 = ~a838 & l346;
assign a2708 = ~a2706 & ~a2704;
assign a2710 = a2672 & a1192;
assign a2712 = a926 & ~l130;
assign a2714 = a2712 & a1178;
assign a2716 = ~a2714 & ~a2680;
assign a2718 = a2716 & ~a2674;
assign a2720 = a2718 & a2710;
assign a2722 = ~a2720 & a2660;
assign a2724 = a2692 & l348;
assign a2726 = ~a2724 & ~a2722;
assign a2728 = ~a2726 & l80;
assign a2730 = l364 & ~l80;
assign a2732 = ~a2730 & ~a2728;
assign a2734 = ~a2732 & a838;
assign a2736 = ~a838 & l348;
assign a2738 = ~a2736 & ~a2734;
assign a2740 = l358 & l258;
assign a2742 = a2740 & a1896;
assign a2744 = a2710 & ~a2664;
assign a2746 = ~a2744 & a2660;
assign a2748 = ~a2746 & ~a2742;
assign a2750 = a2692 & l350;
assign a2752 = ~a2750 & a2748;
assign a2754 = ~a2752 & l80;
assign a2756 = l360 & ~l80;
assign a2758 = ~a2756 & ~a2754;
assign a2760 = ~a2758 & a838;
assign a2762 = ~a838 & l350;
assign a2764 = ~a2762 & ~a2760;
assign a2766 = a952 & ~a924;
assign a2768 = a2766 & a2660;
assign a2770 = a2692 & l352;
assign a2772 = ~a2770 & ~a2768;
assign a2774 = ~a2772 & l80;
assign a2776 = l356 & ~l80;
assign a2778 = ~a2776 & ~a2774;
assign a2780 = ~a2778 & a838;
assign a2782 = ~a838 & l352;
assign a2784 = ~a2782 & ~a2780;
assign a2786 = l80 & i38;
assign a2788 = l362 & ~l80;
assign a2790 = ~a2788 & ~a2786;
assign a2792 = ~a2790 & a838;
assign a2794 = ~a838 & l358;
assign a2796 = ~a2794 & ~a2792;
assign a2798 = ~a1676 & ~l140;
assign a2800 = a2798 & l386;
assign a2802 = l386 & ~l144;
assign a2804 = l398 & ~l144;
assign a2806 = l400 & ~l144;
assign a2808 = ~a2806 & ~a2804;
assign a2810 = a2808 & ~a2802;
assign a2812 = ~a2808 & a2802;
assign a2814 = ~a2812 & ~a2810;
assign a2816 = ~a2814 & ~a2798;
assign a2818 = ~a2816 & ~a2800;
assign a2820 = ~a2818 & l80;
assign a2822 = l422 & ~l80;
assign a2824 = ~a2822 & ~a2820;
assign a2826 = ~a2824 & a838;
assign a2828 = ~a838 & l386;
assign a2830 = ~a2828 & ~a2826;
assign a2832 = a2798 & l388;
assign a2834 = l402 & ~l144;
assign a2836 = ~a2834 & a2810;
assign a2838 = l388 & ~l144;
assign a2840 = ~a2838 & a2836;
assign a2842 = a2838 & ~a2836;
assign a2844 = ~a2842 & ~a2840;
assign a2846 = ~a2844 & ~a2798;
assign a2848 = ~a2846 & ~a2832;
assign a2850 = ~a2848 & l80;
assign a2852 = l420 & ~l80;
assign a2854 = ~a2852 & ~a2850;
assign a2856 = ~a2854 & a838;
assign a2858 = ~a838 & l388;
assign a2860 = ~a2858 & ~a2856;
assign a2862 = a2798 & l390;
assign a2864 = l390 & ~l144;
assign a2866 = ~a2864 & a2840;
assign a2868 = a2864 & ~a2840;
assign a2870 = ~a2868 & ~a2866;
assign a2872 = ~a2870 & ~a2798;
assign a2874 = ~a2872 & ~a2862;
assign a2876 = ~a2874 & l80;
assign a2878 = l418 & ~l80;
assign a2880 = ~a2878 & ~a2876;
assign a2882 = ~a2880 & a838;
assign a2884 = ~a838 & l390;
assign a2886 = ~a2884 & ~a2882;
assign a2888 = a2798 & l392;
assign a2890 = l392 & ~l144;
assign a2892 = ~a2890 & a2866;
assign a2894 = a2890 & ~a2866;
assign a2896 = ~a2894 & ~a2892;
assign a2898 = ~a2896 & ~a2798;
assign a2900 = ~a2898 & ~a2888;
assign a2902 = ~a2900 & l80;
assign a2904 = l416 & ~l80;
assign a2906 = ~a2904 & ~a2902;
assign a2908 = ~a2906 & a838;
assign a2910 = ~a838 & l392;
assign a2912 = ~a2910 & ~a2908;
assign a2914 = a2798 & l394;
assign a2916 = l396 & ~l144;
assign a2918 = ~a2916 & a2892;
assign a2920 = l394 & ~l144;
assign a2922 = a2920 & ~a2918;
assign a2924 = ~a2920 & a2918;
assign a2926 = ~a2924 & ~a2922;
assign a2928 = ~a2926 & ~a2798;
assign a2930 = ~a2928 & ~a2914;
assign a2932 = ~a2930 & l80;
assign a2934 = l414 & ~l80;
assign a2936 = ~a2934 & ~a2932;
assign a2938 = ~a2936 & a838;
assign a2940 = ~a838 & l394;
assign a2942 = ~a2940 & ~a2938;
assign a2944 = a2798 & l396;
assign a2946 = a2916 & ~a2892;
assign a2948 = ~a2946 & ~a2918;
assign a2950 = ~a2948 & ~a2798;
assign a2952 = ~a2950 & ~a2944;
assign a2954 = ~a2952 & l80;
assign a2956 = l412 & ~l80;
assign a2958 = ~a2956 & ~a2954;
assign a2960 = ~a2958 & a838;
assign a2962 = ~a838 & l396;
assign a2964 = ~a2962 & ~a2960;
assign a2966 = a2798 & l398;
assign a2968 = a2804 & l400;
assign a2970 = ~a2968 & ~a2808;
assign a2972 = ~a2970 & ~a2798;
assign a2974 = ~a2972 & ~a2966;
assign a2976 = ~a2974 & l80;
assign a2978 = l410 & ~l80;
assign a2980 = ~a2978 & ~a2976;
assign a2982 = ~a2980 & a838;
assign a2984 = ~a838 & l398;
assign a2986 = ~a2984 & ~a2982;
assign a2988 = a2798 & l400;
assign a2990 = ~a2806 & ~a2798;
assign a2992 = ~a2990 & ~a2988;
assign a2994 = ~a2992 & l80;
assign a2996 = l408 & ~l80;
assign a2998 = ~a2996 & ~a2994;
assign a3000 = ~a2998 & a838;
assign a3002 = ~a838 & l400;
assign a3004 = ~a3002 & ~a3000;
assign a3006 = a2798 & l402;
assign a3008 = a2834 & ~a2810;
assign a3010 = ~a3008 & ~a2836;
assign a3012 = ~a3010 & ~a2798;
assign a3014 = ~a3012 & ~a3006;
assign a3016 = ~a3014 & l80;
assign a3018 = l406 & ~l80;
assign a3020 = ~a3018 & ~a3016;
assign a3022 = ~a3020 & a838;
assign a3024 = ~a838 & l402;
assign a3026 = ~a3024 & ~a3022;
assign a3028 = ~l468 & ~l80;
assign a3030 = l472 & l470;
assign a3032 = ~a3030 & l80;
assign a3034 = ~a816 & l98;
assign a3036 = a3034 & a3032;
assign a3040 = a3038 & a820;
assign a3042 = ~a820 & l460;
assign a3044 = ~a3042 & ~a3040;
assign a3046 = a816 & i6;
assign a3048 = ~a816 & l462;
assign a3050 = ~a3048 & ~a3046;
assign a3052 = ~a3050 & l80;
assign a3054 = l466 & ~l80;
assign a3056 = ~a3054 & ~a3052;
assign a3058 = ~a3056 & a884;
assign a3060 = ~a884 & l462;
assign a3062 = ~a3060 & ~a3058;
assign a3064 = ~l482 & ~l480;
assign a3066 = ~l488 & ~l486;
assign a3068 = a3066 & l484;
assign a3070 = a3068 & a3064;
assign a3072 = a3066 & ~l484;
assign a3074 = a3064 & l490;
assign a3076 = a3074 & a3072;
assign a3078 = a3072 & ~l490;
assign a3080 = a3078 & ~l482;
assign a3082 = ~a3080 & ~a3076;
assign a3084 = a3082 & ~a3070;
assign a3086 = ~l494 & l492;
assign a3088 = a3086 & ~a3084;
assign a3090 = l498 & l496;
assign a3092 = ~a3090 & a3088;
assign a3094 = l494 & ~l492;
assign a3096 = a3094 & ~l498;
assign a3098 = a3096 & l500;
assign a3100 = a3098 & ~l496;
assign a3102 = a3100 & a3070;
assign a3104 = ~a3102 & ~a3092;
assign a3106 = ~l514 & ~l504;
assign a3108 = a3106 & ~l512;
assign a3110 = ~a3108 & ~l510;
assign a3112 = a3078 & l482;
assign a3114 = a3112 & ~l480;
assign a3116 = ~l522 & ~l520;
assign a3118 = a3116 & l518;
assign a3120 = a3118 & ~l516;
assign a3122 = l524 & l516;
assign a3124 = a3116 & ~l518;
assign a3126 = a3124 & a3122;
assign a3128 = ~a3126 & ~a3120;
assign a3130 = ~a3128 & a3114;
assign a3132 = ~l524 & l516;
assign a3134 = ~l522 & l520;
assign a3136 = a3134 & ~l518;
assign a3138 = ~a3136 & ~a3118;
assign a3140 = ~a3138 & a3132;
assign a3142 = a3140 & ~a3084;
assign a3144 = ~a3142 & ~a3130;
assign a3146 = a3144 & a3110;
assign a3148 = ~a3114 & a3084;
assign a3150 = ~a3148 & a3086;
assign a3152 = a3150 & a3146;
assign a3154 = a3152 & l508;
assign a3156 = l506 & ~l470;
assign a3158 = l526 & i8;
assign a3160 = ~a3158 & ~a3156;
assign a3162 = ~a3100 & ~l492;
assign a3164 = ~a3162 & a3114;
assign a3166 = ~a3164 & a3084;
assign a3168 = a3166 & l474;
assign a3170 = ~a3168 & a3160;
assign a3172 = a3170 & ~a3154;
assign a3174 = a3172 & ~l506;
assign a3176 = ~a3174 & l504;
assign a3178 = a3176 & l502;
assign a3180 = l530 & l528;
assign a3182 = a3180 & a3178;
assign a3184 = l532 & l530;
assign a3186 = a3184 & a3178;
assign a3188 = ~a3186 & ~a3182;
assign a3190 = ~a3188 & ~a3104;
assign a3192 = l478 & ~l470;
assign a3194 = a3192 & ~a3190;
assign a3196 = l536 & l534;
assign a3198 = l494 & l492;
assign a3200 = a3090 & a3086;
assign a3202 = ~a3200 & ~a3198;
assign a3204 = a3098 & ~a3082;
assign a3206 = ~a3204 & a3202;
assign a3208 = ~a3206 & ~a3084;
assign a3210 = l488 & ~l482;
assign a3212 = a3210 & l486;
assign a3214 = l490 & l484;
assign a3216 = a3214 & l480;
assign a3218 = a3216 & a3212;
assign a3220 = ~l494 & ~l492;
assign a3222 = ~l500 & l498;
assign a3224 = a3222 & a3220;
assign a3226 = a3224 & l490;
assign a3228 = l482 & l480;
assign a3230 = a3228 & a3066;
assign a3232 = a3230 & l484;
assign a3234 = a3232 & ~a3226;
assign a3236 = ~a3234 & ~a3112;
assign a3238 = a3236 & ~a3218;
assign a3240 = a3210 & ~l486;
assign a3242 = a3240 & l480;
assign a3244 = a3212 & ~l484;
assign a3246 = ~l538 & ~l490;
assign a3248 = ~a3246 & l480;
assign a3250 = a3248 & a3244;
assign a3252 = ~a3250 & ~a3242;
assign a3254 = a3252 & a3238;
assign a3256 = a3230 & a3214;
assign a3258 = a3242 & ~a3214;
assign a3260 = ~a3258 & ~a3256;
assign a3262 = ~a3260 & a3224;
assign a3264 = a3244 & ~l480;
assign a3266 = a3214 & ~l480;
assign a3268 = a3266 & a3240;
assign a3270 = ~a3268 & ~a3264;
assign a3272 = a3270 & ~a3262;
assign a3274 = a3272 & a3254;
assign a3276 = a3274 & ~a3208;
assign a3278 = a3276 & l474;
assign a3280 = ~a3278 & ~a3196;
assign a3282 = a3280 & ~a3194;
assign a3284 = a3282 & ~l478;
assign a3286 = l540 & l80;
assign a3288 = a3286 & a3176;
assign a3290 = a3288 & ~a3284;
assign a3292 = a3198 & ~l498;
assign a3294 = a3292 & ~l500;
assign a3296 = a3076 & ~l174;
assign a3298 = a3296 & a3294;
assign a3300 = a3242 & ~a3224;
assign a3302 = ~a3300 & a3238;
assign a3304 = a3302 & ~a3298;
assign a3306 = l496 & l492;
assign a3308 = a3306 & ~a3304;
assign a3310 = a3086 & ~l498;
assign a3312 = ~a3084 & l500;
assign a3314 = a3312 & a3310;
assign a3316 = a3086 & l498;
assign a3318 = ~a3316 & ~a3292;
assign a3320 = ~a3318 & a3312;
assign a3322 = a3320 & l496;
assign a3324 = ~a3322 & ~a3314;
assign a3326 = a3324 & ~a3308;
assign a3328 = ~a3326 & l532;
assign a3330 = a3310 & l500;
assign a3332 = ~a3330 & ~a3262;
assign a3334 = ~a3332 & ~l532;
assign a3336 = ~a3334 & ~a3328;
assign a3338 = a3134 & l518;
assign a3340 = a3336 & l524;
assign a3342 = ~a3340 & ~l516;
assign a3344 = ~a3342 & ~a3122;
assign a3346 = a3344 & a3338;
assign a3348 = a3110 & l544;
assign a3350 = a3348 & ~a3346;
assign a3352 = a3350 & ~a3336;
assign a3354 = ~a3186 & ~l470;
assign a3356 = a3354 & l542;
assign a3358 = l546 & i10;
assign a3360 = a3198 & l548;
assign a3362 = ~a3360 & ~a3086;
assign a3364 = ~a3362 & a3222;
assign a3366 = ~a3310 & ~a3294;
assign a3368 = a3366 & ~a3364;
assign a3370 = ~a3264 & a3252;
assign a3372 = ~a3370 & ~a3368;
assign a3374 = ~a3372 & ~a3262;
assign a3376 = a3374 & l474;
assign a3378 = ~a3376 & ~a3358;
assign a3380 = a3378 & ~a3356;
assign a3382 = a3380 & ~a3352;
assign a3384 = a3382 & ~l542;
assign a3386 = a3154 & l552;
assign a3388 = l550 & ~l470;
assign a3390 = l556 & l554;
assign a3392 = ~a3390 & ~a3388;
assign a3394 = a3372 & ~a3330;
assign a3396 = ~a3394 & a3166;
assign a3398 = a3396 & l474;
assign a3400 = ~a3398 & a3392;
assign a3402 = a3400 & ~a3386;
assign a3404 = a3402 & ~l550;
assign a3406 = ~a3336 & a3308;
assign a3408 = ~a3406 & a3186;
assign a3410 = ~a3408 & ~a3182;
assign a3412 = l502 & ~l470;
assign a3414 = a3412 & a3410;
assign a3416 = l560 & l558;
assign a3418 = ~l564 & ~l462;
assign a3420 = a3418 & l562;
assign a3422 = ~a3420 & ~a3416;
assign a3424 = ~a3264 & ~a3250;
assign a3426 = a3424 & a3304;
assign a3428 = a3426 & l474;
assign a3430 = ~a3428 & a3422;
assign a3432 = a3430 & ~a3414;
assign a3434 = a3432 & ~l502;
assign a3436 = ~a3434 & ~a3404;
assign a3438 = a3436 & ~a3384;
assign a3440 = a3438 & a3290;
assign a3442 = l566 & ~l80;
assign a3444 = ~a3442 & ~a3440;
assign a3446 = ~a3444 & a820;
assign a3448 = ~a820 & l470;
assign a3450 = ~a3448 & ~a3446;
assign a3452 = l472 & ~l470;
assign a3454 = ~a3452 & ~l474;
assign a3456 = ~a3454 & l80;
assign a3458 = l476 & ~l80;
assign a3460 = ~a3458 & ~a3456;
assign a3462 = ~a3460 & a820;
assign a3464 = ~a820 & l472;
assign a3466 = ~a3464 & ~a3462;
assign a3468 = ~a820 & l474;
assign a3470 = ~a3468 & ~a1350;
assign a3472 = ~a3282 & l80;
assign a3474 = l806 & ~l80;
assign a3476 = ~a3474 & ~a3472;
assign a3478 = ~a3476 & a820;
assign a3480 = ~a820 & l478;
assign a3482 = ~a3480 & ~a3478;
assign a3484 = a816 & i70;
assign a3486 = ~a816 & l480;
assign a3488 = ~a3486 & ~a3484;
assign a3490 = ~a3488 & l80;
assign a3492 = l804 & ~l80;
assign a3494 = ~a3492 & ~a3490;
assign a3496 = ~a3494 & a884;
assign a3498 = ~a884 & l480;
assign a3500 = ~a3498 & ~a3496;
assign a3502 = a816 & i72;
assign a3504 = ~a816 & l482;
assign a3506 = ~a3504 & ~a3502;
assign a3508 = ~a3506 & l80;
assign a3510 = l802 & ~l80;
assign a3512 = ~a3510 & ~a3508;
assign a3514 = ~a3512 & a884;
assign a3516 = ~a884 & l482;
assign a3518 = ~a3516 & ~a3514;
assign a3520 = a1412 & a816;
assign a3522 = ~a816 & l484;
assign a3524 = ~a3522 & ~a3520;
assign a3526 = ~a3524 & l80;
assign a3528 = l800 & ~l80;
assign a3530 = ~a3528 & ~a3526;
assign a3532 = ~a3530 & a884;
assign a3534 = ~a884 & l484;
assign a3536 = ~a3534 & ~a3532;
assign a3538 = a816 & i66;
assign a3540 = ~a816 & l486;
assign a3542 = ~a3540 & ~a3538;
assign a3544 = ~a3542 & l80;
assign a3546 = l798 & ~l80;
assign a3548 = ~a3546 & ~a3544;
assign a3550 = ~a3548 & a884;
assign a3552 = ~a884 & l486;
assign a3554 = ~a3552 & ~a3550;
assign a3556 = a816 & i64;
assign a3558 = ~a816 & l488;
assign a3560 = ~a3558 & ~a3556;
assign a3562 = ~a3560 & l80;
assign a3564 = l796 & ~l80;
assign a3566 = ~a3564 & ~a3562;
assign a3568 = ~a3566 & a884;
assign a3570 = ~a884 & l488;
assign a3572 = ~a3570 & ~a3568;
assign a3574 = a816 & i62;
assign a3576 = ~a816 & l490;
assign a3578 = ~a3576 & ~a3574;
assign a3580 = ~a3578 & l80;
assign a3582 = l794 & ~l80;
assign a3584 = ~a3582 & ~a3580;
assign a3586 = ~a3584 & a884;
assign a3588 = ~a884 & l490;
assign a3590 = ~a3588 & ~a3586;
assign a3592 = a816 & i60;
assign a3594 = ~a816 & l492;
assign a3596 = ~a3594 & ~a3592;
assign a3598 = ~a3596 & l80;
assign a3600 = l792 & ~l80;
assign a3602 = ~a3600 & ~a3598;
assign a3604 = ~a3602 & a884;
assign a3606 = ~a884 & l492;
assign a3608 = ~a3606 & ~a3604;
assign a3610 = a816 & i58;
assign a3612 = ~a816 & l494;
assign a3614 = ~a3612 & ~a3610;
assign a3616 = ~a3614 & l80;
assign a3618 = l790 & ~l80;
assign a3620 = ~a3618 & ~a3616;
assign a3622 = ~a3620 & a884;
assign a3624 = ~a884 & l494;
assign a3626 = ~a3624 & ~a3622;
assign a3628 = a816 & i54;
assign a3630 = ~a816 & l496;
assign a3632 = ~a3630 & ~a3628;
assign a3634 = ~a3632 & l80;
assign a3636 = l788 & ~l80;
assign a3638 = ~a3636 & ~a3634;
assign a3640 = ~a3638 & a884;
assign a3642 = ~a884 & l496;
assign a3644 = ~a3642 & ~a3640;
assign a3646 = a816 & i56;
assign a3648 = ~a816 & l498;
assign a3650 = ~a3648 & ~a3646;
assign a3652 = ~a3650 & l80;
assign a3654 = l786 & ~l80;
assign a3656 = ~a3654 & ~a3652;
assign a3658 = ~a3656 & a884;
assign a3660 = ~a884 & l498;
assign a3662 = ~a3660 & ~a3658;
assign a3664 = a816 & i52;
assign a3666 = ~a816 & l500;
assign a3668 = ~a3666 & ~a3664;
assign a3670 = ~a3668 & l80;
assign a3672 = l784 & ~l80;
assign a3674 = ~a3672 & ~a3670;
assign a3676 = ~a3674 & a884;
assign a3678 = ~a884 & l500;
assign a3680 = ~a3678 & ~a3676;
assign a3682 = ~a3432 & l80;
assign a3684 = l782 & ~l80;
assign a3686 = ~a3684 & ~a3682;
assign a3688 = ~a3686 & a820;
assign a3690 = ~a820 & l502;
assign a3692 = ~a3690 & ~a3688;
assign a3694 = a3354 & l504;
assign a3696 = ~l738 & ~l736;
assign a3698 = ~l742 & ~l740;
assign a3700 = a3698 & a3696;
assign a3702 = ~l746 & ~l744;
assign a3704 = ~l750 & ~l748;
assign a3706 = a3704 & ~l752;
assign a3708 = a3706 & a3702;
assign a3710 = a3708 & a3700;
assign a3712 = a3710 & l512;
assign a3714 = l494 & l480;
assign a3716 = ~a3714 & a3112;
assign a3718 = ~a3716 & ~a3234;
assign a3720 = ~a3718 & l492;
assign a3722 = ~a3720 & a3084;
assign a3724 = a3722 & a3374;
assign a3726 = a3724 & l474;
assign a3728 = ~a3726 & ~a3712;
assign a3730 = a3728 & ~a3694;
assign a3732 = ~a3730 & l80;
assign a3734 = l780 & ~l80;
assign a3736 = ~a3734 & ~a3732;
assign a3738 = ~a3736 & a820;
assign a3740 = ~a820 & l504;
assign a3742 = ~a3740 & ~a3738;
assign a3744 = ~a3172 & l80;
assign a3746 = l778 & ~l80;
assign a3748 = ~a3746 & ~a3744;
assign a3750 = ~a3748 & a820;
assign a3752 = ~a820 & l506;
assign a3754 = ~a3752 & ~a3750;
assign a3756 = ~a3166 & l474;
assign a3758 = ~a3144 & a3110;
assign a3760 = ~a3758 & a3150;
assign a3762 = a3760 & l508;
assign a3764 = a3762 & ~a3152;
assign a3766 = ~a3764 & ~a3756;
assign a3768 = ~a3766 & l80;
assign a3770 = l776 & ~l80;
assign a3772 = ~a3770 & ~a3768;
assign a3774 = ~a3772 & a820;
assign a3776 = ~a820 & l508;
assign a3778 = ~a3776 & ~a3774;
assign a3780 = a3346 & a3110;
assign a3782 = a3780 & l544;
assign a3784 = a3782 & l514;
assign a3786 = l510 & i40;
assign a3788 = ~l600 & ~l582;
assign a3790 = a3788 & ~l608;
assign a3792 = a3790 & ~l546;
assign a3794 = ~a3792 & ~l544;
assign a3796 = ~a3794 & a3786;
assign a3798 = ~a3796 & l510;
assign a3800 = ~a3724 & l474;
assign a3802 = ~a3800 & ~a3798;
assign a3804 = a3802 & ~a3186;
assign a3806 = a3804 & ~a3784;
assign a3808 = ~a3806 & l80;
assign a3810 = l774 & ~l80;
assign a3812 = ~a3810 & ~a3808;
assign a3814 = ~a3812 & a820;
assign a3816 = ~a820 & l510;
assign a3818 = ~a3816 & ~a3814;
assign a3820 = ~a3782 & l514;
assign a3822 = ~a3710 & l512;
assign a3824 = ~a3822 & ~a3820;
assign a3826 = ~a3824 & l80;
assign a3828 = l754 & ~l80;
assign a3830 = ~a3828 & ~a3826;
assign a3832 = ~a3830 & a820;
assign a3834 = ~a820 & l512;
assign a3836 = ~a3834 & ~a3832;
assign a3838 = a3796 & l80;
assign a3840 = l734 & ~l80;
assign a3842 = ~a3840 & ~a3838;
assign a3844 = ~a3842 & a820;
assign a3846 = ~a820 & l514;
assign a3848 = ~a3846 & ~a3844;
assign a3850 = a3796 & i50;
assign a3852 = ~a3796 & l516;
assign a3854 = ~a3852 & ~a3850;
assign a3856 = ~a3854 & l80;
assign a3858 = l732 & ~l80;
assign a3860 = ~a3858 & ~a3856;
assign a3862 = ~a3860 & a820;
assign a3864 = ~a820 & l516;
assign a3866 = ~a3864 & ~a3862;
assign a3868 = a3796 & i48;
assign a3870 = ~a3796 & l518;
assign a3872 = ~a3870 & ~a3868;
assign a3874 = ~a3872 & l80;
assign a3876 = l730 & ~l80;
assign a3878 = ~a3876 & ~a3874;
assign a3880 = ~a3878 & a820;
assign a3882 = ~a820 & l518;
assign a3884 = ~a3882 & ~a3880;
assign a3886 = a3796 & i46;
assign a3888 = ~a3796 & l520;
assign a3890 = ~a3888 & ~a3886;
assign a3892 = ~a3890 & l80;
assign a3894 = l728 & ~l80;
assign a3896 = ~a3894 & ~a3892;
assign a3898 = ~a3896 & a820;
assign a3900 = ~a820 & l520;
assign a3902 = ~a3900 & ~a3898;
assign a3904 = a3796 & i44;
assign a3906 = ~a3796 & l522;
assign a3908 = ~a3906 & ~a3904;
assign a3910 = ~a3908 & l80;
assign a3912 = l726 & ~l80;
assign a3914 = ~a3912 & ~a3910;
assign a3916 = ~a3914 & a820;
assign a3918 = ~a820 & l522;
assign a3920 = ~a3918 & ~a3916;
assign a3922 = a3796 & i42;
assign a3924 = ~a3796 & l524;
assign a3926 = ~a3924 & ~a3922;
assign a3928 = ~a3926 & l80;
assign a3930 = l724 & ~l80;
assign a3932 = ~a3930 & ~a3928;
assign a3934 = ~a3932 & a820;
assign a3936 = ~a820 & l524;
assign a3938 = ~a3936 & ~a3934;
assign a3940 = l526 & ~i8;
assign a3942 = ~a3940 & ~l584;
assign a3944 = ~a3942 & l80;
assign a3946 = l722 & ~l80;
assign a3948 = ~a3946 & ~a3944;
assign a3950 = ~a3948 & a820;
assign a3952 = ~a820 & l526;
assign a3954 = ~a3952 & ~a3950;
assign a3956 = ~l704 & ~l700;
assign a3958 = l702 & ~l698;
assign a3960 = a3958 & a3956;
assign a3962 = l700 & l698;
assign a3964 = l704 & ~l702;
assign a3966 = a3964 & a3962;
assign a3968 = ~a3966 & ~a3960;
assign a3970 = ~a3968 & ~a3166;
assign a3972 = a3098 & a3070;
assign a3974 = ~a3972 & l626;
assign a3976 = a3974 & ~a3970;
assign a3978 = ~l626 & ~l528;
assign a3980 = ~a3978 & a3032;
assign a3982 = a3980 & ~a3976;
assign a3984 = l720 & ~l80;
assign a3986 = ~a3984 & ~a3982;
assign a3988 = ~a3986 & a820;
assign a3990 = ~a820 & l528;
assign a3992 = ~a3990 & ~a3988;
assign a3994 = ~a3374 & l620;
assign a3996 = ~l624 & ~l620;
assign a3998 = a3996 & ~l622;
assign a4000 = ~a3998 & ~a3166;
assign a4002 = ~a4000 & ~a3994;
assign a4004 = l628 & l626;
assign a4006 = a4004 & ~a4002;
assign a4008 = ~l532 & ~l528;
assign a4010 = ~a4008 & l530;
assign a4012 = a4010 & ~a3178;
assign a4014 = ~a4012 & ~a4006;
assign a4016 = ~a4014 & l80;
assign a4018 = l718 & ~l80;
assign a4020 = ~a4018 & ~a4016;
assign a4022 = ~a4020 & a820;
assign a4024 = ~a820 & l530;
assign a4026 = ~a4024 & ~a4022;
assign a4028 = ~a3956 & ~l702;
assign a4030 = a4028 & ~a3962;
assign a4032 = a4030 & ~a3166;
assign a4034 = ~a4032 & l626;
assign a4036 = ~l626 & ~l532;
assign a4038 = ~a4036 & a3032;
assign a4040 = a4038 & ~a4034;
assign a4042 = l706 & ~l80;
assign a4044 = ~a4042 & ~a4040;
assign a4046 = ~a4044 & a820;
assign a4048 = ~a820 & l532;
assign a4050 = ~a4048 & ~a4046;
assign a4052 = ~l536 & l534;
assign a4054 = ~a4052 & ~l688;
assign a4056 = ~a4054 & l80;
assign a4058 = l690 & ~l80;
assign a4060 = ~a4058 & ~a4056;
assign a4062 = ~a4060 & a820;
assign a4064 = ~a820 & l534;
assign a4066 = ~a4064 & ~a4062;
assign a4068 = ~a1976 & a820;
assign a4070 = ~a820 & l536;
assign a4072 = ~a4070 & ~a4068;
assign a4074 = a816 & i34;
assign a4076 = ~a816 & l538;
assign a4078 = ~a4076 & ~a4074;
assign a4080 = ~a4078 & l80;
assign a4082 = l686 & ~l80;
assign a4084 = ~a4082 & ~a4080;
assign a4086 = ~a4084 & a884;
assign a4088 = ~a884 & l538;
assign a4090 = ~a4088 & ~a4086;
assign a4092 = ~a3396 & l616;
assign a4094 = ~a4092 & l474;
assign a4096 = ~l546 & ~l542;
assign a4098 = ~a4096 & l502;
assign a4100 = a4098 & l618;
assign a4102 = l540 & ~l470;
assign a4104 = a4008 & l530;
assign a4106 = ~a4104 & ~a4102;
assign a4108 = a4106 & ~a4100;
assign a4110 = a4108 & ~a4094;
assign a4112 = a4004 & a4002;
assign a4114 = a3154 & l630;
assign a4116 = ~a4114 & ~a4112;
assign a4118 = a4116 & a4110;
assign a4120 = ~a4118 & l80;
assign a4122 = l632 & ~l80;
assign a4124 = ~a4122 & ~a4120;
assign a4126 = ~a4124 & a820;
assign a4128 = ~a820 & l540;
assign a4130 = ~a4128 & ~a4126;
assign a4132 = ~a3382 & l80;
assign a4134 = l614 & ~l80;
assign a4136 = ~a4134 & ~a4132;
assign a4138 = ~a4136 & a820;
assign a4140 = ~a820 & l542;
assign a4142 = ~a4140 & ~a4138;
assign a4144 = ~l602 & l600;
assign a4146 = ~a3110 & l544;
assign a4148 = ~a4146 & ~a4144;
assign a4150 = ~a4148 & l80;
assign a4152 = l604 & ~l80;
assign a4154 = ~a4152 & ~a4150;
assign a4156 = ~a4154 & a820;
assign a4158 = ~a820 & l544;
assign a4160 = ~a4158 & ~a4156;
assign a4162 = l546 & ~i10;
assign a4164 = ~a4162 & ~l582;
assign a4166 = ~a4164 & l80;
assign a4168 = l598 & ~l80;
assign a4170 = ~a4168 & ~a4166;
assign a4172 = ~a4170 & a820;
assign a4174 = ~a820 & l546;
assign a4176 = ~a4174 & ~a4172;
assign a4178 = a816 & i18;
assign a4180 = ~a816 & l548;
assign a4182 = ~a4180 & ~a4178;
assign a4184 = ~a4182 & l80;
assign a4186 = l596 & ~l80;
assign a4188 = ~a4186 & ~a4184;
assign a4190 = ~a4188 & a884;
assign a4192 = ~a884 & l548;
assign a4194 = ~a4192 & ~a4190;
assign a4196 = ~a3402 & l80;
assign a4198 = l594 & ~l80;
assign a4200 = ~a4198 & ~a4196;
assign a4202 = ~a4200 & a820;
assign a4204 = ~a820 & l550;
assign a4206 = ~a4204 & ~a4202;
assign a4208 = ~a3396 & l82;
assign a4210 = ~l584 & ~l582;
assign a4212 = a4210 & l552;
assign a4214 = a4212 & ~a3154;
assign a4216 = ~a4214 & ~a4208;
assign a4218 = ~a4216 & l80;
assign a4220 = l592 & ~l80;
assign a4222 = ~a4220 & ~a4218;
assign a4224 = ~a4222 & a820;
assign a4226 = ~a820 & l552;
assign a4228 = ~a4226 & ~a4224;
assign a4230 = ~l556 & l554;
assign a4232 = ~a4230 & ~l578;
assign a4234 = ~a4232 & l80;
assign a4236 = l580 & ~l80;
assign a4238 = ~a4236 & ~a4234;
assign a4240 = ~a4238 & a820;
assign a4242 = ~a820 & l554;
assign a4244 = ~a4242 & ~a4240;
assign a4246 = ~a2182 & a820;
assign a4248 = ~a820 & l556;
assign a4250 = ~a4248 & ~a4246;
assign a4252 = ~l560 & l558;
assign a4254 = ~a4252 & ~l572;
assign a4256 = ~a4254 & l80;
assign a4258 = l574 & ~l80;
assign a4260 = ~a4258 & ~a4256;
assign a4262 = ~a4260 & a820;
assign a4264 = ~a820 & l558;
assign a4266 = ~a4264 & ~a4262;
assign a4268 = ~a2210 & a820;
assign a4270 = ~a820 & l560;
assign a4272 = ~a4270 & ~a4268;
assign a4274 = ~a3426 & l474;
assign a4276 = ~a4274 & a3410;
assign a4278 = ~a4276 & l80;
assign a4280 = l570 & ~l80;
assign a4282 = ~a4280 & ~a4278;
assign a4284 = ~a4282 & a820;
assign a4286 = ~a820 & l562;
assign a4288 = ~a4286 & ~a4284;
assign a4290 = a816 & i12;
assign a4292 = ~a816 & l564;
assign a4294 = ~a4292 & ~a4290;
assign a4296 = ~a4294 & l80;
assign a4298 = l568 & ~l80;
assign a4300 = ~a4298 & ~a4296;
assign a4302 = ~a4300 & a884;
assign a4304 = ~a884 & l564;
assign a4306 = ~a4304 & ~a4302;
assign a4308 = l562 & l80;
assign a4310 = a4308 & ~a3418;
assign a4312 = l576 & ~l80;
assign a4314 = ~a4312 & ~a4310;
assign a4316 = ~a4314 & a820;
assign a4318 = ~a820 & l572;
assign a4320 = ~a4318 & ~a4316;
assign a4322 = l552 & l80;
assign a4324 = a4322 & ~a4210;
assign a4326 = l586 & ~l80;
assign a4328 = ~a4326 & ~a4324;
assign a4330 = ~a4328 & a820;
assign a4332 = ~a820 & l578;
assign a4334 = ~a4332 & ~a4330;
assign a4336 = a3336 & l80;
assign a4338 = a4336 & a3350;
assign a4340 = l590 & ~l80;
assign a4342 = ~a4340 & ~a4338;
assign a4344 = ~a4342 & a820;
assign a4346 = ~a820 & l582;
assign a4348 = ~a4346 & ~a4344;
assign a4350 = l508 & l80;
assign a4352 = a4350 & ~a3760;
assign a4354 = l588 & ~l80;
assign a4356 = ~a4354 & ~a4352;
assign a4358 = ~a4356 & a820;
assign a4360 = ~a820 & l584;
assign a4362 = ~a4360 & ~a4358;
assign a4364 = l602 & l600;
assign a4366 = ~a4364 & ~l608;
assign a4368 = a4366 & ~a3782;
assign a4370 = ~a4368 & l80;
assign a4372 = l610 & ~l80;
assign a4374 = ~a4372 & ~a4370;
assign a4376 = ~a4374 & a820;
assign a4378 = ~a820 & l600;
assign a4380 = ~a4378 & ~a4376;
assign a4382 = a3780 & i20;
assign a4384 = ~a4382 & ~l602;
assign a4386 = ~a3780 & i22;
assign a4388 = ~l460 & l80;
assign a4390 = a4388 & ~a4386;
assign a4392 = a4390 & ~a4384;
assign a4394 = l606 & ~l80;
assign a4396 = ~a4394 & ~a4392;
assign a4398 = ~a4396 & a820;
assign a4400 = ~a820 & l602;
assign a4402 = ~a4400 & ~a4398;
assign a4404 = a3186 & l542;
assign a4406 = ~a3374 & l474;
assign a4408 = ~a4406 & ~a4404;
assign a4410 = ~a4408 & l80;
assign a4412 = l612 & ~l80;
assign a4414 = ~a4412 & ~a4410;
assign a4416 = ~a4414 & a820;
assign a4418 = ~a820 & l608;
assign a4420 = ~a4418 & ~a4416;
assign a4422 = ~a2394 & a820;
assign a4424 = ~a820 & l616;
assign a4426 = ~a4424 & ~a4422;
assign a4428 = ~a4098 & l618;
assign a4430 = ~a4428 & a3188;
assign a4432 = ~a4430 & l80;
assign a4434 = l684 & ~l80;
assign a4436 = ~a4434 & ~a4432;
assign a4438 = ~a4436 & a820;
assign a4440 = ~a820 & l618;
assign a4442 = ~a4440 & ~a4438;
assign a4444 = ~a2406 & a820;
assign a4446 = ~a820 & l620;
assign a4448 = ~a4446 & ~a4444;
assign a4450 = ~a2418 & a820;
assign a4452 = ~a820 & l622;
assign a4454 = ~a4452 & ~a4450;
assign a4456 = ~a2430 & a820;
assign a4458 = ~a820 & l624;
assign a4460 = ~a4458 & ~a4456;
assign a4462 = l638 & l80;
assign a4464 = l640 & ~l80;
assign a4466 = ~a4464 & ~a4462;
assign a4468 = ~a4466 & a820;
assign a4470 = ~a820 & l626;
assign a4472 = ~a4470 & ~a4468;
assign a4474 = ~a3154 & l630;
assign a4476 = a4474 & ~a3404;
assign a4478 = l628 & ~l626;
assign a4480 = ~a4478 & ~a4476;
assign a4482 = ~a4480 & l80;
assign a4484 = l636 & ~l80;
assign a4486 = ~a4484 & ~a4482;
assign a4488 = ~a4486 & a820;
assign a4490 = ~a820 & l628;
assign a4492 = ~a4490 & ~a4488;
assign a4494 = a4092 & l474;
assign a4496 = a4474 & a3404;
assign a4498 = ~a4496 & ~a4494;
assign a4500 = ~a4498 & l80;
assign a4502 = l634 & ~l80;
assign a4504 = ~a4502 & ~a4500;
assign a4506 = ~a4504 & a820;
assign a4508 = ~a820 & l630;
assign a4510 = ~a4508 & ~a4506;
assign a4512 = l642 & l80;
assign a4514 = l644 & ~l80;
assign a4516 = ~a4514 & ~a4512;
assign a4518 = ~a4516 & a820;
assign a4520 = ~a820 & l638;
assign a4522 = ~a4520 & ~a4518;
assign a4524 = l646 & l80;
assign a4526 = l648 & ~l80;
assign a4528 = ~a4526 & ~a4524;
assign a4530 = ~a4528 & a820;
assign a4532 = ~a820 & l642;
assign a4534 = ~a4532 & ~a4530;
assign a4536 = l650 & l80;
assign a4538 = l652 & ~l80;
assign a4540 = ~a4538 & ~a4536;
assign a4542 = ~a4540 & a820;
assign a4544 = ~a820 & l646;
assign a4546 = ~a4544 & ~a4542;
assign a4548 = l654 & l80;
assign a4550 = l656 & ~l80;
assign a4552 = ~a4550 & ~a4548;
assign a4554 = ~a4552 & a820;
assign a4556 = ~a820 & l650;
assign a4558 = ~a4556 & ~a4554;
assign a4560 = l658 & l80;
assign a4562 = l660 & ~l80;
assign a4564 = ~a4562 & ~a4560;
assign a4566 = ~a4564 & a820;
assign a4568 = ~a820 & l654;
assign a4570 = ~a4568 & ~a4566;
assign a4572 = l662 & l80;
assign a4574 = l664 & ~l80;
assign a4576 = ~a4574 & ~a4572;
assign a4578 = ~a4576 & a820;
assign a4580 = ~a820 & l658;
assign a4582 = ~a4580 & ~a4578;
assign a4584 = l666 & l80;
assign a4586 = l668 & ~l80;
assign a4588 = ~a4586 & ~a4584;
assign a4590 = ~a4588 & a820;
assign a4592 = ~a820 & l662;
assign a4594 = ~a4592 & ~a4590;
assign a4596 = l670 & l80;
assign a4598 = l672 & ~l80;
assign a4600 = ~a4598 & ~a4596;
assign a4602 = ~a4600 & a820;
assign a4604 = ~a820 & l666;
assign a4606 = ~a4604 & ~a4602;
assign a4608 = l674 & l80;
assign a4610 = l676 & ~l80;
assign a4612 = ~a4610 & ~a4608;
assign a4614 = ~a4612 & a820;
assign a4616 = ~a820 & l670;
assign a4618 = ~a4616 & ~a4614;
assign a4620 = l678 & l80;
assign a4622 = l680 & ~l80;
assign a4624 = ~a4622 & ~a4620;
assign a4626 = ~a4624 & a820;
assign a4628 = ~a820 & l674;
assign a4630 = ~a4628 & ~a4626;
assign a4632 = a4476 & l80;
assign a4634 = l682 & ~l80;
assign a4636 = ~a4634 & ~a4632;
assign a4638 = ~a4636 & a820;
assign a4640 = ~a820 & l678;
assign a4642 = ~a4640 & ~a4638;
assign a4644 = ~l618 & ~l540;
assign a4646 = ~a4644 & a3436;
assign a4648 = l692 & l80;
assign a4650 = a4648 & a4646;
assign a4652 = l694 & ~l80;
assign a4654 = ~a4652 & ~a4650;
assign a4656 = ~a4654 & a820;
assign a4658 = ~a820 & l688;
assign a4660 = ~a4658 & ~a4656;
assign a4662 = ~a4646 & l692;
assign a4664 = a3190 & l478;
assign a4666 = ~a3276 & l474;
assign a4668 = ~a4666 & ~a4664;
assign a4670 = a4668 & ~a4662;
assign a4672 = ~a4670 & l80;
assign a4674 = l696 & ~l80;
assign a4676 = ~a4674 & ~a4672;
assign a4678 = ~a4676 & a820;
assign a4680 = ~a820 & l692;
assign a4682 = ~a4680 & ~a4678;
assign a4684 = l714 & l620;
assign a4686 = a4684 & a4006;
assign a4688 = ~a4006 & l474;
assign a4690 = a3320 & ~l496;
assign a4692 = ~a4690 & a3324;
assign a4694 = ~a3220 & ~l496;
assign a4696 = a4694 & ~a3304;
assign a4698 = ~a4696 & a4692;
assign a4700 = ~a4698 & a4688;
assign a4702 = ~a4700 & ~a4686;
assign a4704 = ~a4006 & ~l474;
assign a4706 = a4704 & l698;
assign a4708 = ~a4706 & a4702;
assign a4710 = ~a4708 & l80;
assign a4712 = l716 & ~l80;
assign a4714 = ~a4712 & ~a4710;
assign a4716 = ~a4714 & a820;
assign a4718 = ~a820 & l698;
assign a4720 = ~a4718 & ~a4716;
assign a4722 = ~a3296 & a3294;
assign a4724 = ~a4722 & ~a3364;
assign a4726 = ~a4724 & ~a3084;
assign a4728 = a4726 & ~l496;
assign a4730 = ~a4728 & ~a3308;
assign a4732 = ~a4696 & ~a4690;
assign a4734 = a4732 & a4730;
assign a4736 = ~a4734 & a4688;
assign a4738 = a4704 & l700;
assign a4740 = ~a4738 & ~a4736;
assign a4742 = ~a4740 & l80;
assign a4744 = l712 & ~l80;
assign a4746 = ~a4744 & ~a4742;
assign a4748 = ~a4746 & a820;
assign a4750 = ~a820 & l700;
assign a4752 = ~a4750 & ~a4748;
assign a4754 = a3312 & a3096;
assign a4756 = a4754 & a4688;
assign a4758 = a4704 & l702;
assign a4760 = ~a4758 & ~a4756;
assign a4762 = ~a4760 & l80;
assign a4764 = l710 & ~l80;
assign a4766 = ~a4764 & ~a4762;
assign a4768 = ~a4766 & a820;
assign a4770 = ~a820 & l702;
assign a4772 = ~a4770 & ~a4768;
assign a4774 = ~l500 & ~l498;
assign a4776 = a4774 & a3088;
assign a4778 = ~a4776 & ~a4726;
assign a4780 = a4778 & a4692;
assign a4782 = ~a4780 & a4688;
assign a4784 = a4704 & l704;
assign a4786 = ~a4784 & ~a4782;
assign a4788 = ~a4786 & l80;
assign a4790 = l708 & ~l80;
assign a4792 = ~a4790 & ~a4788;
assign a4794 = ~a4792 & a820;
assign a4796 = ~a820 & l704;
assign a4798 = ~a4796 & ~a4794;
assign a4800 = ~a2790 & a820;
assign a4802 = ~a820 & l714;
assign a4804 = ~a4802 & ~a4800;
assign a4806 = ~a3820 & ~l512;
assign a4808 = a4806 & l736;
assign a4810 = l736 & ~l514;
assign a4812 = l748 & ~l514;
assign a4814 = l750 & ~l514;
assign a4816 = ~a4814 & ~a4812;
assign a4818 = a4816 & ~a4810;
assign a4820 = ~a4816 & a4810;
assign a4822 = ~a4820 & ~a4818;
assign a4824 = ~a4822 & ~a4806;
assign a4826 = ~a4824 & ~a4808;
assign a4828 = ~a4826 & l80;
assign a4830 = l772 & ~l80;
assign a4832 = ~a4830 & ~a4828;
assign a4834 = ~a4832 & a820;
assign a4836 = ~a820 & l736;
assign a4838 = ~a4836 & ~a4834;
assign a4840 = a4806 & l738;
assign a4842 = l752 & ~l514;
assign a4844 = ~a4842 & a4818;
assign a4846 = l738 & ~l514;
assign a4848 = ~a4846 & a4844;
assign a4850 = a4846 & ~a4844;
assign a4852 = ~a4850 & ~a4848;
assign a4854 = ~a4852 & ~a4806;
assign a4856 = ~a4854 & ~a4840;
assign a4858 = ~a4856 & l80;
assign a4860 = l770 & ~l80;
assign a4862 = ~a4860 & ~a4858;
assign a4864 = ~a4862 & a820;
assign a4866 = ~a820 & l738;
assign a4868 = ~a4866 & ~a4864;
assign a4870 = a4806 & l740;
assign a4872 = l740 & ~l514;
assign a4874 = ~a4872 & a4848;
assign a4876 = a4872 & ~a4848;
assign a4878 = ~a4876 & ~a4874;
assign a4880 = ~a4878 & ~a4806;
assign a4882 = ~a4880 & ~a4870;
assign a4884 = ~a4882 & l80;
assign a4886 = l768 & ~l80;
assign a4888 = ~a4886 & ~a4884;
assign a4890 = ~a4888 & a820;
assign a4892 = ~a820 & l740;
assign a4894 = ~a4892 & ~a4890;
assign a4896 = a4806 & l742;
assign a4898 = l742 & ~l514;
assign a4900 = ~a4898 & a4874;
assign a4902 = a4898 & ~a4874;
assign a4904 = ~a4902 & ~a4900;
assign a4906 = ~a4904 & ~a4806;
assign a4908 = ~a4906 & ~a4896;
assign a4910 = ~a4908 & l80;
assign a4912 = l766 & ~l80;
assign a4914 = ~a4912 & ~a4910;
assign a4916 = ~a4914 & a820;
assign a4918 = ~a820 & l742;
assign a4920 = ~a4918 & ~a4916;
assign a4922 = a4806 & l744;
assign a4924 = l746 & ~l514;
assign a4926 = ~a4924 & a4900;
assign a4928 = l744 & ~l514;
assign a4930 = a4928 & ~a4926;
assign a4932 = ~a4928 & a4926;
assign a4934 = ~a4932 & ~a4930;
assign a4936 = ~a4934 & ~a4806;
assign a4938 = ~a4936 & ~a4922;
assign a4940 = ~a4938 & l80;
assign a4942 = l764 & ~l80;
assign a4944 = ~a4942 & ~a4940;
assign a4946 = ~a4944 & a820;
assign a4948 = ~a820 & l744;
assign a4950 = ~a4948 & ~a4946;
assign a4952 = a4806 & l746;
assign a4954 = a4924 & ~a4900;
assign a4956 = ~a4954 & ~a4926;
assign a4958 = ~a4956 & ~a4806;
assign a4960 = ~a4958 & ~a4952;
assign a4962 = ~a4960 & l80;
assign a4964 = l762 & ~l80;
assign a4966 = ~a4964 & ~a4962;
assign a4968 = ~a4966 & a820;
assign a4970 = ~a820 & l746;
assign a4972 = ~a4970 & ~a4968;
assign a4974 = a4806 & l748;
assign a4976 = a4812 & l750;
assign a4978 = ~a4976 & ~a4816;
assign a4980 = ~a4978 & ~a4806;
assign a4982 = ~a4980 & ~a4974;
assign a4984 = ~a4982 & l80;
assign a4986 = l760 & ~l80;
assign a4988 = ~a4986 & ~a4984;
assign a4990 = ~a4988 & a820;
assign a4992 = ~a820 & l748;
assign a4994 = ~a4992 & ~a4990;
assign a4996 = a4806 & l750;
assign a4998 = ~a4814 & ~a4806;
assign a5000 = ~a4998 & ~a4996;
assign a5002 = ~a5000 & l80;
assign a5004 = l758 & ~l80;
assign a5006 = ~a5004 & ~a5002;
assign a5008 = ~a5006 & a820;
assign a5010 = ~a820 & l750;
assign a5012 = ~a5010 & ~a5008;
assign a5014 = a4806 & l752;
assign a5016 = a4842 & ~a4818;
assign a5018 = ~a5016 & ~a4844;
assign a5020 = ~a5018 & ~a4806;
assign a5022 = ~a5020 & ~a5014;
assign a5024 = ~a5022 & l80;
assign a5026 = l756 & ~l80;
assign a5028 = ~a5026 & ~a5024;
assign a5030 = ~a5028 & a820;
assign a5032 = ~a820 & l752;
assign a5034 = ~a5032 & ~a5030;
assign p0 = ~a814;

assert property (~p0);

endmodule
