module ms33 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62;

output p0;

wire na586,a598,a608,a626,a634,a644,a674,a680,a684,a692,a710,a718,a728,a752,a758,
a762,a770,a788,a796,a806,a826,a832,a836,ni62,a850,a866,a872,a1056,na1058,a1066,
a1120,a1130,a1190,a1196,a1214,a1222,a1256,a1262,a1270,a1276,a1324,a1330,a1340,a1348,a1374,
a1380,a1388,a1394,a1442,a1448,a1458,a1466,a1492,a1498,a1506,a1512,a1540,na878,na1546,na1552,
a1598,a1604,a1610,a1616,a1622,a1628,a1634,a1640,a1646,a1652,a1656,a1660,a1664,a1670,a1674,
a1684,a1698,a1700,a1702,a1710,a1714,a1724,a1738,a1742,a1752,a1766,a1778,a1784,a1788,a1818,
a1824,a1900,a1906,a1916,a1922,a1930,a1934,a1940,a1948,a1954,a1960,a1966,a1972,a1978,a1984,
a1890,a1992,a2000,a2016,a2022,a2030,a2036,a2046,a2052,a2060,a2064,a2070,a2076,a2084,a2090,
a2100,a2106,a2114,a2118,a2124,a2130,a2138,a2144,a2154,a2160,a2168,a2172,na1118,a2218,a2224,
a2230,a2236,a2242,a2248,a2254,c1,a348,a350,a352,a354,a356,a358,a360,a362,a364,
a366,a368,a370,a372,a374,a376,a378,a380,a382,a384,a386,a388,a390,a392,a394,
a396,a398,a400,a402,a404,a406,a408,a410,a412,a414,a416,a418,a420,a422,a424,
a426,a428,a430,a432,a434,a436,a438,a440,a442,a444,a446,a448,a450,a452,a454,
a456,a458,a460,a462,a464,a466,a468,a470,a472,a474,a476,a478,a480,a482,a484,
a486,a488,a490,a492,a494,a496,a498,a500,a502,a504,a506,a508,a510,a512,a514,
a516,a518,a520,a522,a524,a526,a528,a530,a532,a534,a536,a538,a540,a542,a544,
a546,a548,a550,a552,a554,a556,a558,a560,a562,a564,a566,a568,a570,a572,a574,
a576,a578,a580,a582,a584,a586,a588,a590,a592,a594,a596,a600,a602,a604,a606,
a610,a612,a614,a616,a618,a620,a622,a624,a628,a630,a632,a636,a638,a640,a642,
a646,a648,a650,a652,a654,a656,a658,a660,a662,a664,a666,a668,a670,a672,a676,
a678,a682,a686,a688,a690,a694,a696,a698,a700,a702,a704,a706,a708,a712,a714,
a716,a720,a722,a724,a726,a730,a732,a734,a736,a738,a740,a742,a744,a746,a748,
a750,a754,a756,a760,a764,a766,a768,a772,a774,a776,a778,a780,a782,a784,a786,
a790,a792,a794,a798,a800,a802,a804,a808,a810,a812,a814,a816,a818,a820,a822,
a824,a828,a830,a834,a838,a840,a842,a844,a846,a848,a852,a854,a856,a858,a860,
a862,a864,a868,a870,a874,a876,a878,a880,a882,a884,a886,a888,a890,a892,a894,
a896,a898,a900,a902,a904,a906,a908,a910,a912,a914,a916,a918,a920,a922,a924,
a926,a928,a930,a932,a934,a936,a938,a940,a942,a944,a946,a948,a950,a952,a954,
a956,a958,a960,a962,a964,a966,a968,a970,a972,a974,a976,a978,a980,a982,a984,
a986,a988,a990,a992,a994,a996,a998,a1000,a1002,a1004,a1006,a1008,a1010,a1012,a1014,
a1016,a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,a1038,a1040,a1042,a1044,
a1046,a1048,a1050,a1052,a1054,a1058,a1060,a1062,a1064,a1068,a1070,a1072,a1074,a1076,a1078,
a1080,a1082,a1084,a1086,a1088,a1090,a1092,a1094,a1096,a1098,a1100,a1102,a1104,a1106,a1108,
a1110,a1112,a1114,a1116,a1118,a1122,a1124,a1126,a1128,a1132,a1134,a1136,a1138,a1140,a1142,
a1144,a1146,a1148,a1150,a1152,a1154,a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1170,a1172,
a1174,a1176,a1178,a1180,a1182,a1184,a1186,a1188,a1192,a1194,a1198,a1200,a1202,a1204,a1206,
a1208,a1210,a1212,a1216,a1218,a1220,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,
a1242,a1244,a1246,a1248,a1250,a1252,a1254,a1258,a1260,a1264,a1266,a1268,a1272,a1274,a1278,
a1280,a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,
a1310,a1312,a1314,a1316,a1318,a1320,a1322,a1326,a1328,a1332,a1334,a1336,a1338,a1342,a1344,
a1346,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,a1368,a1370,a1372,a1376,a1378,
a1382,a1384,a1386,a1390,a1392,a1396,a1398,a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,
a1416,a1418,a1420,a1422,a1424,a1426,a1428,a1430,a1432,a1434,a1436,a1438,a1440,a1444,a1446,
a1450,a1452,a1454,a1456,a1460,a1462,a1464,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1482,
a1484,a1486,a1488,a1490,a1494,a1496,a1500,a1502,a1504,a1508,a1510,a1514,a1516,a1518,a1520,
a1522,a1524,a1526,a1528,a1530,a1532,a1534,a1536,a1538,a1542,a1544,a1546,a1548,a1550,a1552,
a1554,a1556,a1558,a1560,a1562,a1564,a1566,a1568,a1570,a1572,a1574,a1576,a1578,a1580,a1582,
a1584,a1586,a1588,a1590,a1592,a1594,a1596,a1600,a1602,a1606,a1608,a1612,a1614,a1618,a1620,
a1624,a1626,a1630,a1632,a1636,a1638,a1642,a1644,a1648,a1650,a1654,a1658,a1662,a1666,a1668,
a1672,a1676,a1678,a1680,a1682,a1686,a1688,a1690,a1692,a1694,a1696,a1704,a1706,a1708,a1712,
a1716,a1718,a1720,a1722,a1726,a1728,a1730,a1732,a1734,a1736,a1740,a1744,a1746,a1748,a1750,
a1754,a1756,a1758,a1760,a1762,a1764,a1768,a1770,a1772,a1774,a1776,a1780,a1782,a1786,a1790,
a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1820,a1822,
a1826,a1828,a1830,a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,a1848,a1850,a1852,a1854,
a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,a1882,a1884,
a1886,a1888,a1892,a1894,a1896,a1898,a1902,a1904,a1908,a1910,a1912,a1914,a1918,a1920,a1924,
a1926,a1928,a1932,a1936,a1938,a1942,a1944,a1946,a1950,a1952,a1956,a1958,a1962,a1964,a1968,
a1970,a1974,a1976,a1980,a1982,a1986,a1988,a1990,a1994,a1996,a1998,a2002,a2004,a2006,a2008,
a2010,a2012,a2014,a2018,a2020,a2024,a2026,a2028,a2032,a2034,a2038,a2040,a2042,a2044,a2048,
a2050,a2054,a2056,a2058,a2062,a2066,a2068,a2072,a2074,a2078,a2080,a2082,a2086,a2088,a2092,
a2094,a2096,a2098,a2102,a2104,a2108,a2110,a2112,a2116,a2120,a2122,a2126,a2128,a2132,a2134,
a2136,a2140,a2142,a2146,a2148,a2150,a2152,a2156,a2158,a2162,a2164,a2166,a2170,a2174,a2176,
a2178,a2180,a2182,a2184,a2186,a2188,a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,
a2208,a2210,a2212,a2214,a2216,a2220,a2222,a2226,a2228,a2232,a2234,a2238,a2240,a2244,a2246,
a2250,a2252,p0;

reg l64,l66,l68,l70,l72,l74,l76,l78,l80,l82,l84,l86,l88,l90,l92,
l94,l96,l98,l100,l102,l104,l106,l108,l110,l112,l114,l116,l118,l120,l122,
l124,l126,l128,l130,l132,l134,l136,l138,l140,l142,l144,l146,l148,l150,l152,
l154,l156,l158,l160,l162,l164,l166,l168,l170,l172,l174,l176,l178,l180,l182,
l184,l186,l188,l190,l192,l194,l196,l198,l200,l202,l204,l206,l208,l210,l212,
l214,l216,l218,l220,l222,l224,l226,l228,l230,l232,l234,l236,l238,l240,l242,
l244,l246,l248,l250,l252,l254,l256,l258,l260,l262,l264,l266,l268,l270,l272,
l274,l276,l278,l280,l282,l284,l286,l288,l290,l292,l294,l296,l298,l300,l302,
l304,l306,l308,l310,l312,l314,l316,l318,l320,l322,l324,l326,l328,l330,l332,
l334,l336,l338,l340,l342,l344,l346;

initial
begin
   l64 = 0;
   l66 = 0;
   l68 = 0;
   l70 = 0;
   l72 = 0;
   l74 = 0;
   l76 = 0;
   l78 = 0;
   l80 = 0;
   l82 = 0;
   l84 = 0;
   l86 = 0;
   l88 = 0;
   l90 = 0;
   l92 = 0;
   l94 = 0;
   l96 = 0;
   l98 = 0;
   l100 = 0;
   l102 = 0;
   l104 = 0;
   l106 = 0;
   l108 = 0;
   l110 = 0;
   l112 = 0;
   l114 = 0;
   l116 = 0;
   l118 = 0;
   l120 = 0;
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
end

always @(posedge na586)
   l64 <= na586;

always @(posedge a598)
   l66 <= a598;

always @(posedge a608)
   l68 <= a608;

always @(posedge a626)
   l70 <= a626;

always @(posedge a634)
   l72 <= a634;

always @(posedge a644)
   l74 <= a644;

always @(posedge a674)
   l76 <= a674;

always @(posedge a680)
   l78 <= a680;

always @(posedge a684)
   l80 <= a684;

always @(posedge a692)
   l82 <= a692;

always @(posedge a710)
   l84 <= a710;

always @(posedge a718)
   l86 <= a718;

always @(posedge a728)
   l88 <= a728;

always @(posedge a752)
   l90 <= a752;

always @(posedge a758)
   l92 <= a758;

always @(posedge a762)
   l94 <= a762;

always @(posedge a770)
   l96 <= a770;

always @(posedge a788)
   l98 <= a788;

always @(posedge a796)
   l100 <= a796;

always @(posedge a806)
   l102 <= a806;

always @(posedge a826)
   l104 <= a826;

always @(posedge a832)
   l106 <= a832;

always @(posedge a836)
   l108 <= a836;

always @(posedge ni62)
   l110 <= ni62;

always @(posedge a850)
   l112 <= a850;

always @(posedge a866)
   l114 <= a866;

always @(posedge a872)
   l116 <= a872;

always @(posedge a1056)
   l118 <= a1056;

always @(posedge na1058)
   l120 <= na1058;

always @(posedge a1066)
   l122 <= a1066;

always @(posedge a1120)
   l124 <= a1120;

always @(posedge a1130)
   l126 <= a1130;

always @(posedge a1190)
   l128 <= a1190;

always @(posedge a1196)
   l130 <= a1196;

always @(posedge a1214)
   l132 <= a1214;

always @(posedge a1222)
   l134 <= a1222;

always @(posedge a1256)
   l136 <= a1256;

always @(posedge a1262)
   l138 <= a1262;

always @(posedge a1270)
   l140 <= a1270;

always @(posedge a1276)
   l142 <= a1276;

always @(posedge a1324)
   l144 <= a1324;

always @(posedge a1330)
   l146 <= a1330;

always @(posedge a1340)
   l148 <= a1340;

always @(posedge a1348)
   l150 <= a1348;

always @(posedge a1374)
   l152 <= a1374;

always @(posedge a1380)
   l154 <= a1380;

always @(posedge a1388)
   l156 <= a1388;

always @(posedge a1394)
   l158 <= a1394;

always @(posedge a1442)
   l160 <= a1442;

always @(posedge a1448)
   l162 <= a1448;

always @(posedge a1458)
   l164 <= a1458;

always @(posedge a1466)
   l166 <= a1466;

always @(posedge a1492)
   l168 <= a1492;

always @(posedge a1498)
   l170 <= a1498;

always @(posedge a1506)
   l172 <= a1506;

always @(posedge a1512)
   l174 <= a1512;

always @(posedge a1540)
   l176 <= a1540;

always @(posedge na878)
   l178 <= na878;

always @(posedge na1546)
   l180 <= na1546;

always @(posedge na1552)
   l182 <= na1552;

always @(posedge a1598)
   l184 <= a1598;

always @(posedge a1604)
   l186 <= a1604;

always @(posedge a1610)
   l188 <= a1610;

always @(posedge a1616)
   l190 <= a1616;

always @(posedge a1622)
   l192 <= a1622;

always @(posedge a1628)
   l194 <= a1628;

always @(posedge a1634)
   l196 <= a1634;

always @(posedge a1640)
   l198 <= a1640;

always @(posedge a1646)
   l200 <= a1646;

always @(posedge a1652)
   l202 <= a1652;

always @(posedge a1656)
   l204 <= a1656;

always @(posedge a1660)
   l206 <= a1660;

always @(posedge a1664)
   l208 <= a1664;

always @(posedge a1670)
   l210 <= a1670;

always @(posedge a1674)
   l212 <= a1674;

always @(posedge a1684)
   l214 <= a1684;

always @(posedge a1698)
   l216 <= a1698;

always @(posedge a1700)
   l218 <= a1700;

always @(posedge l222)
   l220 <= l222;

always @(posedge a1702)
   l222 <= a1702;

always @(posedge a1710)
   l224 <= a1710;

always @(posedge a1714)
   l226 <= a1714;

always @(posedge a1724)
   l228 <= a1724;

always @(posedge a1738)
   l230 <= a1738;

always @(posedge a1742)
   l232 <= a1742;

always @(posedge a1752)
   l234 <= a1752;

always @(posedge a1766)
   l236 <= a1766;

always @(posedge a1778)
   l238 <= a1778;

always @(posedge a1784)
   l240 <= a1784;

always @(posedge a1788)
   l242 <= a1788;

always @(posedge a1818)
   l244 <= a1818;

always @(posedge a1824)
   l246 <= a1824;

always @(posedge a1900)
   l248 <= a1900;

always @(posedge a1906)
   l250 <= a1906;

always @(posedge a1916)
   l252 <= a1916;

always @(posedge a1922)
   l254 <= a1922;

always @(posedge a1930)
   l256 <= a1930;

always @(posedge a1934)
   l258 <= a1934;

always @(posedge a1940)
   l260 <= a1940;

always @(posedge a1948)
   l262 <= a1948;

always @(posedge a1954)
   l264 <= a1954;

always @(posedge a1960)
   l266 <= a1960;

always @(posedge a1966)
   l268 <= a1966;

always @(posedge a1972)
   l270 <= a1972;

always @(posedge a1978)
   l272 <= a1978;

always @(posedge a1984)
   l274 <= a1984;

always @(posedge a1890)
   l276 <= a1890;

always @(posedge a1992)
   l278 <= a1992;

always @(posedge a2000)
   l280 <= a2000;

always @(posedge a2016)
   l282 <= a2016;

always @(posedge a2022)
   l284 <= a2022;

always @(posedge a2030)
   l286 <= a2030;

always @(posedge a2036)
   l288 <= a2036;

always @(posedge a2046)
   l290 <= a2046;

always @(posedge a2052)
   l292 <= a2052;

always @(posedge a2060)
   l294 <= a2060;

always @(posedge a2064)
   l296 <= a2064;

always @(posedge a2070)
   l298 <= a2070;

always @(posedge a2076)
   l300 <= a2076;

always @(posedge a2084)
   l302 <= a2084;

always @(posedge a2090)
   l304 <= a2090;

always @(posedge a2100)
   l306 <= a2100;

always @(posedge a2106)
   l308 <= a2106;

always @(posedge a2114)
   l310 <= a2114;

always @(posedge a2118)
   l312 <= a2118;

always @(posedge a2124)
   l314 <= a2124;

always @(posedge a2130)
   l316 <= a2130;

always @(posedge a2138)
   l318 <= a2138;

always @(posedge a2144)
   l320 <= a2144;

always @(posedge a2154)
   l322 <= a2154;

always @(posedge a2160)
   l324 <= a2160;

always @(posedge a2168)
   l326 <= a2168;

always @(posedge a2172)
   l328 <= a2172;

always @(posedge na1118)
   l330 <= na1118;

always @(posedge a2218)
   l332 <= a2218;

always @(posedge a2224)
   l334 <= a2224;

always @(posedge a2230)
   l336 <= a2230;

always @(posedge a2236)
   l338 <= a2236;

always @(posedge a2242)
   l340 <= a2242;

always @(posedge a2248)
   l342 <= a2248;

always @(posedge a2254)
   l344 <= a2254;

always @(posedge c1)
   l346 <= c1;


assign na586 = ~a586;
assign a598 = ~a596 & ~a594;
assign a608 = ~a606 & ~a604;
assign a626 = ~a624 & ~a622;
assign a634 = ~a632 & ~a630;
assign a644 = ~a642 & ~a640;
assign a674 = ~a672 & ~a646;
assign a680 = ~a678 & ~a676;
assign a684 = ~a682 & ~a620;
assign a692 = ~a690 & ~a688;
assign a710 = ~a708 & ~a706;
assign a718 = ~a716 & ~a714;
assign a728 = ~a726 & ~a724;
assign a752 = ~a750 & ~a730;
assign a758 = ~a756 & ~a754;
assign a762 = ~a760 & ~a704;
assign a770 = ~a768 & ~a766;
assign a788 = ~a786 & ~a784;
assign a796 = ~a794 & ~a792;
assign a806 = ~a804 & ~a802;
assign a826 = ~a824 & ~a808;
assign a832 = ~a830 & ~a828;
assign a836 = ~a834 & ~a782;
assign ni62 = ~i62;
assign a850 = ~a848 & ~a840;
assign a866 = ~a864 & ~a858;
assign a872 = ~a870 & ~a868;
assign a1056 = ~a1054 & ~a1050;
assign na1058 = ~a1058;
assign a1066 = ~a1064 & ~a1060;
assign a1120 = ~a1118 & ~a1078;
assign a1130 = ~a1128 & ~a1122;
assign a1190 = ~a1188 & ~a1132;
assign a1196 = ~a1194 & ~a1192;
assign a1214 = ~a1212 & ~a1200;
assign a1222 = ~a1220 & ~a1218;
assign a1256 = ~a1254 & a1250;
assign a1262 = ~a1260 & ~a1258;
assign a1270 = ~a1268 & ~a1264;
assign a1276 = ~a1274 & ~a1272;
assign a1324 = ~a1322 & ~a1278;
assign a1330 = ~a1328 & ~a1326;
assign a1340 = ~a1338 & ~a1334;
assign a1348 = ~a1346 & ~a1344;
assign a1374 = ~a1372 & a1368;
assign a1380 = ~a1378 & ~a1376;
assign a1388 = ~a1386 & ~a1382;
assign a1394 = ~a1392 & ~a1390;
assign a1442 = ~a1440 & ~a1396;
assign a1448 = ~a1446 & ~a1444;
assign a1458 = ~a1456 & ~a1452;
assign a1466 = ~a1464 & ~a1462;
assign a1492 = ~a1490 & a1486;
assign a1498 = ~a1496 & ~a1494;
assign a1506 = ~a1504 & ~a1500;
assign a1512 = ~a1510 & ~a1508;
assign a1540 = ~a1538 & a1522;
assign na878 = ~a878;
assign na1546 = ~a1546;
assign na1552 = ~a1552;
assign a1598 = ~a1596 & ~a1554;
assign a1604 = ~a1602 & ~a1600;
assign a1610 = ~a1608 & ~a1606;
assign a1616 = ~a1614 & ~a1612;
assign a1622 = ~a1620 & ~a1618;
assign a1628 = ~a1626 & ~a1624;
assign a1634 = ~a1632 & ~a1630;
assign a1640 = ~a1638 & ~a1636;
assign a1646 = ~a1644 & ~a1642;
assign a1652 = ~a1650 & ~a1648;
assign a1656 = ~a1654 & ~a820;
assign a1660 = ~a1658 & ~a668;
assign a1664 = ~a1662 & ~a746;
assign a1670 = ~a1668 & ~a1118;
assign a1674 = ~a1672 & ~a750;
assign a1684 = ~a1682 & ~a1680;
assign a1698 = ~a1696 & a1694;
assign a1700 = a1666 & ~a650;
assign a1702 = a1124 & l224;
assign a1710 = ~a1708 & ~a1704;
assign a1714 = ~a1712 & ~a672;
assign a1724 = ~a1722 & ~a1720;
assign a1738 = ~a1736 & a1734;
assign a1742 = ~a1740 & ~a824;
assign a1752 = ~a1750 & ~a1748;
assign a1766 = ~a1764 & a1762;
assign a1778 = ~a1776 & a1774;
assign a1784 = a1782 & a1670;
assign a1788 = ~a1786 & a1670;
assign a1818 = ~a1816 & ~a1806;
assign a1824 = ~a1822 & ~a1820;
assign a1900 = ~a1898 & ~a574;
assign a1906 = ~a1904 & ~a1902;
assign a1916 = a1914 & a1912;
assign a1922 = ~a1920 & ~a1918;
assign a1930 = a1928 & a1914;
assign a1934 = ~a1932 & a1914;
assign a1940 = ~a1938 & ~a1936;
assign a1948 = ~a1946 & ~a1942;
assign a1954 = ~a1952 & ~a1950;
assign a1960 = ~a1958 & ~a1956;
assign a1966 = ~a1964 & ~a1962;
assign a1972 = ~a1970 & ~a1968;
assign a1978 = ~a1976 & ~a1974;
assign a1984 = ~a1982 & ~a1980;
assign a1890 = ~a1888 & ~a574;
assign a1992 = ~a1990 & ~a1988;
assign a2000 = ~a1998 & ~a1994;
assign a2016 = ~a2014 & ~a2002;
assign a2022 = ~a2020 & ~a2018;
assign a2030 = ~a2028 & ~a1434;
assign a2036 = ~a2034 & ~a2032;
assign a2046 = a2044 & a2042;
assign a2052 = ~a2050 & ~a2048;
assign a2060 = a2058 & a2044;
assign a2064 = ~a2062 & ~a1440;
assign a2070 = ~a2068 & ~a2066;
assign a2076 = ~a2074 & ~a2072;
assign a2084 = ~a2082 & ~a1316;
assign a2090 = ~a2088 & ~a2086;
assign a2100 = a2098 & a2096;
assign a2106 = ~a2104 & ~a2102;
assign a2114 = a2112 & a2098;
assign a2118 = ~a2116 & ~a1322;
assign a2124 = ~a2122 & ~a2120;
assign a2130 = ~a2128 & ~a2126;
assign a2138 = ~a2136 & ~a1182;
assign a2144 = ~a2142 & ~a2140;
assign a2154 = a2152 & a2150;
assign a2160 = ~a2158 & ~a2156;
assign a2168 = a2166 & a2152;
assign a2172 = ~a2170 & ~a1188;
assign na1118 = ~a1118;
assign a2218 = ~a2216 & ~a2174;
assign a2224 = ~a2222 & ~a2220;
assign a2230 = ~a2228 & ~a2226;
assign a2236 = ~a2234 & ~a2232;
assign a2242 = ~a2240 & ~a2238;
assign a2248 = ~a2246 & ~a2244;
assign a2254 = ~a2252 & ~a2250;
assign c1 = 1;
assign a348 = l114 & l112;
assign a350 = ~l346 & ~i14;
assign a352 = l346 & l110;
assign a354 = ~a352 & ~a350;
assign a356 = ~l346 & i10;
assign a358 = l346 & l102;
assign a360 = ~a358 & ~a356;
assign a362 = i12 & i10;
assign a364 = a362 & ~l346;
assign a366 = l346 & l98;
assign a368 = ~a366 & ~a364;
assign a370 = l346 & ~l104;
assign a372 = ~a370 & a368;
assign a374 = ~a372 & l96;
assign a376 = ~l346 & ~i10;
assign a378 = l346 & l108;
assign a380 = ~a378 & ~a376;
assign a382 = ~a380 & ~l100;
assign a384 = ~a382 & ~l96;
assign a386 = ~a384 & ~a374;
assign a388 = l346 & ~l106;
assign a390 = a388 & ~l96;
assign a392 = ~a380 & l96;
assign a394 = ~a392 & ~a390;
assign a396 = a394 & a386;
assign a398 = a388 & l96;
assign a400 = a370 & ~l96;
assign a402 = ~a400 & ~a398;
assign a404 = ~a402 & ~a396;
assign a406 = ~a404 & ~a360;
assign a408 = l100 & l96;
assign a410 = ~a368 & ~l96;
assign a412 = ~a410 & ~a408;
assign a414 = a412 & a406;
assign a416 = ~l346 & i6;
assign a418 = l346 & l88;
assign a420 = ~a418 & ~a416;
assign a422 = i8 & i6;
assign a424 = a422 & ~l346;
assign a426 = l346 & l84;
assign a428 = ~a426 & ~a424;
assign a430 = l346 & ~l90;
assign a432 = ~a430 & a428;
assign a434 = ~a432 & l82;
assign a436 = ~l346 & ~i6;
assign a438 = l346 & l94;
assign a440 = ~a438 & ~a436;
assign a442 = ~a440 & ~l86;
assign a444 = ~a442 & ~l82;
assign a446 = ~a444 & ~a434;
assign a448 = l346 & ~l92;
assign a450 = a448 & ~l82;
assign a452 = ~a440 & l82;
assign a454 = ~a452 & ~a450;
assign a456 = a454 & a446;
assign a458 = a448 & l82;
assign a460 = a430 & ~l82;
assign a462 = ~a460 & ~a458;
assign a464 = ~a462 & ~a456;
assign a466 = ~a464 & ~a420;
assign a468 = l86 & l82;
assign a470 = ~a428 & ~l82;
assign a472 = ~a470 & ~a468;
assign a474 = a472 & a466;
assign a476 = ~a474 & ~a414;
assign a478 = ~l346 & i2;
assign a480 = l346 & l74;
assign a482 = ~a480 & ~a478;
assign a484 = i4 & i2;
assign a486 = a484 & ~l346;
assign a488 = l346 & l70;
assign a490 = ~a488 & ~a486;
assign a492 = l346 & ~l76;
assign a494 = ~a492 & a490;
assign a496 = ~a494 & l68;
assign a498 = ~l346 & ~i2;
assign a500 = l346 & l80;
assign a502 = ~a500 & ~a498;
assign a504 = ~a502 & ~l72;
assign a506 = ~a504 & ~l68;
assign a508 = ~a506 & ~a496;
assign a510 = l346 & ~l78;
assign a512 = a510 & ~l68;
assign a514 = ~a502 & l68;
assign a516 = ~a514 & ~a512;
assign a518 = a516 & a508;
assign a520 = a510 & l68;
assign a522 = a492 & ~l68;
assign a524 = ~a522 & ~a520;
assign a526 = ~a524 & ~a518;
assign a528 = ~a526 & ~a482;
assign a530 = l72 & l68;
assign a532 = ~a490 & ~l68;
assign a534 = ~a532 & ~a530;
assign a536 = a534 & a528;
assign a538 = ~a536 & a476;
assign a540 = ~a538 & a354;
assign a542 = l346 & ~l64;
assign a544 = l346 & ~l66;
assign a546 = a544 & a542;
assign a548 = ~a546 & a540;
assign a550 = a548 & a348;
assign a552 = a550 & l116;
assign a554 = ~l256 & ~l254;
assign a556 = ~l258 & l254;
assign a558 = l346 & ~l250;
assign a560 = ~a558 & l252;
assign a562 = ~a560 & ~a556;
assign a564 = a562 & ~a554;
assign a566 = a558 & ~l252;
assign a568 = ~a566 & a564;
assign a570 = l346 & ~l246;
assign a572 = a570 & ~l248;
assign a574 = ~a572 & a568;
assign a576 = a574 & ~a548;
assign a578 = ~a574 & a548;
assign a580 = ~a578 & ~a576;
assign a582 = ~a580 & a542;
assign a584 = a580 & ~a542;
assign a586 = ~a584 & ~a582;
assign a588 = a578 & a542;
assign a590 = a576 & ~a542;
assign a592 = ~a590 & ~a588;
assign a594 = ~a592 & ~a544;
assign a596 = ~a590 & a544;
assign a600 = l346 & ~l210;
assign a602 = a600 & l188;
assign a604 = a602 & l68;
assign a606 = ~a602 & ~l68;
assign a610 = l346 & l228;
assign a612 = ~a610 & ~a498;
assign a614 = l346 & ~l230;
assign a616 = a614 & ~a612;
assign a618 = ~a616 & i22;
assign a620 = a618 & ~a502;
assign a622 = a620 & ~i26;
assign a624 = ~a620 & a490;
assign a628 = a618 & a502;
assign a630 = a628 & ~i26;
assign a632 = ~a628 & ~l72;
assign a636 = ~a618 & a602;
assign a638 = ~a636 & ~a482;
assign a640 = ~a638 & a612;
assign a642 = ~a618 & a482;
assign a646 = ~a620 & a492;
assign a648 = l346 & ~l226;
assign a650 = l346 & ~l126;
assign a652 = a650 & a602;
assign a654 = l346 & ~l204;
assign a656 = l346 & ~l208;
assign a658 = a656 & ~a414;
assign a660 = ~a658 & ~a654;
assign a662 = a476 & ~l206;
assign a664 = ~a662 & a660;
assign a666 = ~a664 & a536;
assign a668 = a666 & a548;
assign a670 = ~a668 & ~a652;
assign a672 = ~a670 & ~a648;
assign a676 = ~a628 & a510;
assign a678 = ~a670 & a648;
assign a682 = ~a618 & a502;
assign a686 = a600 & l190;
assign a688 = a686 & l82;
assign a690 = ~a686 & ~l82;
assign a694 = l346 & l214;
assign a696 = ~a694 & ~a436;
assign a698 = l346 & ~l216;
assign a700 = a698 & ~a696;
assign a702 = ~a700 & i18;
assign a704 = a702 & ~a440;
assign a706 = a704 & ~i28;
assign a708 = ~a704 & a428;
assign a712 = a702 & a440;
assign a714 = a712 & ~i28;
assign a716 = ~a712 & ~l86;
assign a720 = ~a702 & a686;
assign a722 = ~a720 & ~a420;
assign a724 = ~a722 & a696;
assign a726 = ~a702 & a420;
assign a730 = ~a704 & a430;
assign a732 = l346 & ~l212;
assign a734 = a686 & a650;
assign a736 = a658 & ~a536;
assign a738 = a654 & ~a536;
assign a740 = ~a738 & l206;
assign a742 = a740 & ~a736;
assign a744 = ~a742 & a474;
assign a746 = a744 & a548;
assign a748 = ~a746 & ~a734;
assign a750 = ~a748 & ~a732;
assign a754 = ~a712 & a448;
assign a756 = ~a748 & a732;
assign a760 = ~a702 & a440;
assign a764 = a600 & l186;
assign a766 = a764 & l96;
assign a768 = ~a764 & ~l96;
assign a772 = l346 & l234;
assign a774 = ~a772 & ~a376;
assign a776 = l346 & ~l236;
assign a778 = a776 & ~a774;
assign a780 = ~a778 & i24;
assign a782 = a780 & ~a380;
assign a784 = a782 & ~i30;
assign a786 = ~a782 & a368;
assign a790 = a780 & a380;
assign a792 = a790 & ~i30;
assign a794 = ~a790 & ~l100;
assign a798 = ~a780 & a764;
assign a800 = ~a798 & ~a360;
assign a802 = ~a800 & a774;
assign a804 = ~a780 & a360;
assign a808 = ~a782 & a370;
assign a810 = l346 & ~l232;
assign a812 = a764 & a650;
assign a814 = ~a740 & ~a474;
assign a816 = ~a814 & ~a656;
assign a818 = ~a816 & a414;
assign a820 = a818 & a548;
assign a822 = ~a820 & ~a812;
assign a824 = ~a822 & ~a810;
assign a828 = ~a790 & a388;
assign a830 = ~a822 & a810;
assign a834 = ~a780 & a380;
assign a838 = a548 & ~a348;
assign a840 = ~a838 & ~l112;
assign a842 = l346 & ~l122;
assign a844 = l346 & ~l120;
assign a846 = a844 & l118;
assign a848 = a846 & ~a842;
assign a852 = ~l116 & l114;
assign a854 = ~a852 & l112;
assign a856 = a854 & a838;
assign a858 = ~a856 & ~l114;
assign a860 = l346 & ~l118;
assign a862 = a860 & a844;
assign a864 = a862 & ~a842;
assign a868 = ~a550 & ~l116;
assign a870 = a846 & a842;
assign a874 = ~l346 & i16;
assign a876 = l346 & l178;
assign a878 = ~a876 & ~a874;
assign a880 = l346 & ~l174;
assign a882 = a880 & l82;
assign a884 = l346 & ~l172;
assign a886 = a884 & ~l82;
assign a888 = ~a886 & ~a882;
assign a890 = l346 & ~l168;
assign a892 = ~a890 & ~l170;
assign a894 = l346 & ~l166;
assign a896 = a894 & l82;
assign a898 = l346 & ~l164;
assign a900 = a898 & ~l82;
assign a902 = ~a900 & ~a896;
assign a904 = ~a902 & ~a892;
assign a906 = ~a904 & a888;
assign a908 = a472 & ~a462;
assign a910 = a908 & ~a906;
assign a912 = ~a472 & a354;
assign a914 = ~a912 & ~a910;
assign a916 = l346 & ~l162;
assign a918 = a916 & l82;
assign a920 = l346 & ~l160;
assign a922 = a920 & ~l82;
assign a924 = ~a922 & ~a918;
assign a926 = ~a924 & ~a914;
assign a928 = a926 & ~a420;
assign a930 = l346 & ~l158;
assign a932 = a930 & l96;
assign a934 = l346 & ~l156;
assign a936 = a934 & ~l96;
assign a938 = ~a936 & ~a932;
assign a940 = l346 & ~l152;
assign a942 = ~a940 & ~l154;
assign a944 = l346 & ~l150;
assign a946 = a944 & l96;
assign a948 = l346 & ~l148;
assign a950 = a948 & ~l96;
assign a952 = ~a950 & ~a946;
assign a954 = ~a952 & ~a942;
assign a956 = ~a954 & a938;
assign a958 = a412 & ~a402;
assign a960 = a958 & ~a956;
assign a962 = ~a412 & a354;
assign a964 = ~a962 & ~a960;
assign a966 = l346 & ~l146;
assign a968 = a966 & l96;
assign a970 = l346 & ~l144;
assign a972 = a970 & ~l96;
assign a974 = ~a972 & ~a968;
assign a976 = ~a974 & ~a964;
assign a978 = a976 & ~a360;
assign a980 = ~a978 & ~a928;
assign a982 = l346 & ~l142;
assign a984 = a982 & l68;
assign a986 = l346 & ~l140;
assign a988 = a986 & ~l68;
assign a990 = ~a988 & ~a984;
assign a992 = l346 & ~l136;
assign a994 = ~a992 & ~l138;
assign a996 = l346 & ~l134;
assign a998 = a996 & l68;
assign a1000 = l346 & ~l132;
assign a1002 = a1000 & ~l68;
assign a1004 = ~a1002 & ~a998;
assign a1006 = ~a1004 & ~a994;
assign a1008 = ~a1006 & a990;
assign a1010 = a534 & ~a524;
assign a1012 = a1010 & ~a1008;
assign a1014 = ~a534 & a354;
assign a1016 = ~a1014 & ~a1012;
assign a1018 = l346 & ~l130;
assign a1020 = a1018 & l68;
assign a1022 = l346 & l128;
assign a1024 = ~a1022 & ~a498;
assign a1026 = a1024 & ~l68;
assign a1028 = ~a1026 & ~a1020;
assign a1030 = ~a1028 & ~a1016;
assign a1032 = a1030 & ~a482;
assign a1034 = ~a1032 & a980;
assign a1036 = ~a1034 & ~l176;
assign a1038 = ~a1036 & a878;
assign a1040 = a1038 & ~l180;
assign a1042 = a1040 & ~l182;
assign a1044 = l346 & ~l124;
assign a1046 = ~a1044 & ~a650;
assign a1048 = a1046 & a1042;
assign a1050 = a1048 & a860;
assign a1052 = l346 & ~l332;
assign a1054 = a1052 & ~a1048;
assign a1058 = l346 & ~l330;
assign a1060 = a1048 & a842;
assign a1062 = l346 & ~l184;
assign a1064 = a1062 & ~a1048;
assign a1068 = l346 & ~l242;
assign a1070 = l346 & ~l240;
assign a1072 = a1070 & l238;
assign a1074 = a1072 & ~a1068;
assign a1076 = a1074 & ~a1048;
assign a1078 = ~a1076 & a1044;
assign a1080 = ~a978 & l190;
assign a1082 = ~a1080 & ~l186;
assign a1084 = l346 & ~l188;
assign a1086 = ~a1084 & a980;
assign a1088 = ~a1086 & a1082;
assign a1090 = ~a1088 & a1032;
assign a1092 = a1090 & a1010;
assign a1094 = ~a1032 & l186;
assign a1096 = ~a1094 & a1084;
assign a1098 = ~a1096 & ~a928;
assign a1100 = ~a1098 & ~l190;
assign a1102 = ~a1100 & a978;
assign a1104 = a1102 & a958;
assign a1106 = ~a1104 & ~a1092;
assign a1108 = a1080 & ~a1032;
assign a1110 = ~a1108 & a1096;
assign a1112 = ~a1110 & a928;
assign a1114 = a1112 & a908;
assign a1116 = ~a1114 & a1106;
assign a1118 = ~a1116 & a1036;
assign a1122 = ~a1076 & a650;
assign a1124 = l346 & ~l218;
assign a1126 = a1124 & l220;
assign a1128 = a1126 & l182;
assign a1132 = a1024 & ~a620;
assign a1134 = l346 & l328;
assign a1136 = ~a1134 & ~a498;
assign a1138 = ~l346 & ~i54;
assign a1140 = l346 & l324;
assign a1142 = ~a1140 & ~a1138;
assign a1144 = ~l346 & ~i50;
assign a1146 = l346 & l316;
assign a1148 = ~a1146 & ~a1144;
assign a1150 = ~l346 & ~i52;
assign a1152 = l346 & l320;
assign a1154 = ~a1152 & ~a1150;
assign a1156 = ~a1154 & ~a1148;
assign a1158 = a1156 & ~a1142;
assign a1160 = a1158 & a618;
assign a1162 = ~a1142 & l326;
assign a1164 = a1142 & ~l326;
assign a1166 = ~a1164 & ~a1162;
assign a1168 = ~a1154 & l322;
assign a1170 = a1154 & ~l322;
assign a1172 = ~a1170 & ~a1168;
assign a1174 = a1172 & a1166;
assign a1176 = ~a1148 & l318;
assign a1178 = a1148 & ~l318;
assign a1180 = ~a1178 & ~a1176;
assign a1182 = a1180 & a1174;
assign a1184 = a1182 & ~a1158;
assign a1186 = ~a1184 & ~a1160;
assign a1188 = ~a1186 & ~a1136;
assign a1192 = a1018 & ~a628;
assign a1194 = ~a1186 & a1136;
assign a1198 = ~a672 & ~a620;
assign a1200 = a1198 & a1000;
assign a1202 = l346 & ~l244;
assign a1204 = a1202 & ~l260;
assign a1206 = a1204 & a574;
assign a1208 = ~a1206 & a1202;
assign a1210 = a1208 & a668;
assign a1212 = a1210 & a672;
assign a1216 = ~a678 & ~a628;
assign a1218 = a1216 & a996;
assign a1220 = a1210 & a678;
assign a1224 = a992 & l138;
assign a1226 = ~a1224 & ~a994;
assign a1228 = l346 & ~l280;
assign a1230 = a1228 & a844;
assign a1232 = a1230 & ~a1084;
assign a1234 = l346 & ~l314;
assign a1236 = l346 & ~l262;
assign a1238 = a1236 & a574;
assign a1240 = a1238 & a1234;
assign a1242 = ~a1240 & a1232;
assign a1244 = a1242 & ~a1226;
assign a1246 = a1240 & ~a1232;
assign a1248 = a1246 & a1226;
assign a1250 = ~a1248 & ~a1244;
assign a1252 = ~a1246 & ~a1242;
assign a1254 = a1252 & a992;
assign a1258 = ~a1252 & l138;
assign a1260 = a1252 & ~l138;
assign a1264 = a1198 & a986;
assign a1266 = ~a1208 & a668;
assign a1268 = a1266 & a672;
assign a1272 = a1216 & a982;
assign a1274 = a1266 & a678;
assign a1278 = a970 & ~a782;
assign a1280 = l346 & ~l312;
assign a1282 = l346 & ~l308;
assign a1284 = l346 & ~l304;
assign a1286 = ~a1284 & l300;
assign a1288 = a1286 & ~a1282;
assign a1290 = a1288 & a780;
assign a1292 = ~a1282 & l310;
assign a1294 = a1282 & ~l310;
assign a1296 = ~a1294 & ~a1292;
assign a1298 = ~a1284 & l306;
assign a1300 = a1284 & ~l306;
assign a1302 = ~a1300 & ~a1298;
assign a1304 = a1302 & a1296;
assign a1306 = l346 & l302;
assign a1308 = ~a1306 & ~a356;
assign a1310 = ~a1308 & l300;
assign a1312 = a1308 & ~l300;
assign a1314 = ~a1312 & ~a1310;
assign a1316 = a1314 & a1304;
assign a1318 = a1316 & ~a1288;
assign a1320 = ~a1318 & ~a1290;
assign a1322 = ~a1320 & ~a1280;
assign a1326 = a966 & ~a790;
assign a1328 = ~a1320 & a1280;
assign a1332 = ~a824 & ~a782;
assign a1334 = a1332 & a948;
assign a1336 = a1208 & a820;
assign a1338 = a1336 & a824;
assign a1342 = ~a830 & ~a790;
assign a1344 = a1342 & a944;
assign a1346 = a1336 & a830;
assign a1350 = a940 & l154;
assign a1352 = ~a1350 & ~a942;
assign a1354 = a1230 & l186;
assign a1356 = l346 & ~l298;
assign a1358 = a1356 & a1238;
assign a1360 = ~a1358 & a1354;
assign a1362 = a1360 & ~a1352;
assign a1364 = a1358 & ~a1354;
assign a1366 = a1364 & a1352;
assign a1368 = ~a1366 & ~a1362;
assign a1370 = ~a1364 & ~a1360;
assign a1372 = a1370 & a940;
assign a1376 = ~a1370 & l154;
assign a1378 = a1370 & ~l154;
assign a1382 = a1332 & a934;
assign a1384 = ~a1208 & a820;
assign a1386 = a1384 & a824;
assign a1390 = a1342 & a930;
assign a1392 = a1384 & a830;
assign a1396 = a920 & ~a704;
assign a1398 = l346 & ~l296;
assign a1400 = l346 & ~l284;
assign a1402 = l346 & ~l292;
assign a1404 = ~a1402 & l288;
assign a1406 = a1404 & ~a1400;
assign a1408 = a1406 & a702;
assign a1410 = ~l290 & ~l288;
assign a1412 = l290 & l288;
assign a1414 = ~a1412 & ~a1410;
assign a1416 = ~a1402 & l294;
assign a1418 = a1402 & ~l294;
assign a1420 = ~a1418 & ~a1416;
assign a1422 = a1420 & a1414;
assign a1424 = l346 & l286;
assign a1426 = ~a1424 & ~a416;
assign a1428 = ~a1426 & ~a1400;
assign a1430 = a1426 & a1400;
assign a1432 = ~a1430 & ~a1428;
assign a1434 = a1432 & a1422;
assign a1436 = a1434 & ~a1406;
assign a1438 = ~a1436 & ~a1408;
assign a1440 = ~a1438 & ~a1398;
assign a1444 = a916 & ~a712;
assign a1446 = ~a1438 & a1398;
assign a1450 = ~a750 & ~a704;
assign a1452 = a1450 & a898;
assign a1454 = a1208 & a746;
assign a1456 = a1454 & a750;
assign a1460 = ~a756 & ~a712;
assign a1462 = a1460 & a894;
assign a1464 = a1454 & a756;
assign a1468 = a890 & l170;
assign a1470 = ~a1468 & ~a892;
assign a1472 = a1230 & l190;
assign a1474 = l346 & ~l278;
assign a1476 = a1474 & a1238;
assign a1478 = ~a1476 & a1472;
assign a1480 = a1478 & ~a1470;
assign a1482 = a1476 & ~a1472;
assign a1484 = a1482 & a1470;
assign a1486 = ~a1484 & ~a1480;
assign a1488 = ~a1482 & ~a1478;
assign a1490 = a1488 & a890;
assign a1494 = ~a1488 & l170;
assign a1496 = a1488 & ~l170;
assign a1500 = a1450 & a884;
assign a1502 = ~a1208 & a746;
assign a1504 = a1502 & a750;
assign a1508 = a1460 & a880;
assign a1510 = a1502 & a756;
assign a1514 = ~l220 & l180;
assign a1516 = a1074 & a1044;
assign a1518 = ~a1516 & ~a1514;
assign a1520 = a1034 & ~l176;
assign a1522 = ~a1520 & a1518;
assign a1524 = a1074 & a650;
assign a1526 = a978 & l190;
assign a1528 = a1032 & l186;
assign a1530 = ~a1528 & ~a1526;
assign a1532 = a1112 & ~a1084;
assign a1534 = ~a1532 & a1530;
assign a1536 = ~a1534 & ~a1116;
assign a1538 = a1536 & a1524;
assign a1542 = l220 & l180;
assign a1544 = ~a1536 & a1524;
assign a1546 = ~a1544 & ~a1542;
assign a1548 = ~a1126 & l182;
assign a1550 = a1116 & a1036;
assign a1552 = ~a1550 & ~a1548;
assign a1554 = a1062 & a1048;
assign a1556 = l346 & ~l202;
assign a1558 = a1556 & l82;
assign a1560 = l346 & ~l200;
assign a1562 = a1560 & ~l82;
assign a1564 = ~a1562 & ~a1558;
assign a1566 = ~a1564 & a1114;
assign a1568 = l346 & ~l198;
assign a1570 = a1568 & l68;
assign a1572 = l346 & ~l196;
assign a1574 = a1572 & ~l68;
assign a1576 = ~a1574 & ~a1570;
assign a1578 = ~a1576 & a1092;
assign a1580 = ~a1578 & ~a1566;
assign a1582 = l346 & ~l194;
assign a1584 = a1582 & l96;
assign a1586 = l346 & ~l192;
assign a1588 = a1586 & ~l96;
assign a1590 = ~a1588 & ~a1584;
assign a1592 = ~a1590 & a1104;
assign a1594 = ~a1592 & a1580;
assign a1596 = ~a1594 & ~a1048;
assign a1600 = ~a1102 & a1036;
assign a1602 = ~a1036 & ~l186;
assign a1606 = ~a1090 & a1036;
assign a1608 = a1084 & ~a1036;
assign a1612 = ~a1112 & a1036;
assign a1614 = ~a1036 & ~l190;
assign a1618 = a1586 & a1332;
assign a1620 = a824 & a348;
assign a1624 = a1582 & a1342;
assign a1626 = a830 & a348;
assign a1630 = a1572 & a1198;
assign a1632 = a672 & a348;
assign a1636 = a1568 & a1216;
assign a1638 = a678 & a348;
assign a1642 = a1560 & a1450;
assign a1644 = a750 & a348;
assign a1648 = a1556 & a1460;
assign a1650 = a756 & a348;
assign a1654 = a654 & ~a548;
assign a1658 = ~a548 & ~l206;
assign a1662 = a656 & ~a548;
assign a1666 = ~a1550 & ~l182;
assign a1668 = ~a1666 & a1126;
assign a1672 = a748 & a732;
assign a1676 = a702 & ~a686;
assign a1678 = ~a1676 & ~a720;
assign a1680 = ~a1678 & ~a696;
assign a1682 = a1678 & a696;
assign a1686 = ~a698 & a696;
assign a1688 = ~a1686 & ~a700;
assign a1690 = ~a1688 & a1676;
assign a1692 = a1688 & a720;
assign a1694 = ~a1692 & ~a1690;
assign a1696 = a1678 & a698;
assign a1704 = ~a1702 & l222;
assign a1706 = a1124 & i20;
assign a1708 = ~a1706 & ~l224;
assign a1712 = a670 & a648;
assign a1716 = a618 & ~a602;
assign a1718 = ~a1716 & ~a636;
assign a1720 = ~a1718 & ~a612;
assign a1722 = a1718 & a612;
assign a1726 = ~a614 & a612;
assign a1728 = ~a1726 & ~a616;
assign a1730 = ~a1728 & a1716;
assign a1732 = a1728 & a636;
assign a1734 = ~a1732 & ~a1730;
assign a1736 = a1718 & a614;
assign a1740 = a822 & a810;
assign a1744 = a780 & ~a764;
assign a1746 = ~a1744 & ~a798;
assign a1748 = ~a1746 & ~a774;
assign a1750 = a1746 & a774;
assign a1754 = ~a776 & a774;
assign a1756 = ~a1754 & ~a778;
assign a1758 = ~a1756 & a1744;
assign a1760 = a1756 & a798;
assign a1762 = ~a1760 & ~a1758;
assign a1764 = a1746 & a776;
assign a1768 = l346 & ~l238;
assign a1770 = ~a1070 & ~a1046;
assign a1772 = a1770 & ~a1768;
assign a1774 = ~a1772 & a1670;
assign a1776 = ~a1770 & a1768;
assign a1780 = a1070 & a1046;
assign a1782 = ~a1780 & ~a1770;
assign a1786 = ~a1772 & a1068;
assign a1790 = ~a1236 & a574;
assign a1792 = a544 & l64;
assign a1794 = a1792 & a1206;
assign a1796 = ~a1794 & a1202;
assign a1798 = ~a1796 & a548;
assign a1800 = a1798 & ~a1790;
assign a1802 = ~a1798 & a1790;
assign a1804 = ~a1802 & ~a1800;
assign a1806 = a1804 & a1202;
assign a1808 = ~a1202 & l260;
assign a1810 = ~a1808 & ~a1204;
assign a1812 = ~a1810 & ~a1800;
assign a1814 = a1810 & ~a1802;
assign a1816 = ~a1814 & ~a1812;
assign a1820 = ~a574 & a570;
assign a1822 = a574 & i36;
assign a1826 = ~l258 & ~l256;
assign a1828 = a1826 & ~l252;
assign a1830 = ~a1828 & ~l248;
assign a1832 = a1828 & ~l248;
assign a1834 = ~a484 & ~l346;
assign a1836 = l346 & l274;
assign a1838 = ~a1836 & ~a1834;
assign a1840 = ~a1838 & ~a616;
assign a1842 = l346 & ~l272;
assign a1844 = ~a1842 & a616;
assign a1846 = ~a1844 & ~a1840;
assign a1848 = ~a1846 & a602;
assign a1850 = ~a422 & ~l346;
assign a1852 = l346 & l270;
assign a1854 = ~a1852 & ~a1850;
assign a1856 = ~a1854 & ~a700;
assign a1858 = l346 & ~l268;
assign a1860 = ~a1858 & a700;
assign a1862 = ~a1860 & ~a1856;
assign a1864 = ~a1862 & a686;
assign a1866 = ~a1864 & ~a1848;
assign a1868 = ~a362 & ~l346;
assign a1870 = l346 & l266;
assign a1872 = ~a1870 & ~a1868;
assign a1874 = ~a1872 & ~a778;
assign a1876 = l346 & ~l264;
assign a1878 = ~a1876 & a778;
assign a1880 = ~a1878 & ~a1874;
assign a1882 = ~a1880 & a764;
assign a1884 = ~a1882 & a1866;
assign a1886 = ~a1884 & ~a1832;
assign a1888 = ~a1886 & ~l276;
assign a1892 = ~a1890 & l276;
assign a1894 = ~a1884 & a1832;
assign a1896 = ~a1894 & ~a1892;
assign a1898 = a1896 & ~a1830;
assign a1902 = ~a574 & a558;
assign a1904 = a574 & i34;
assign a1908 = l252 & l248;
assign a1910 = ~l252 & ~l248;
assign a1912 = ~a1910 & ~a1908;
assign a1914 = a1896 & ~a574;
assign a1918 = a574 & ~i32;
assign a1920 = ~a574 & ~l254;
assign a1924 = a1908 & l256;
assign a1926 = ~a1908 & ~l256;
assign a1928 = ~a1926 & ~a1924;
assign a1932 = ~a1924 & ~l258;
assign a1936 = ~a1804 & l260;
assign a1938 = a1804 & ~l260;
assign a1942 = a1236 & ~a574;
assign a1944 = a1792 & a1204;
assign a1946 = a1944 & a578;
assign a1950 = a1876 & ~a780;
assign a1952 = a1872 & a780;
assign a1956 = a1872 & ~a780;
assign a1958 = a780 & i30;
assign a1962 = a1858 & ~a702;
assign a1964 = a1854 & a702;
assign a1968 = a1854 & ~a702;
assign a1970 = a702 & i28;
assign a1974 = a1842 & ~a618;
assign a1976 = a1838 & a618;
assign a1980 = a1838 & ~a618;
assign a1982 = a618 & i26;
assign a1986 = ~a1946 & ~a1238;
assign a1988 = a1986 & a1474;
assign a1990 = a1946 & a744;
assign a1994 = a1228 & a1048;
assign a1996 = l346 & ~l282;
assign a1998 = a1996 & ~a1048;
assign a2002 = a1996 & a1048;
assign a2004 = a1092 & ~a1004;
assign a2006 = a1114 & ~a902;
assign a2008 = ~a2006 & ~a2004;
assign a2010 = a1104 & ~a952;
assign a2012 = ~a2010 & a2008;
assign a2014 = ~a2012 & ~a1048;
assign a2018 = ~a1434 & a1400;
assign a2020 = a1434 & i42;
assign a2024 = ~l294 & ~l290;
assign a2026 = ~a2024 & a1426;
assign a2028 = ~a2026 & ~a702;
assign a2032 = ~a1434 & ~l288;
assign a2034 = a1434 & i40;
assign a2038 = a1426 & ~l290;
assign a2040 = ~a1426 & l290;
assign a2042 = ~a2040 & ~a2038;
assign a2044 = ~a1434 & ~a702;
assign a2048 = ~a1434 & a1402;
assign a2050 = a1434 & i38;
assign a2054 = a2040 & l294;
assign a2056 = ~a2040 & ~l294;
assign a2058 = ~a2056 & ~a2054;
assign a2062 = a1438 & a1398;
assign a2066 = a1986 & a1356;
assign a2068 = a1946 & a818;
assign a2072 = ~a1316 & ~l300;
assign a2074 = a1316 & i48;
assign a2078 = ~l310 & ~l306;
assign a2080 = ~a2078 & a1308;
assign a2082 = ~a2080 & ~a780;
assign a2086 = ~a1316 & a1284;
assign a2088 = a1316 & i46;
assign a2092 = a1308 & ~l306;
assign a2094 = ~a1308 & l306;
assign a2096 = ~a2094 & ~a2092;
assign a2098 = ~a1316 & ~a780;
assign a2102 = ~a1316 & a1282;
assign a2104 = a1316 & i44;
assign a2108 = a2094 & l310;
assign a2110 = ~a2094 & ~l310;
assign a2112 = ~a2110 & ~a2108;
assign a2116 = a1320 & a1280;
assign a2120 = a1986 & a1234;
assign a2122 = a1946 & a666;
assign a2126 = ~a1182 & a1148;
assign a2128 = a1182 & i60;
assign a2132 = ~l326 & ~l322;
assign a2134 = ~a2132 & ~l318;
assign a2136 = ~a2134 & ~a618;
assign a2140 = ~a1182 & a1154;
assign a2142 = a1182 & i58;
assign a2146 = l322 & l318;
assign a2148 = ~l322 & ~l318;
assign a2150 = ~a2148 & ~a2146;
assign a2152 = ~a1182 & ~a618;
assign a2156 = ~a1182 & a1142;
assign a2158 = a1182 & i56;
assign a2162 = ~a2146 & ~l326;
assign a2164 = a2146 & l326;
assign a2166 = ~a2164 & ~a2162;
assign a2170 = a1186 & a1136;
assign a2174 = a1052 & a1048;
assign a2176 = l346 & ~l344;
assign a2178 = a2176 & l82;
assign a2180 = l346 & ~l342;
assign a2182 = a2180 & ~l82;
assign a2184 = ~a2182 & ~a2178;
assign a2186 = ~a2184 & a1114;
assign a2188 = l346 & ~l340;
assign a2190 = a2188 & l68;
assign a2192 = l346 & ~l338;
assign a2194 = a2192 & ~l68;
assign a2196 = ~a2194 & ~a2190;
assign a2198 = ~a2196 & a1092;
assign a2200 = ~a2198 & ~a2186;
assign a2202 = l346 & ~l336;
assign a2204 = a2202 & l96;
assign a2206 = l346 & ~l334;
assign a2208 = a2206 & ~l96;
assign a2210 = ~a2208 & ~a2204;
assign a2212 = ~a2210 & a1104;
assign a2214 = ~a2212 & a2200;
assign a2216 = ~a2214 & ~a1048;
assign a2220 = a2206 & a1332;
assign a2222 = a854 & a824;
assign a2226 = a2202 & a1342;
assign a2228 = a854 & a830;
assign a2232 = a2192 & a1198;
assign a2234 = a854 & a672;
assign a2238 = a2188 & a1216;
assign a2240 = a854 & a678;
assign a2244 = a2180 & a1450;
assign a2246 = a854 & a750;
assign a2250 = a2176 & a1460;
assign a2252 = a854 & a756;
assign p0 = a552;

assert property (~p0);

endmodule
