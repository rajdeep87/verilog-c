module m6s10 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98;

output p0;

wire a4234,c1,a4248,na776,z0,z1,z2,z3,z4,z5,na4252,a4286,a4306,a4342,a4480,
a4508,a4532,a4556,na4580,na4604,na4620,na4634,a4686,a4726,a4754,a4774,a4794,a4812,na4878,na4970,
a4976,a4982,a4988,na4992,a4996,a5016,a4224,a5024,a5032,a5040,a5048,a5052,a762,na5110,a5114,
a4390,a5066,a5060,z6,na5128,a5100,a3798,a5146,a5154,a5156,a5212,a5216,na5224,a5234,a5262,
a5206,a5302,a5312,a5328,a5282,na5288,z7,z8,z9,z10,z11,na5348,na5340,a3782,na5368,
na5360,a3752,a5078,na5240,a5376,a5398,na5466,na5476,a5392,a5386,a5478,a5490,na5430,na5492,a5496,
a5498,a5306,na5506,a5510,na5512,a5462,z12,na5568,na5578,na5584,a5594,a5602,a5606,a5612,a4404,
na5618,a5628,a5630,na5638,a5640,na5642,a402,a404,a406,a408,a410,a412,a414,a416,a418,
a420,a422,a424,a426,a428,a430,a432,a434,a436,a438,a440,a442,a444,a446,a448,
a450,a452,a454,a456,a458,a460,a462,a464,a466,a468,a470,a472,a474,a476,a478,
a480,a482,a484,a486,a488,a490,a492,a494,a496,a498,a500,a502,a504,a506,a508,
a510,a512,a514,a516,a518,a520,a522,a524,a526,a528,a530,a532,a534,a536,a538,
a540,a542,a544,a546,a548,a550,a552,a554,a556,a558,a560,a562,a564,a566,a568,
a570,a572,a574,a576,a578,a580,a582,a584,a586,a588,a590,a592,a594,a596,a598,
a600,a602,a604,a606,a608,a610,a612,a614,a616,a618,a620,a622,a624,a626,a628,
a630,a632,a634,a636,a638,a640,a642,a644,a646,a648,a650,a652,a654,a656,a658,
a660,a662,a664,a666,a668,a670,a672,a674,a676,a678,a680,a682,a684,a686,a688,
a690,a692,a694,a696,a698,a700,a702,a704,a706,a708,a710,a712,a714,a716,a718,
a720,a722,a724,a726,a728,a730,a732,a734,a736,a738,a740,a742,a744,a746,a748,
a750,a752,a754,a756,a758,a760,a764,a766,a768,a770,a772,a774,a776,a778,a780,
a782,a784,a786,a788,a790,a792,a794,a796,a798,a800,a802,a804,a806,a808,a810,
a812,a814,a816,a818,a820,a822,a824,a826,a828,a830,a832,a834,a836,a838,a840,
a842,a844,a846,a848,a850,a852,a854,a856,a858,a860,a862,a864,a866,a868,a870,
a872,a874,a876,a878,a880,a882,a884,a886,a888,a890,a892,a894,a896,a898,a900,
a902,a904,a906,a908,a910,a912,a914,a916,a918,a920,a922,a924,a926,a928,a930,
a932,a934,a936,a938,a940,a942,a944,a946,a948,a950,a952,a954,a956,a958,a960,
a962,a964,a966,a968,a970,a972,a974,a976,a978,a980,a982,a984,a986,a988,a990,
a992,a994,a996,a998,a1000,a1002,a1004,a1006,a1008,a1010,a1012,a1014,a1016,a1018,a1020,
a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,a1038,a1040,a1042,a1044,a1046,a1048,a1050,
a1052,a1054,a1056,a1058,a1060,a1062,a1064,a1066,a1068,a1070,a1072,a1074,a1076,a1078,a1080,
a1082,a1084,a1086,a1088,a1090,a1092,a1094,a1096,a1098,a1100,a1102,a1104,a1106,a1108,a1110,
a1112,a1114,a1116,a1118,a1120,a1122,a1124,a1126,a1128,a1130,a1132,a1134,a1136,a1138,a1140,
a1142,a1144,a1146,a1148,a1150,a1152,a1154,a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1170,
a1172,a1174,a1176,a1178,a1180,a1182,a1184,a1186,a1188,a1190,a1192,a1194,a1196,a1198,a1200,
a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,a1218,a1220,a1222,a1224,a1226,a1228,a1230,
a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,a1248,a1250,a1252,a1254,a1256,a1258,a1260,
a1262,a1264,a1266,a1268,a1270,a1272,a1274,a1276,a1278,a1280,a1282,a1284,a1286,a1288,a1290,
a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,a1310,a1312,a1314,a1316,a1318,a1320,
a1322,a1324,a1326,a1328,a1330,a1332,a1334,a1336,a1338,a1340,a1342,a1344,a1346,a1348,a1350,
a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,a1368,a1370,a1372,a1374,a1376,a1378,a1380,
a1382,a1384,a1386,a1388,a1390,a1392,a1394,a1396,a1398,a1400,a1402,a1404,a1406,a1408,a1410,
a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1426,a1428,a1430,a1432,a1434,a1436,a1438,a1440,
a1442,a1444,a1446,a1448,a1450,a1452,a1454,a1456,a1458,a1460,a1462,a1464,a1466,a1468,a1470,
a1472,a1474,a1476,a1478,a1480,a1482,a1484,a1486,a1488,a1490,a1492,a1494,a1496,a1498,a1500,
a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,a1518,a1520,a1522,a1524,a1526,a1528,a1530,
a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,a1548,a1550,a1552,a1554,a1556,a1558,a1560,
a1562,a1564,a1566,a1568,a1570,a1572,a1574,a1576,a1578,a1580,a1582,a1584,a1586,a1588,a1590,
a1592,a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,a1610,a1612,a1614,a1616,a1618,a1620,
a1622,a1624,a1626,a1628,a1630,a1632,a1634,a1636,a1638,a1640,a1642,a1644,a1646,a1648,a1650,
a1652,a1654,a1656,a1658,a1660,a1662,a1664,a1666,a1668,a1670,a1672,a1674,a1676,a1678,a1680,
a1682,a1684,a1686,a1688,a1690,a1692,a1694,a1696,a1698,a1700,a1702,a1704,a1706,a1708,a1710,
a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,a1732,a1734,a1736,a1738,a1740,
a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,a1758,a1760,a1762,a1764,a1766,a1768,a1770,
a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,a1790,a1792,a1794,a1796,a1798,a1800,
a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,a1822,a1824,a1826,a1828,a1830,
a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,a1848,a1850,a1852,a1854,a1856,a1858,a1860,
a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,a1882,a1884,a1886,a1888,a1890,
a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,a1910,a1912,a1914,a1916,a1918,a1920,
a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,a1938,a1940,a1942,a1944,a1946,a1948,a1950,
a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,a1972,a1974,a1976,a1978,a1980,
a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,a1998,a2000,a2002,a2004,a2006,a2008,a2010,
a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,a2030,a2032,a2034,a2036,a2038,a2040,
a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,a2058,a2060,a2062,a2064,a2066,a2068,a2070,
a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,a2090,a2092,a2094,a2096,a2098,a2100,
a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,a2120,a2122,a2124,a2126,a2128,a2130,
a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,a2152,a2154,a2156,a2158,a2160,
a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,a2178,a2180,a2182,a2184,a2186,a2188,a2190,
a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,a2208,a2210,a2212,a2214,a2216,a2218,a2220,
a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,a2238,a2240,a2242,a2244,a2246,a2248,a2250,
a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,a2268,a2270,a2272,a2274,a2276,a2278,a2280,
a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,a2298,a2300,a2302,a2304,a2306,a2308,a2310,
a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,a2328,a2330,a2332,a2334,a2336,a2338,a2340,
a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,a2358,a2360,a2362,a2364,a2366,a2368,a2370,
a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,a2388,a2390,a2392,a2394,a2396,a2398,a2400,
a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,a2420,a2422,a2424,a2426,a2428,a2430,
a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,a2448,a2450,a2452,a2454,a2456,a2458,a2460,
a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,a2478,a2480,a2482,a2484,a2486,a2488,a2490,
a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,a2508,a2510,a2512,a2514,a2516,a2518,a2520,
a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,a2540,a2542,a2544,a2546,a2548,a2550,
a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,a2572,a2574,a2576,a2578,a2580,
a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,a2602,a2604,a2606,a2608,a2610,
a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,a2630,a2632,a2634,a2636,a2638,a2640,
a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,a2662,a2664,a2666,a2668,a2670,
a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,a2692,a2694,a2696,a2698,a2700,
a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,a2718,a2720,a2722,a2724,a2726,a2728,a2730,
a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,a2752,a2754,a2756,a2758,a2760,
a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,a2782,a2784,a2786,a2788,a2790,
a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,a2810,a2812,a2814,a2816,a2818,a2820,
a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,a2840,a2842,a2844,a2846,a2848,a2850,
a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,a2870,a2872,a2874,a2876,a2878,a2880,
a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,a2900,a2902,a2904,a2906,a2908,a2910,
a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2930,a2932,a2934,a2936,a2938,a2940,
a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,a2960,a2962,a2964,a2966,a2968,a2970,
a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,a2988,a2990,a2992,a2994,a2996,a2998,a3000,
a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,a3022,a3024,a3026,a3028,a3030,
a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,a3048,a3050,a3052,a3054,a3056,a3058,a3060,
a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,a3078,a3080,a3082,a3084,a3086,a3088,a3090,
a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,a3112,a3114,a3116,a3118,a3120,
a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,a3142,a3144,a3146,a3148,a3150,
a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,a3172,a3174,a3176,a3178,a3180,
a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3200,a3202,a3204,a3206,a3208,a3210,
a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,a3228,a3230,a3232,a3234,a3236,a3238,a3240,
a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,a3262,a3264,a3266,a3268,a3270,
a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,a3288,a3290,a3292,a3294,a3296,a3298,a3300,
a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,a3324,a3326,a3328,a3330,
a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,a3354,a3356,a3358,a3360,
a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3382,a3384,a3386,a3388,a3390,
a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,a3408,a3410,a3412,a3414,a3416,a3418,a3420,
a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,a3438,a3440,a3442,a3444,a3446,a3448,a3450,
a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,a3468,a3470,a3472,a3474,a3476,a3478,a3480,
a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,a3498,a3500,a3502,a3504,a3506,a3508,a3510,
a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,a3528,a3530,a3532,a3534,a3536,a3538,a3540,
a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,a3558,a3560,a3562,a3564,a3566,a3568,a3570,
a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,a3588,a3590,a3592,a3594,a3596,a3598,a3600,
a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,a3618,a3620,a3622,a3624,a3626,a3628,a3630,
a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3648,a3650,a3652,a3654,a3656,a3658,a3660,
a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,a3678,a3680,a3682,a3684,a3686,a3688,a3690,
a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,a3712,a3714,a3716,a3718,a3720,
a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,a3738,a3740,a3742,a3744,a3746,a3748,a3750,
a3754,a3756,a3758,a3760,a3762,a3764,a3766,a3768,a3770,a3772,a3774,a3776,a3778,a3780,a3784,
a3786,a3788,a3790,a3792,a3794,a3796,a3800,a3802,a3804,a3806,a3808,a3810,a3812,a3814,a3816,
a3818,a3820,a3822,a3824,a3826,a3828,a3830,a3832,a3834,a3836,a3838,a3840,a3842,a3844,a3846,
a3848,a3850,a3852,a3854,a3856,a3858,a3860,a3862,a3864,a3866,a3868,a3870,a3872,a3874,a3876,
a3878,a3880,a3882,a3884,a3886,a3888,a3890,a3892,a3894,a3896,a3898,a3900,a3902,a3904,a3906,
a3908,a3910,a3912,a3914,a3916,a3918,a3920,a3922,a3924,a3926,a3928,a3930,a3932,a3934,a3936,
a3938,a3940,a3942,a3944,a3946,a3948,a3950,a3952,a3954,a3956,a3958,a3960,a3962,a3964,a3966,
a3968,a3970,a3972,a3974,a3976,a3978,a3980,a3982,a3984,a3986,a3988,a3990,a3992,a3994,a3996,
a3998,a4000,a4002,a4004,a4006,a4008,a4010,a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,
a4028,a4030,a4032,a4034,a4036,a4038,a4040,a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,
a4058,a4060,a4062,a4064,a4066,a4068,a4070,a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,
a4088,a4090,a4092,a4094,a4096,a4098,a4100,a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,
a4118,a4120,a4122,a4124,a4126,a4128,a4130,a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4146,
a4148,a4150,a4152,a4154,a4156,a4158,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,
a4178,a4180,a4182,a4184,a4186,a4188,a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,
a4208,a4210,a4212,a4214,a4216,a4218,a4220,a4222,a4226,a4228,a4230,a4232,a4236,a4238,a4240,
a4242,a4244,a4246,a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,
a4274,a4276,a4278,a4280,a4282,a4284,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,
a4308,a4310,a4312,a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,a4334,a4336,
a4338,a4340,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,a4368,
a4370,a4372,a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4392,a4394,a4396,a4398,a4400,
a4402,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,a4432,
a4434,a4436,a4438,a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,a4458,a4460,a4462,
a4464,a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4482,a4484,a4486,a4488,a4490,a4492,a4494,
a4496,a4498,a4500,a4502,a4504,a4506,a4510,a4512,a4514,a4516,a4518,a4520,a4522,a4524,a4526,
a4528,a4530,a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,a4554,a4558,a4560,
a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,a4578,a4580,a4582,a4584,a4586,a4588,a4590,
a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,a4612,a4614,a4616,a4618,a4620,
a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,a4642,a4644,a4646,a4648,a4650,
a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,a4672,a4674,a4676,a4678,a4680,
a4682,a4684,a4688,a4690,a4692,a4694,a4696,a4698,a4700,a4702,a4704,a4706,a4708,a4710,a4712,
a4714,a4716,a4718,a4720,a4722,a4724,a4728,a4730,a4732,a4734,a4736,a4738,a4740,a4742,a4744,
a4746,a4748,a4750,a4752,a4756,a4758,a4760,a4762,a4764,a4766,a4768,a4770,a4772,a4776,a4778,
a4780,a4782,a4784,a4786,a4788,a4790,a4792,a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,
a4814,a4816,a4818,a4820,a4822,a4824,a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,
a4844,a4846,a4848,a4850,a4852,a4854,a4856,a4858,a4860,a4862,a4864,a4866,a4868,a4870,a4872,
a4874,a4876,a4878,a4880,a4882,a4884,a4886,a4888,a4890,a4892,a4894,a4896,a4898,a4900,a4902,
a4904,a4906,a4908,a4910,a4912,a4914,a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,
a4934,a4936,a4938,a4940,a4942,a4944,a4946,a4948,a4950,a4952,a4954,a4956,a4958,a4960,a4962,
a4964,a4966,a4968,a4970,a4972,a4974,a4978,a4980,a4984,a4986,a4990,a4992,a4994,a4998,a5000,
a5002,a5004,a5006,a5008,a5010,a5012,a5014,a5018,a5020,a5022,a5026,a5028,a5030,a5034,a5036,
a5038,a5042,a5044,a5046,a5050,a5054,a5056,a5058,a5062,a5064,a5068,a5070,a5072,a5074,a5076,
a5080,a5082,a5084,a5086,a5088,a5090,a5092,a5094,a5096,a5098,a5102,a5104,a5106,a5108,a5110,
a5112,a5116,a5118,a5120,a5122,a5124,a5126,a5128,a5130,a5132,a5134,a5136,a5138,a5140,a5142,
a5144,a5148,a5150,a5152,a5158,a5160,a5162,a5164,a5166,a5168,a5170,a5172,a5174,a5176,a5178,
a5180,a5182,a5184,a5186,a5188,a5190,a5192,a5194,a5196,a5198,a5200,a5202,a5204,a5208,a5210,
a5214,a5218,a5220,a5222,a5224,a5226,a5228,a5230,a5232,a5236,a5238,a5240,a5242,a5244,a5246,
a5248,a5250,a5252,a5254,a5256,a5258,a5260,a5264,a5266,a5268,a5270,a5272,a5274,a5276,a5278,
a5280,a5284,a5286,a5288,a5290,a5292,a5294,a5296,a5298,a5300,a5304,a5308,a5310,a5314,a5316,
a5318,a5320,a5322,a5324,a5326,a5330,a5332,a5334,a5336,a5338,a5340,a5342,a5344,a5346,a5348,
a5350,a5352,a5354,a5356,a5358,a5360,a5362,a5364,a5366,a5368,a5370,a5372,a5374,a5378,a5380,
a5382,a5384,a5388,a5390,a5394,a5396,a5400,a5402,a5404,a5406,a5408,a5410,a5412,a5414,a5416,
a5418,a5420,a5422,a5424,a5426,a5428,a5430,a5432,a5434,a5436,a5438,a5440,a5442,a5444,a5446,
a5448,a5450,a5452,a5454,a5456,a5458,a5460,a5464,a5466,a5468,a5470,a5472,a5474,a5476,a5480,
a5482,a5484,a5486,a5488,a5492,a5494,a5500,a5502,a5504,a5506,a5508,a5512,a5514,a5516,a5518,
a5520,a5522,a5524,a5526,a5528,a5530,a5532,a5534,a5536,a5538,a5540,a5542,a5544,a5546,a5548,
a5550,a5552,a5554,a5556,a5558,a5560,a5562,a5564,a5566,a5568,a5570,a5572,a5574,a5576,a5578,
a5580,a5582,a5584,a5586,a5588,a5590,a5592,a5596,a5598,a5600,a5604,a5608,a5610,a5614,a5616,
a5618,a5620,a5622,a5624,a5626,a5632,a5634,a5636,a5638,a5642,a5644,a5646,a5648,a5650,p0;

reg l100,l102,l104,l106,l108,l110,l112,l114,l116,l118,l120,l122,l124,l126,l128,
l130,l132,l134,l136,l138,l140,l142,l144,l146,l148,l150,l152,l154,l156,l158,
l160,l162,l164,l166,l168,l170,l172,l174,l176,l178,l180,l182,l184,l186,l188,
l190,l192,l194,l196,l198,l200,l202,l204,l206,l208,l210,l212,l214,l216,l218,
l220,l222,l224,l226,l228,l230,l232,l234,l236,l238,l240,l242,l244,l246,l248,
l250,l252,l254,l256,l258,l260,l262,l264,l266,l268,l270,l272,l274,l276,l278,
l280,l282,l284,l286,l288,l290,l292,l294,l296,l298,l300,l302,l304,l306,l308,
l310,l312,l314,l316,l318,l320,l322,l324,l326,l328,l330,l332,l334,l336,l338,
l340,l342,l344,l346,l348,l350,l352,l354,l356,l358,l360,l362,l364,l366,l368,
l370,l372,l374,l376,l378,l380,l382,l384,l386,l388,l390,l392,l394,l396,l398,
l400;

initial
begin
   l100 = 0;
   l102 = 0;
   l104 = 0;
   l106 = 0;
   l108 = 0;
   l110 = 0;
   l112 = 0;
   l114 = 0;
   l116 = 0;
   l118 = 0;
   l120 = 0;
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
   l392 = 0;
   l394 = 0;
   l396 = 0;
   l398 = 0;
   l400 = 0;
end

always @(posedge a4234)
   l100 <= a4234;

always @(posedge c1)
   l102 <= c1;

always @(posedge a4248)
   l104 <= a4248;

always @(posedge l114)
   l106 <= l114;

always @(posedge na776)
   l108 <= na776;

always @(posedge z0)
   l110 <= z0;

always @(posedge z1)
   l112 <= z1;

always @(posedge z2)
   l114 <= z2;

always @(posedge l122)
   l116 <= l122;

always @(posedge z3)
   l118 <= z3;

always @(posedge z4)
   l120 <= z4;

always @(posedge z5)
   l122 <= z5;

always @(posedge na4252)
   l124 <= na4252;

always @(posedge a4286)
   l126 <= a4286;

always @(posedge a4306)
   l128 <= a4306;

always @(posedge a4342)
   l130 <= a4342;

always @(posedge a4480)
   l132 <= a4480;

always @(posedge a4508)
   l134 <= a4508;

always @(posedge a4532)
   l136 <= a4532;

always @(posedge a4556)
   l138 <= a4556;

always @(posedge na4580)
   l140 <= na4580;

always @(posedge na4604)
   l142 <= na4604;

always @(posedge na4620)
   l144 <= na4620;

always @(posedge na4634)
   l146 <= na4634;

always @(posedge a4686)
   l148 <= a4686;

always @(posedge a4726)
   l150 <= a4726;

always @(posedge a4754)
   l152 <= a4754;

always @(posedge a4774)
   l154 <= a4774;

always @(posedge a4794)
   l156 <= a4794;

always @(posedge a4812)
   l158 <= a4812;

always @(posedge l364)
   l160 <= l364;

always @(posedge na4878)
   l162 <= na4878;

always @(posedge na4970)
   l164 <= na4970;

always @(posedge a4976)
   l166 <= a4976;

always @(posedge a4982)
   l168 <= a4982;

always @(posedge a4988)
   l170 <= a4988;

always @(posedge l316)
   l172 <= l316;

always @(posedge l304)
   l174 <= l304;

always @(posedge na4992)
   l176 <= na4992;

always @(posedge l284)
   l178 <= l284;

always @(posedge l272)
   l180 <= l272;

always @(posedge l202)
   l182 <= l202;

always @(posedge a4996)
   l184 <= a4996;

always @(posedge a5016)
   l186 <= a5016;

always @(posedge a4224)
   l188 <= a4224;

always @(posedge a5024)
   l190 <= a5024;

always @(posedge a5032)
   l192 <= a5032;

always @(posedge a5040)
   l194 <= a5040;

always @(posedge a5048)
   l196 <= a5048;

always @(posedge a5052)
   l198 <= a5052;

always @(posedge a762)
   l200 <= a762;

always @(posedge l204)
   l202 <= l204;

always @(posedge l206)
   l204 <= l206;

always @(posedge l208)
   l206 <= l208;

always @(posedge na5110)
   l208 <= na5110;

always @(posedge a5114)
   l210 <= a5114;

always @(posedge l232)
   l212 <= l232;

always @(posedge a4390)
   l214 <= a4390;

always @(posedge a5066)
   l216 <= a5066;

always @(posedge a5060)
   l218 <= a5060;

always @(posedge z6)
   l220 <= z6;

always @(posedge na5128)
   l222 <= na5128;

always @(posedge a5100)
   l224 <= a5100;

always @(posedge a3798)
   l226 <= a3798;

always @(posedge a5146)
   l228 <= a5146;

always @(posedge a5154)
   l230 <= a5154;

always @(posedge l234)
   l232 <= l234;

always @(posedge l236)
   l234 <= l236;

always @(posedge l238)
   l236 <= l238;

always @(posedge a5156)
   l238 <= a5156;

always @(posedge a5212)
   l240 <= a5212;

always @(posedge a5216)
   l242 <= a5216;

always @(posedge na5224)
   l244 <= na5224;

always @(posedge a5234)
   l246 <= a5234;

always @(posedge a5262)
   l248 <= a5262;

always @(posedge a5206)
   l250 <= a5206;

always @(posedge a5302)
   l252 <= a5302;

always @(posedge a5312)
   l254 <= a5312;

always @(posedge a5328)
   l256 <= a5328;

always @(posedge a5282)
   l258 <= a5282;

always @(posedge na5288)
   l260 <= na5288;

always @(posedge z7)
   l262 <= z7;

always @(posedge z8)
   l264 <= z8;

always @(posedge z9)
   l266 <= z9;

always @(posedge z10)
   l268 <= z10;

always @(posedge z11)
   l270 <= z11;

always @(posedge l274)
   l272 <= l274;

always @(posedge l276)
   l274 <= l276;

always @(posedge l278)
   l276 <= l278;

always @(posedge na5348)
   l278 <= na5348;

always @(posedge na5340)
   l280 <= na5340;

always @(posedge a3782)
   l282 <= a3782;

always @(posedge l286)
   l284 <= l286;

always @(posedge l288)
   l286 <= l288;

always @(posedge l290)
   l288 <= l290;

always @(posedge na5368)
   l290 <= na5368;

always @(posedge na5360)
   l292 <= na5360;

always @(posedge a3752)
   l294 <= a3752;

always @(posedge l298)
   l296 <= l298;

always @(posedge l300)
   l298 <= l300;

always @(posedge l302)
   l300 <= l302;

always @(posedge a5078)
   l302 <= a5078;

always @(posedge l306)
   l304 <= l306;

always @(posedge l308)
   l306 <= l308;

always @(posedge l310)
   l308 <= l310;

always @(posedge l312)
   l310 <= l312;

always @(posedge l314)
   l312 <= l314;

always @(posedge na5240)
   l314 <= na5240;

always @(posedge l318)
   l316 <= l318;

always @(posedge l320)
   l318 <= l320;

always @(posedge a5376)
   l320 <= a5376;

always @(posedge a5398)
   l322 <= a5398;

always @(posedge na5466)
   l324 <= na5466;

always @(posedge l348)
   l326 <= l348;

always @(posedge na5476)
   l328 <= na5476;

always @(posedge a5392)
   l330 <= a5392;

always @(posedge a5386)
   l332 <= a5386;

always @(posedge a5478)
   l334 <= a5478;

always @(posedge a5490)
   l336 <= a5490;

always @(posedge na5430)
   l338 <= na5430;

always @(posedge na5492)
   l340 <= na5492;

always @(posedge a5496)
   l342 <= a5496;

always @(posedge a5498)
   l344 <= a5498;

always @(posedge a5306)
   l346 <= a5306;

always @(posedge na5506)
   l348 <= na5506;

always @(posedge a5510)
   l350 <= a5510;

always @(posedge l358)
   l352 <= l358;

always @(posedge na5512)
   l354 <= na5512;

always @(posedge a5462)
   l356 <= a5462;

always @(posedge z12)
   l358 <= z12;

always @(posedge na5568)
   l360 <= na5568;

always @(posedge na5578)
   l362 <= na5578;

always @(posedge l366)
   l364 <= l366;

always @(posedge l368)
   l366 <= l368;

always @(posedge l370)
   l368 <= l370;

always @(posedge l372)
   l370 <= l372;

always @(posedge l374)
   l372 <= l374;

always @(posedge l376)
   l374 <= l376;

always @(posedge na5584)
   l376 <= na5584;

always @(posedge a5594)
   l378 <= a5594;

always @(posedge a5602)
   l380 <= a5602;

always @(posedge a5606)
   l382 <= a5606;

always @(posedge a5612)
   l384 <= a5612;

always @(posedge a4404)
   l386 <= a4404;

always @(posedge l390)
   l388 <= l390;

always @(posedge na5618)
   l390 <= na5618;

always @(posedge a5628)
   l392 <= a5628;

always @(posedge a5630)
   l394 <= a5630;

always @(posedge na5638)
   l396 <= na5638;

always @(posedge a5640)
   l398 <= a5640;

always @(posedge na5642)
   l400 <= na5642;


assign a4234 = a4232 & ~a4224;
assign c1 = 1;
assign a4248 = a4246 & a4240;
assign na776 = ~a776;
assign z0 = l108;
assign z1 = l106;
assign z2 = l110;
assign z3 = l116;
assign z4 = l112;
assign z5 = l120;
assign na4252 = ~a4252;
assign a4286 = ~a4284 & ~a4254;
assign a4306 = ~a4304 & ~a4288;
assign a4342 = ~a4340 & ~a4308;
assign a4480 = ~a4478 & ~a4380;
assign a4508 = ~a4506 & ~a4486;
assign a4532 = ~a4530 & ~a4514;
assign a4556 = ~a4554 & ~a4538;
assign na4580 = ~a4580;
assign na4604 = ~a4604;
assign na4620 = ~a4620;
assign na4634 = ~a4634;
assign a4686 = a4684 & ~a4636;
assign a4726 = a4724 & ~a4688;
assign a4754 = a4752 & ~a4728;
assign a4774 = a4772 & ~a4756;
assign a4794 = a4792 & ~a4776;
assign a4812 = a4810 & ~a4796;
assign na4878 = ~a4878;
assign na4970 = ~a4970;
assign a4976 = ~a4974 & ~a4972;
assign a4982 = ~a4980 & ~a4978;
assign a4988 = ~a4986 & ~a4984;
assign na4992 = ~a4992;
assign a4996 = ~a4994 & ~l112;
assign a5016 = ~a5014 & ~a4964;
assign a4224 = ~a4222 & a4212;
assign a5024 = a5022 & ~a4234;
assign a5032 = a5030 & ~a4234;
assign a5040 = a5038 & ~a4234;
assign a5048 = a5046 & ~a4234;
assign a5052 = a5050 & ~a762;
assign a762 = ~a760 & ~a402;
assign na5110 = ~a5110;
assign a5114 = ~a5112 & ~l212;
assign a4390 = a4388 & a792;
assign a5066 = a5064 & a3808;
assign a5060 = ~a5058 & ~a5056;
assign z6 = l216;
assign na5128 = ~a5128;
assign a5100 = ~a5098 & ~a5096;
assign a3798 = ~a3796 & ~a3792;
assign a5146 = ~a5144 & ~a4234;
assign a5154 = ~a5152 & ~a4400;
assign a5156 = ~l240 & l106;
assign a5212 = ~a5210 & ~a5206;
assign a5216 = ~a5214 & a5202;
assign na5224 = ~a5224;
assign a5234 = ~a5232 & ~a5228;
assign a5262 = ~a5260 & ~a5248;
assign a5206 = ~a5204 & ~a5164;
assign a5302 = a5300 & a5282;
assign a5312 = a5310 & a5308;
assign a5328 = a5326 & a5308;
assign a5282 = ~a5280 & a5264;
assign na5288 = ~a5288;
assign z7 = l260;
assign z8 = l262;
assign z9 = l264;
assign z10 = l266;
assign z11 = l268;
assign na5348 = ~a5348;
assign na5340 = ~a5340;
assign a3782 = a3780 & ~a3764;
assign na5368 = ~a5368;
assign na5360 = ~a5360;
assign a3752 = a3750 & ~a3720;
assign a5078 = a5076 & ~a5054;
assign na5240 = ~a5240;
assign a5376 = ~a5374 & ~a5370;
assign a5398 = ~a5396 & i92;
assign na5466 = ~a5466;
assign na5476 = ~a5476;
assign a5392 = ~a5390 & ~a5388;
assign a5386 = a5384 & ~a5378;
assign a5478 = a5436 & ~a5420;
assign a5490 = ~a5488 & ~a5486;
assign na5430 = ~a5430;
assign na5492 = ~a5492;
assign a5496 = ~a5494 & ~a5456;
assign a5498 = a5456 & a5438;
assign a5306 = ~a5304 & ~a3810;
assign na5506 = ~a5506;
assign a5510 = a5508 & a5140;
assign na5512 = ~a5512;
assign a5462 = ~a5460 & ~l352;
assign z12 = l326;
assign na5568 = ~a5568;
assign na5578 = ~a5578;
assign na5584 = ~a5584;
assign a5594 = a5592 & a4240;
assign a5602 = a5600 & ~a762;
assign a5606 = a5604 & ~l384;
assign a5612 = ~a5610 & ~a5608;
assign a4404 = a4402 & a4390;
assign na5618 = ~a5618;
assign a5628 = a5626 & ~l384;
assign a5630 = ~a4404 & ~l396;
assign na5638 = ~a5638;
assign a5640 = ~a4404 & ~l400;
assign na5642 = ~a5642;
assign a402 = l102 & ~l100;
assign a404 = ~i12 & i10;
assign a406 = a404 & i8;
assign a408 = a406 & i14;
assign a410 = a408 & ~i6;
assign a412 = a410 & ~i16;
assign a414 = a408 & i6;
assign a416 = a406 & ~i14;
assign a418 = i12 & i10;
assign a420 = a418 & i6;
assign a422 = ~i12 & ~i10;
assign a424 = a422 & i8;
assign a426 = ~a424 & ~a420;
assign a428 = a426 & ~a416;
assign a430 = a428 & ~a414;
assign a432 = a430 & ~a412;
assign a434 = ~a432 & i18;
assign a436 = a404 & ~i8;
assign a438 = a436 & i20;
assign a440 = a438 & ~i14;
assign a442 = a440 & ~i6;
assign a444 = a442 & i16;
assign a446 = a422 & ~i8;
assign a448 = a446 & ~i20;
assign a450 = a448 & i22;
assign a452 = ~a450 & ~a444;
assign a454 = ~a452 & ~i18;
assign a456 = ~a454 & ~a434;
assign a458 = ~a456 & i24;
assign a460 = a410 & i16;
assign a462 = a440 & i6;
assign a464 = ~a462 & ~a460;
assign a466 = a442 & ~i16;
assign a468 = a438 & i14;
assign a470 = a446 & i20;
assign a472 = ~a470 & ~a468;
assign a474 = a472 & ~a466;
assign a476 = a474 & a464;
assign a478 = ~a476 & i18;
assign a480 = a478 & ~i24;
assign a482 = ~a480 & ~a458;
assign a484 = ~a482 & ~i26;
assign a486 = a418 & ~i6;
assign a488 = i12 & ~i10;
assign a490 = ~a488 & ~a486;
assign a492 = ~a490 & i26;
assign a494 = ~a492 & ~a484;
assign a496 = a436 & ~i20;
assign a498 = a496 & i22;
assign a500 = ~a498 & a494;
assign a502 = a448 & ~i22;
assign a504 = a502 & i28;
assign a506 = ~a504 & a500;
assign a508 = a496 & ~i22;
assign a510 = a502 & ~i28;
assign a512 = ~a510 & ~a508;
assign a514 = a512 & a506;
assign a516 = a514 & i4;
assign a518 = ~i12 & ~i8;
assign a520 = a518 & ~i20;
assign a522 = a520 & ~i22;
assign a524 = a522 & ~i28;
assign a526 = ~a524 & i10;
assign a528 = a526 & i30;
assign a530 = ~i16 & ~i14;
assign a532 = ~a530 & i6;
assign a534 = ~a532 & i14;
assign a536 = i12 & i6;
assign a538 = ~a532 & i16;
assign a540 = a534 & ~a518;
assign a542 = ~a534 & ~a520;
assign a544 = ~a542 & ~a540;
assign a546 = ~a544 & a538;
assign a548 = a534 & ~a522;
assign a550 = ~a534 & ~a524;
assign a552 = ~a550 & ~a548;
assign a554 = ~a552 & ~a538;
assign a556 = ~a554 & ~a546;
assign a558 = ~a556 & ~i6;
assign a560 = ~a558 & ~a536;
assign a562 = ~a560 & a534;
assign a564 = ~a562 & ~a524;
assign a566 = ~i36 & ~i32;
assign a568 = ~a566 & i34;
assign a570 = ~a568 & i32;
assign a572 = ~a564 & a526;
assign a574 = a560 & ~a524;
assign a576 = ~a574 & ~a558;
assign a578 = ~a576 & ~a546;
assign a580 = a578 & a572;
assign a582 = ~a580 & ~a522;
assign a584 = ~i24 & ~i18;
assign a586 = ~a584 & i26;
assign a588 = ~a586 & i24;
assign a590 = ~a586 & i18;
assign a592 = a572 & a546;
assign a594 = ~a592 & ~a518;
assign a596 = a594 & a588;
assign a598 = a564 & a526;
assign a600 = a598 & a546;
assign a602 = ~a600 & ~a520;
assign a604 = a602 & ~a588;
assign a606 = ~a604 & ~a596;
assign a608 = ~a606 & a590;
assign a610 = a588 & a582;
assign a612 = a598 & ~a546;
assign a614 = a612 & ~a576;
assign a616 = ~a614 & ~a524;
assign a618 = a616 & ~a588;
assign a620 = ~a618 & ~a610;
assign a622 = ~a620 & ~a590;
assign a624 = ~a622 & ~a608;
assign a626 = ~a624 & ~i26;
assign a628 = ~a626 & ~a492;
assign a630 = ~a628 & a588;
assign a632 = a628 & ~a616;
assign a634 = ~a632 & ~a630;
assign a636 = a512 & ~a492;
assign a638 = a636 & ~a608;
assign a640 = a638 & a634;
assign a642 = a640 & a582;
assign a644 = a642 & a570;
assign a646 = ~a568 & i36;
assign a648 = ~a646 & a644;
assign a650 = ~a634 & a608;
assign a652 = ~a650 & ~a492;
assign a654 = a652 & a594;
assign a656 = a654 & a570;
assign a658 = a652 & a602;
assign a660 = a634 & a608;
assign a662 = ~a660 & a658;
assign a664 = a662 & ~a570;
assign a666 = ~a664 & ~a656;
assign a668 = ~a666 & a646;
assign a670 = ~a668 & ~a648;
assign a672 = ~a490 & ~i26;
assign a674 = a672 & i34;
assign a676 = ~a674 & a670;
assign a678 = ~a676 & a570;
assign a680 = ~a662 & ~a654;
assign a682 = a680 & ~a642;
assign a684 = a682 & a672;
assign a686 = ~a684 & a676;
assign a688 = a662 & ~a642;
assign a690 = ~a688 & a686;
assign a692 = ~a690 & ~a678;
assign a694 = a692 & ~a564;
assign a696 = a676 & ~a642;
assign a698 = a696 & ~a680;
assign a700 = ~a698 & ~a668;
assign a702 = a700 & a546;
assign a704 = ~a702 & ~a694;
assign a706 = ~a700 & ~a546;
assign a708 = ~a706 & ~a704;
assign a710 = a682 & a676;
assign a712 = ~a710 & ~a674;
assign a714 = a712 & a576;
assign a716 = ~a714 & ~a708;
assign a718 = ~a712 & ~a576;
assign a720 = ~a718 & ~a716;
assign a722 = ~a720 & a528;
assign a724 = ~a722 & a516;
assign a726 = a512 & i38;
assign a728 = a634 & ~a564;
assign a730 = ~a608 & a546;
assign a732 = ~a730 & ~a728;
assign a734 = a608 & ~a546;
assign a736 = ~a734 & ~a732;
assign a738 = a636 & a576;
assign a740 = ~a738 & ~a736;
assign a742 = ~a636 & ~a576;
assign a744 = ~a742 & ~a740;
assign a746 = ~a744 & a528;
assign a748 = ~a746 & a726;
assign a750 = ~a748 & a724;
assign a752 = a750 & i40;
assign a754 = a748 & i42;
assign a756 = ~a754 & ~a752;
assign a758 = ~a756 & i2;
assign a760 = ~a758 & ~l102;
assign a764 = ~l104 & l102;
assign a766 = a750 & ~i40;
assign a768 = a748 & ~i42;
assign a770 = ~a768 & ~a766;
assign a772 = a770 & ~a528;
assign a774 = ~a772 & ~l102;
assign a776 = ~a774 & ~a764;
assign a778 = a776 & ~l106;
assign a780 = ~l114 & ~l112;
assign a782 = a780 & ~l110;
assign a784 = a782 & ~l108;
assign a786 = a784 & a778;
assign a788 = ~l118 & ~l116;
assign a790 = ~l122 & ~l120;
assign a792 = a790 & a788;
assign a794 = a792 & a786;
assign a796 = a794 & ~a762;
assign a798 = ~l124 & l102;
assign a800 = ~a756 & ~l102;
assign a802 = ~a800 & ~a798;
assign a804 = a802 & a796;
assign a806 = ~l130 & l102;
assign a808 = ~a518 & ~l102;
assign a810 = ~a808 & ~a806;
assign a812 = ~l148 & l102;
assign a814 = ~a712 & a692;
assign a816 = a814 & a752;
assign a818 = a754 & a492;
assign a820 = ~a818 & ~a816;
assign a822 = ~a820 & ~l102;
assign a824 = ~a822 & ~a812;
assign a826 = a824 & a810;
assign a828 = ~a824 & ~a810;
assign a830 = ~a828 & ~a826;
assign a832 = ~l126 & l102;
assign a834 = ~a522 & a518;
assign a836 = a834 & ~l102;
assign a838 = ~a836 & ~a832;
assign a840 = ~l150 & l102;
assign a842 = a752 & ~a700;
assign a844 = a754 & a608;
assign a846 = ~a844 & ~a842;
assign a848 = ~a846 & ~l102;
assign a850 = ~a848 & ~a840;
assign a852 = a850 & ~a838;
assign a854 = ~a850 & a838;
assign a856 = ~a854 & ~a852;
assign a858 = ~l128 & l102;
assign a860 = a522 & i28;
assign a862 = ~a860 & a520;
assign a864 = ~a862 & a518;
assign a866 = ~a864 & ~i12;
assign a868 = ~a866 & ~l102;
assign a870 = ~a868 & ~a858;
assign a872 = ~l152 & l102;
assign a874 = ~a700 & ~a692;
assign a876 = a712 & a700;
assign a878 = ~a876 & ~a874;
assign a880 = ~a878 & a752;
assign a882 = ~a634 & a512;
assign a884 = a882 & a754;
assign a886 = ~a884 & ~a880;
assign a888 = ~a886 & ~l102;
assign a890 = ~a888 & ~a872;
assign a892 = a890 & ~a870;
assign a894 = ~a890 & a870;
assign a896 = ~a894 & ~a892;
assign a898 = a896 & ~a802;
assign a900 = a898 & a856;
assign a902 = a900 & ~a830;
assign a904 = ~l154 & l102;
assign a906 = a770 & a528;
assign a908 = ~a564 & a546;
assign a910 = ~a908 & ~a536;
assign a912 = ~a910 & a906;
assign a914 = a814 & a766;
assign a916 = ~a914 & ~a912;
assign a918 = a768 & a492;
assign a920 = ~a918 & a916;
assign a922 = ~a920 & ~l102;
assign a924 = ~a922 & ~a904;
assign a926 = a924 & a810;
assign a928 = ~a924 & ~a810;
assign a930 = ~a928 & ~a926;
assign a932 = ~l156 & l102;
assign a934 = a564 & a546;
assign a936 = a562 & ~a546;
assign a938 = ~a936 & ~a934;
assign a940 = ~a938 & a906;
assign a942 = a766 & ~a700;
assign a944 = ~a942 & ~a940;
assign a946 = a768 & a608;
assign a948 = ~a946 & a944;
assign a950 = ~a948 & ~l102;
assign a952 = ~a950 & ~a932;
assign a954 = a952 & ~a838;
assign a956 = ~a952 & a838;
assign a958 = ~a956 & ~a954;
assign a960 = ~l158 & l102;
assign a962 = a906 & ~a562;
assign a964 = ~a878 & a766;
assign a966 = ~a964 & ~a962;
assign a968 = a882 & a768;
assign a970 = ~a968 & a966;
assign a972 = ~a970 & ~l102;
assign a974 = ~a972 & ~a960;
assign a976 = a974 & ~a870;
assign a978 = ~a974 & a870;
assign a980 = ~a978 & ~a976;
assign a982 = a980 & ~a796;
assign a984 = a982 & a958;
assign a986 = a984 & ~a930;
assign a988 = ~a986 & ~l160;
assign a990 = a988 & ~a902;
assign a992 = a870 & a838;
assign a994 = a992 & a810;
assign a996 = ~l132 & l102;
assign a998 = a750 & a720;
assign a1000 = a748 & a744;
assign a1002 = ~a1000 & ~a998;
assign a1004 = ~a1002 & a580;
assign a1006 = a1004 & ~l102;
assign a1008 = ~a1006 & ~a996;
assign a1010 = ~a1008 & a994;
assign a1012 = a838 & a810;
assign a1014 = a1012 & ~a870;
assign a1016 = ~l134 & l102;
assign a1018 = ~a1002 & a600;
assign a1020 = a1018 & ~l102;
assign a1022 = ~a1020 & ~a1016;
assign a1024 = ~a1022 & a1014;
assign a1026 = ~a838 & a810;
assign a1028 = a1026 & a870;
assign a1030 = ~l136 & l102;
assign a1032 = ~a1002 & a592;
assign a1034 = a1032 & ~l102;
assign a1036 = ~a1034 & ~a1030;
assign a1038 = ~a1036 & a1028;
assign a1040 = ~a870 & ~a838;
assign a1042 = a1040 & a810;
assign a1044 = ~l138 & l102;
assign a1046 = ~a1002 & a420;
assign a1048 = a1046 & ~l102;
assign a1050 = ~a1048 & ~a1044;
assign a1052 = ~a1050 & a1042;
assign a1054 = a992 & ~a810;
assign a1056 = a1054 & l140;
assign a1058 = ~a870 & ~a810;
assign a1060 = a1058 & a838;
assign a1062 = a1060 & l142;
assign a1064 = ~a838 & ~a810;
assign a1066 = a1064 & a870;
assign a1068 = a1066 & l144;
assign a1070 = ~a1066 & l146;
assign a1072 = ~a1070 & ~a1068;
assign a1074 = ~a1072 & ~a1060;
assign a1076 = ~a1074 & ~a1062;
assign a1078 = ~a1076 & ~a1054;
assign a1080 = ~a1078 & ~a1056;
assign a1082 = ~a1080 & ~a1042;
assign a1084 = ~a1082 & ~a1052;
assign a1086 = ~a1084 & ~a1028;
assign a1088 = ~a1086 & ~a1038;
assign a1090 = ~a1088 & ~a1014;
assign a1092 = ~a1090 & ~a1024;
assign a1094 = ~a1092 & ~a994;
assign a1096 = ~a1094 & ~a1010;
assign a1098 = a994 & l146;
assign a1100 = a1014 & ~a1008;
assign a1102 = a1028 & ~a1022;
assign a1104 = a1042 & ~a1036;
assign a1106 = a1054 & ~a1050;
assign a1108 = a1060 & l140;
assign a1110 = a1066 & l142;
assign a1112 = ~a1066 & l144;
assign a1114 = ~a1112 & ~a1110;
assign a1116 = ~a1114 & ~a1060;
assign a1118 = ~a1116 & ~a1108;
assign a1120 = ~a1118 & ~a1054;
assign a1122 = ~a1120 & ~a1106;
assign a1124 = ~a1122 & ~a1042;
assign a1126 = ~a1124 & ~a1104;
assign a1128 = ~a1126 & ~a1028;
assign a1130 = ~a1128 & ~a1102;
assign a1132 = ~a1130 & ~a1014;
assign a1134 = ~a1132 & ~a1100;
assign a1136 = ~a1134 & ~a994;
assign a1138 = ~a1136 & ~a1098;
assign a1140 = ~a1138 & ~a1096;
assign a1142 = ~a896 & ~a802;
assign a1144 = a1040 & ~a830;
assign a1146 = a870 & a856;
assign a1148 = ~a870 & ~a856;
assign a1150 = ~a1148 & ~a1146;
assign a1152 = ~a1040 & a830;
assign a1154 = ~a1152 & ~a1150;
assign a1156 = a1154 & ~a1144;
assign a1158 = a1156 & a1142;
assign a1160 = ~a980 & ~a796;
assign a1162 = a1040 & ~a930;
assign a1164 = a958 & a870;
assign a1166 = ~a958 & ~a870;
assign a1168 = ~a1166 & ~a1164;
assign a1170 = ~a1040 & a930;
assign a1172 = ~a1170 & ~a1168;
assign a1174 = a1172 & ~a1162;
assign a1176 = a1174 & a1160;
assign a1178 = ~a1176 & ~a1158;
assign a1180 = a1178 & ~a1140;
assign a1182 = a1180 & a990;
assign a1184 = a1138 & a1096;
assign a1186 = ~a1022 & a994;
assign a1188 = ~a1036 & a1014;
assign a1190 = ~a1050 & a1028;
assign a1192 = a1042 & l140;
assign a1194 = a1054 & l142;
assign a1196 = a1060 & l144;
assign a1198 = a1066 & l146;
assign a1200 = ~a1066 & ~a1008;
assign a1202 = ~a1200 & ~a1198;
assign a1204 = ~a1202 & ~a1060;
assign a1206 = ~a1204 & ~a1196;
assign a1208 = ~a1206 & ~a1054;
assign a1210 = ~a1208 & ~a1194;
assign a1212 = ~a1210 & ~a1042;
assign a1214 = ~a1212 & ~a1192;
assign a1216 = ~a1214 & ~a1028;
assign a1218 = ~a1216 & ~a1190;
assign a1220 = ~a1218 & ~a1014;
assign a1222 = ~a1220 & ~a1188;
assign a1224 = ~a1222 & ~a994;
assign a1226 = ~a1224 & ~a1186;
assign a1228 = ~a1226 & ~a1184;
assign a1230 = ~a1064 & ~a1012;
assign a1232 = a1230 & a824;
assign a1234 = ~a1230 & ~a824;
assign a1236 = ~a1234 & ~a856;
assign a1238 = a1236 & ~a1232;
assign a1240 = a1238 & a898;
assign a1242 = a1230 & a924;
assign a1244 = ~a1230 & ~a924;
assign a1246 = ~a1244 & ~a958;
assign a1248 = a1246 & ~a1242;
assign a1250 = a1248 & a982;
assign a1252 = ~a1250 & ~a1240;
assign a1254 = a1252 & ~a1228;
assign a1256 = a1254 & a1182;
assign a1258 = a1226 & a1184;
assign a1260 = ~a1036 & a994;
assign a1262 = ~a1050 & a1014;
assign a1264 = a1028 & l140;
assign a1266 = a1042 & l142;
assign a1268 = a1054 & l144;
assign a1270 = a1060 & l146;
assign a1272 = a1066 & ~a1008;
assign a1274 = ~a1066 & ~a1022;
assign a1276 = ~a1274 & ~a1272;
assign a1278 = ~a1276 & ~a1060;
assign a1280 = ~a1278 & ~a1270;
assign a1282 = ~a1280 & ~a1054;
assign a1284 = ~a1282 & ~a1268;
assign a1286 = ~a1284 & ~a1042;
assign a1288 = ~a1286 & ~a1266;
assign a1290 = ~a1288 & ~a1028;
assign a1292 = ~a1290 & ~a1264;
assign a1294 = ~a1292 & ~a1014;
assign a1296 = ~a1294 & ~a1262;
assign a1298 = ~a1296 & ~a994;
assign a1300 = ~a1298 & ~a1260;
assign a1302 = ~a1300 & ~a1258;
assign a1304 = ~a992 & ~a810;
assign a1306 = ~a1304 & ~a994;
assign a1308 = a1306 & a824;
assign a1310 = ~a1306 & ~a824;
assign a1312 = ~a1310 & ~a1308;
assign a1314 = a1312 & a1150;
assign a1316 = a1314 & a1142;
assign a1318 = a1306 & a924;
assign a1320 = ~a1306 & ~a924;
assign a1322 = ~a1320 & ~a1318;
assign a1324 = a1322 & a1168;
assign a1326 = a1324 & a1160;
assign a1328 = ~a1326 & ~a1316;
assign a1330 = a1328 & ~a1302;
assign a1332 = a1330 & a1256;
assign a1334 = ~a1050 & a994;
assign a1336 = a1014 & l140;
assign a1338 = a1028 & l142;
assign a1340 = a1042 & l144;
assign a1342 = a1054 & l146;
assign a1344 = a1060 & ~a1008;
assign a1346 = a1066 & ~a1022;
assign a1348 = ~a1066 & ~a1036;
assign a1350 = ~a1348 & ~a1346;
assign a1352 = ~a1350 & ~a1060;
assign a1354 = ~a1352 & ~a1344;
assign a1356 = ~a1354 & ~a1054;
assign a1358 = ~a1356 & ~a1342;
assign a1360 = ~a1358 & ~a1042;
assign a1362 = ~a1360 & ~a1340;
assign a1364 = ~a1362 & ~a1028;
assign a1366 = ~a1364 & ~a1338;
assign a1368 = ~a1366 & ~a1014;
assign a1370 = ~a1368 & ~a1336;
assign a1372 = ~a1370 & ~a994;
assign a1374 = ~a1372 & ~a1334;
assign a1376 = a1300 & a1258;
assign a1378 = ~a1376 & ~a1374;
assign a1380 = a900 & a830;
assign a1382 = a984 & a930;
assign a1384 = ~a1382 & ~a1380;
assign a1386 = a1384 & ~a1378;
assign a1388 = a1386 & a1332;
assign a1390 = a1388 & i50;
assign a1392 = ~a1390 & ~i48;
assign a1394 = ~a1392 & a1332;
assign a1396 = ~a1394 & ~i46;
assign a1398 = ~a1396 & a1256;
assign a1400 = ~a1398 & ~i44;
assign a1402 = ~a1400 & a1182;
assign a1404 = ~a1402 & ~i52;
assign a1406 = ~a1404 & a990;
assign a1408 = a802 & ~a796;
assign a1410 = a1408 & ~a810;
assign a1412 = ~a802 & ~a796;
assign a1414 = a1412 & ~a850;
assign a1416 = a1414 & ~a810;
assign a1418 = a1416 & a824;
assign a1420 = ~a1418 & ~a1410;
assign a1422 = ~a1420 & a838;
assign a1424 = a1422 & ~a924;
assign a1426 = a1424 & a952;
assign a1428 = a1412 & a850;
assign a1430 = a1428 & ~a810;
assign a1432 = a1430 & ~a824;
assign a1434 = a1432 & a838;
assign a1436 = a1434 & ~a924;
assign a1438 = a1436 & a952;
assign a1440 = a1438 & a890;
assign a1442 = ~a1440 & ~a1426;
assign a1444 = ~a1442 & a974;
assign a1446 = a1434 & a924;
assign a1448 = a1446 & ~a952;
assign a1450 = ~a802 & a796;
assign a1452 = a1450 & a850;
assign a1454 = a1452 & ~a810;
assign a1456 = a1454 & ~a824;
assign a1458 = a1456 & a838;
assign a1460 = ~a1458 & ~a1448;
assign a1462 = ~a1460 & a890;
assign a1464 = a1422 & a924;
assign a1466 = a1464 & ~a952;
assign a1468 = ~a810 & a804;
assign a1470 = a1450 & ~a850;
assign a1472 = a1470 & ~a810;
assign a1474 = a1472 & a824;
assign a1476 = ~a1474 & ~a1468;
assign a1478 = ~a1476 & a838;
assign a1480 = ~a1478 & ~a1466;
assign a1482 = a1480 & ~a1462;
assign a1484 = a1482 & ~a1444;
assign a1486 = ~a1484 & ~a870;
assign a1488 = a1486 & ~i50;
assign a1490 = a1430 & a824;
assign a1492 = a1490 & a838;
assign a1494 = a1492 & ~a924;
assign a1496 = a1494 & a952;
assign a1498 = a1496 & ~a890;
assign a1500 = a1498 & a974;
assign a1502 = a1446 & a952;
assign a1504 = a1502 & a890;
assign a1506 = a1504 & ~a974;
assign a1508 = ~a1506 & ~a1500;
assign a1510 = a1464 & a952;
assign a1512 = a1492 & a924;
assign a1514 = a1512 & a952;
assign a1516 = a1514 & ~a890;
assign a1518 = ~a1516 & ~a1510;
assign a1520 = ~a1518 & ~a974;
assign a1522 = a1512 & ~a952;
assign a1524 = a1454 & a824;
assign a1526 = a1524 & a838;
assign a1528 = ~a1526 & ~a1522;
assign a1530 = ~a1528 & ~a890;
assign a1532 = ~a1530 & ~a1520;
assign a1534 = a1532 & a1508;
assign a1536 = ~a1534 & ~a870;
assign a1538 = ~a1536 & ~a1488;
assign a1540 = ~a1538 & l146;
assign a1542 = a1486 & i50;
assign a1544 = a1542 & l146;
assign a1546 = a1544 & ~a1008;
assign a1548 = ~a1546 & ~a1540;
assign a1550 = a1544 & a1008;
assign a1552 = ~a1518 & a974;
assign a1554 = a1528 & ~a1514;
assign a1556 = ~a1554 & a890;
assign a1558 = ~a1556 & ~a1552;
assign a1560 = a1496 & a890;
assign a1562 = ~a1560 & ~a1504;
assign a1564 = ~a1562 & a974;
assign a1566 = ~a1564 & a1558;
assign a1568 = ~a1566 & ~a870;
assign a1570 = ~a1568 & ~a1550;
assign a1572 = a1570 & a1548;
assign a1574 = ~a1572 & ~l142;
assign a1576 = a1574 & l144;
assign a1578 = ~a1558 & a870;
assign a1580 = a1532 & a1480;
assign a1582 = ~a1580 & a870;
assign a1584 = a1582 & ~i50;
assign a1586 = ~a1584 & ~a1578;
assign a1588 = ~a1586 & a1050;
assign a1590 = a1582 & i50;
assign a1592 = a1590 & l146;
assign a1594 = a1592 & a1050;
assign a1596 = ~a1594 & ~a1588;
assign a1598 = ~a1596 & l142;
assign a1600 = a1590 & ~l146;
assign a1602 = a1600 & a1050;
assign a1604 = a1602 & l142;
assign a1606 = ~a1604 & ~a1598;
assign a1608 = ~a1606 & l144;
assign a1610 = ~a1494 & ~a1424;
assign a1612 = ~a1610 & ~a952;
assign a1614 = a1416 & ~a824;
assign a1616 = a1614 & a838;
assign a1618 = a1616 & ~a924;
assign a1620 = a1618 & ~a952;
assign a1622 = a1620 & ~a890;
assign a1624 = ~a1622 & ~a1612;
assign a1626 = ~a1624 & ~a974;
assign a1628 = a1616 & a924;
assign a1630 = a1472 & ~a824;
assign a1632 = a1630 & a838;
assign a1634 = ~a1632 & ~a1628;
assign a1636 = ~a1634 & ~a890;
assign a1638 = ~a1636 & ~a1626;
assign a1640 = ~a1638 & a870;
assign a1642 = a1640 & a1050;
assign a1644 = a1642 & l142;
assign a1646 = ~a1644 & ~a1608;
assign a1648 = a1646 & ~a1576;
assign a1650 = ~a1648 & ~l140;
assign a1652 = ~a1432 & ~a1410;
assign a1654 = ~a1652 & ~a838;
assign a1656 = a1654 & ~a924;
assign a1658 = a1656 & ~a952;
assign a1660 = a1614 & ~a838;
assign a1662 = a1660 & ~a924;
assign a1664 = a1662 & ~a952;
assign a1666 = a1664 & a890;
assign a1668 = ~a1666 & ~a1658;
assign a1670 = ~a1668 & a974;
assign a1672 = a1662 & a952;
assign a1674 = a1630 & ~a838;
assign a1676 = ~a1674 & ~a1672;
assign a1678 = ~a1676 & a890;
assign a1680 = a1656 & a952;
assign a1682 = ~a1468 & ~a1456;
assign a1684 = ~a1682 & ~a838;
assign a1686 = ~a1684 & ~a1680;
assign a1688 = a1686 & ~a1678;
assign a1690 = a1688 & ~a1670;
assign a1692 = ~a1690 & ~a870;
assign a1694 = a1692 & ~i50;
assign a1696 = a1418 & ~a838;
assign a1698 = a1696 & ~a924;
assign a1700 = a1698 & ~a952;
assign a1702 = a1700 & ~a890;
assign a1704 = a1702 & a974;
assign a1706 = a1660 & a924;
assign a1708 = a1706 & ~a952;
assign a1710 = a1708 & a890;
assign a1712 = a1710 & ~a974;
assign a1714 = ~a1712 & ~a1704;
assign a1716 = a1654 & a924;
assign a1718 = a1716 & ~a952;
assign a1720 = a1696 & a924;
assign a1722 = a1720 & ~a952;
assign a1724 = a1722 & ~a890;
assign a1726 = ~a1724 & ~a1718;
assign a1728 = ~a1726 & ~a974;
assign a1730 = a1698 & a952;
assign a1732 = a1474 & ~a838;
assign a1734 = ~a1732 & ~a1730;
assign a1736 = ~a1734 & ~a890;
assign a1738 = ~a1736 & ~a1728;
assign a1740 = a1738 & a1714;
assign a1742 = ~a1740 & ~a870;
assign a1744 = ~a1742 & ~a1694;
assign a1746 = ~a1744 & ~l146;
assign a1748 = a1746 & ~a1008;
assign a1750 = a1692 & i50;
assign a1752 = a1750 & ~l146;
assign a1754 = a1752 & ~a1008;
assign a1756 = a1754 & ~a1036;
assign a1758 = ~a1756 & ~a1748;
assign a1760 = ~a1758 & ~l144;
assign a1762 = a1408 & a810;
assign a1764 = a1414 & a810;
assign a1766 = a1764 & ~a824;
assign a1768 = ~a1766 & ~a1762;
assign a1770 = ~a1768 & a838;
assign a1772 = a1770 & a924;
assign a1774 = a1428 & a810;
assign a1776 = a1774 & ~a824;
assign a1778 = a1776 & a838;
assign a1780 = a1778 & a924;
assign a1782 = ~a1780 & ~a1772;
assign a1784 = ~a1782 & ~a952;
assign a1786 = a1764 & a824;
assign a1788 = a1786 & a838;
assign a1790 = a1788 & a924;
assign a1792 = a1790 & ~a952;
assign a1794 = a1792 & ~a890;
assign a1796 = ~a1794 & ~a1784;
assign a1798 = ~a1796 & ~a974;
assign a1800 = a1788 & ~a924;
assign a1802 = a1470 & a810;
assign a1804 = a1802 & a824;
assign a1806 = a1804 & a838;
assign a1808 = ~a1806 & ~a1800;
assign a1810 = ~a1808 & ~a890;
assign a1812 = ~a1810 & ~a1798;
assign a1814 = ~a1812 & a870;
assign a1816 = a1814 & ~l146;
assign a1818 = a1816 & a1008;
assign a1820 = ~a1818 & ~a1760;
assign a1822 = a1770 & ~a924;
assign a1824 = a1822 & ~a952;
assign a1826 = a810 & a804;
assign a1828 = a1802 & ~a824;
assign a1830 = ~a1828 & ~a1826;
assign a1832 = ~a1830 & a838;
assign a1834 = ~a1832 & ~a1824;
assign a1836 = a1822 & a952;
assign a1838 = a1778 & ~a924;
assign a1840 = a1838 & a952;
assign a1842 = a1840 & ~a890;
assign a1844 = ~a1842 & ~a1836;
assign a1846 = ~a1844 & ~a974;
assign a1848 = a1838 & ~a952;
assign a1850 = a1452 & a810;
assign a1852 = a1850 & ~a824;
assign a1854 = a1852 & a838;
assign a1856 = ~a1854 & ~a1848;
assign a1858 = ~a1856 & ~a890;
assign a1860 = ~a1858 & ~a1846;
assign a1862 = a1860 & a1834;
assign a1864 = ~a1862 & a870;
assign a1866 = a1864 & i50;
assign a1868 = a1866 & ~l146;
assign a1870 = a1868 & a1008;
assign a1872 = a1870 & ~a1036;
assign a1874 = a1872 & a1050;
assign a1876 = a1754 & a1036;
assign a1878 = a1876 & ~l144;
assign a1880 = ~a1878 & ~a1874;
assign a1882 = ~a1844 & a974;
assign a1884 = a1856 & ~a1840;
assign a1886 = ~a1884 & a890;
assign a1888 = ~a1886 & ~a1882;
assign a1890 = ~a1888 & a870;
assign a1892 = a1864 & ~i50;
assign a1894 = ~a1892 & ~a1890;
assign a1896 = ~a1894 & ~l146;
assign a1898 = a1896 & a1008;
assign a1900 = a1898 & ~a1036;
assign a1902 = a1872 & ~a1050;
assign a1904 = ~a1902 & ~a1900;
assign a1906 = a1904 & a1880;
assign a1908 = a1906 & a1820;
assign a1910 = ~a1908 & ~a1022;
assign a1912 = a1774 & a824;
assign a1914 = ~a1912 & ~a1762;
assign a1916 = ~a1914 & ~a838;
assign a1918 = a1916 & ~a924;
assign a1920 = a1918 & ~a952;
assign a1922 = a1766 & ~a838;
assign a1924 = a1922 & ~a924;
assign a1926 = a1924 & ~a952;
assign a1928 = a1926 & ~a890;
assign a1930 = ~a1928 & ~a1920;
assign a1932 = ~a1930 & a974;
assign a1934 = a1922 & a924;
assign a1936 = a1934 & a952;
assign a1938 = a1828 & ~a838;
assign a1940 = ~a1938 & ~a1936;
assign a1942 = a1940 & ~a1926;
assign a1944 = ~a1942 & a890;
assign a1946 = ~a1944 & ~a1932;
assign a1948 = a1786 & ~a838;
assign a1950 = a1948 & ~a924;
assign a1952 = a1950 & ~a952;
assign a1954 = a1952 & a890;
assign a1956 = a1934 & ~a952;
assign a1958 = a1956 & a890;
assign a1960 = ~a1958 & ~a1954;
assign a1962 = ~a1960 & a974;
assign a1964 = ~a1962 & a1946;
assign a1966 = ~a1964 & ~a870;
assign a1968 = a1966 & a1036;
assign a1970 = a1968 & a1050;
assign a1972 = a1916 & a924;
assign a1974 = a1972 & ~a952;
assign a1976 = a1948 & a924;
assign a1978 = a1976 & ~a952;
assign a1980 = a1978 & a890;
assign a1982 = ~a1980 & ~a1974;
assign a1984 = ~a1982 & a974;
assign a1986 = a1976 & a952;
assign a1988 = a1804 & ~a838;
assign a1990 = ~a1988 & ~a1986;
assign a1992 = ~a1990 & a890;
assign a1994 = a1972 & a952;
assign a1996 = a1850 & a824;
assign a1998 = ~a1996 & ~a1826;
assign a2000 = ~a1998 & ~a838;
assign a2002 = ~a2000 & ~a1994;
assign a2004 = a2002 & ~a1992;
assign a2006 = a2004 & ~a1984;
assign a2008 = ~a2006 & ~a870;
assign a2010 = a2008 & i50;
assign a2012 = a2010 & a1036;
assign a2014 = a2012 & a1050;
assign a2016 = a2014 & l142;
assign a2018 = a2016 & ~l144;
assign a2020 = ~a2018 & ~a1970;
assign a2022 = a2016 & l144;
assign a2024 = a2008 & ~i50;
assign a2026 = a1954 & ~a974;
assign a2028 = a1956 & ~a890;
assign a2030 = a2028 & a974;
assign a2032 = ~a2030 & ~a2026;
assign a2034 = ~a1930 & ~a974;
assign a2036 = ~a1940 & ~a890;
assign a2038 = ~a2036 & ~a2034;
assign a2040 = a2038 & a2032;
assign a2042 = ~a2040 & ~a870;
assign a2044 = ~a2042 & ~a2024;
assign a2046 = ~a2044 & a1036;
assign a2048 = a2046 & a1050;
assign a2050 = a2048 & l142;
assign a2052 = ~a2050 & ~a2022;
assign a2054 = a2052 & a2020;
assign a2056 = ~a2054 & l140;
assign a2058 = ~a2056 & ~a1910;
assign a2060 = a2058 & ~a1650;
assign a2062 = a1598 & ~l144;
assign a2064 = ~a1538 & ~l146;
assign a2066 = a2064 & ~l142;
assign a2068 = a1542 & ~l146;
assign a2070 = a2068 & ~a1008;
assign a2072 = a2070 & ~l142;
assign a2074 = ~a2072 & ~a2066;
assign a2076 = ~a2074 & l144;
assign a2078 = ~a2076 & ~a2062;
assign a2080 = ~a2078 & ~l140;
assign a2082 = a2014 & ~l142;
assign a2084 = a2082 & l144;
assign a2086 = a2048 & ~l142;
assign a2088 = ~a2086 & ~a2084;
assign a2090 = ~a2088 & l140;
assign a2092 = ~a1726 & a974;
assign a2094 = a1734 & ~a1722;
assign a2096 = ~a2094 & a890;
assign a2098 = ~a2096 & ~a2092;
assign a2100 = ~a2098 & a870;
assign a2102 = a1738 & a1686;
assign a2104 = ~a2102 & a870;
assign a2106 = a2104 & ~i50;
assign a2108 = ~a2106 & ~a2100;
assign a2110 = ~a2108 & l146;
assign a2112 = a2110 & a1008;
assign a2114 = a2112 & ~l142;
assign a2116 = a2114 & ~l144;
assign a2118 = ~a2116 & ~a2090;
assign a2120 = a2118 & ~a2080;
assign a2122 = a2038 & a2002;
assign a2124 = ~a2122 & a870;
assign a2126 = a2124 & i50;
assign a2128 = a2126 & a1036;
assign a2130 = a2128 & ~a1050;
assign a2132 = a2130 & l142;
assign a2134 = a2124 & ~i50;
assign a2136 = ~a1946 & a870;
assign a2138 = ~a2136 & ~a2134;
assign a2140 = ~a2138 & a1036;
assign a2142 = a2140 & ~a1050;
assign a2144 = ~a2142 & ~a2132;
assign a2146 = ~a2144 & ~l140;
assign a2148 = a1772 & a952;
assign a2150 = a1912 & a838;
assign a2152 = a2150 & a924;
assign a2154 = a2152 & a952;
assign a2156 = a2154 & a890;
assign a2158 = ~a2156 & ~a2148;
assign a2160 = ~a2158 & a974;
assign a2162 = a2150 & ~a924;
assign a2164 = a2162 & ~a952;
assign a2166 = a1996 & a838;
assign a2168 = ~a2166 & ~a2164;
assign a2170 = ~a2168 & a890;
assign a2172 = ~a2170 & a1834;
assign a2174 = a2172 & ~a2160;
assign a2176 = ~a2174 & ~a870;
assign a2178 = a2176 & i50;
assign a2180 = a2178 & a1008;
assign a2182 = a2180 & ~a1036;
assign a2184 = a2182 & a1050;
assign a2186 = a2184 & l140;
assign a2188 = a2176 & ~i50;
assign a2190 = a2162 & a952;
assign a2192 = a2190 & a890;
assign a2194 = a2192 & ~a974;
assign a2196 = a1780 & a952;
assign a2198 = a2196 & ~a890;
assign a2200 = a2198 & a974;
assign a2202 = ~a2200 & ~a2194;
assign a2204 = a2202 & a1860;
assign a2206 = ~a2204 & ~a870;
assign a2208 = ~a2206 & ~a2188;
assign a2210 = ~a2208 & a1008;
assign a2212 = a2210 & ~a1036;
assign a2214 = a2212 & a1050;
assign a2216 = ~a2214 & ~a2186;
assign a2218 = a2216 & ~a1760;
assign a2220 = a2218 & ~a2146;
assign a2222 = ~a2220 & a1022;
assign a2224 = a1898 & a1036;
assign a2226 = a1870 & a1036;
assign a2228 = a2226 & ~a1050;
assign a2230 = a2104 & i50;
assign a2232 = a2230 & l146;
assign a2234 = a2232 & a1008;
assign a2236 = a2234 & ~l142;
assign a2238 = a2236 & ~l144;
assign a2240 = ~a2238 & ~a2228;
assign a2242 = a2240 & ~a2224;
assign a2244 = ~a2242 & ~a1022;
assign a2246 = ~a2244 & ~a2222;
assign a2248 = a2246 & a2120;
assign a2250 = ~a2248 & ~i48;
assign a2252 = a2130 & ~l142;
assign a2254 = ~a2252 & a2144;
assign a2256 = ~a2254 & l140;
assign a2258 = a1776 & ~a838;
assign a2260 = a2258 & ~a924;
assign a2262 = a2260 & a952;
assign a2264 = a2262 & ~a890;
assign a2266 = ~a1924 & ~a1918;
assign a2268 = ~a2266 & a952;
assign a2270 = ~a2268 & ~a2264;
assign a2272 = ~a2270 & ~a974;
assign a2274 = a2258 & a924;
assign a2276 = a2274 & a952;
assign a2278 = a2260 & ~a952;
assign a2280 = a1852 & ~a838;
assign a2282 = ~a2280 & ~a2278;
assign a2284 = a2282 & ~a2276;
assign a2286 = ~a2284 & ~a890;
assign a2288 = ~a2286 & ~a2272;
assign a2290 = ~a2288 & a870;
assign a2292 = a2290 & a1036;
assign a2294 = a2292 & ~a1050;
assign a2296 = ~a2294 & ~a2256;
assign a2298 = ~a2212 & ~a2182;
assign a2300 = ~a2298 & ~a1050;
assign a2302 = a2196 & a890;
assign a2304 = ~a2302 & ~a2192;
assign a2306 = ~a2304 & a974;
assign a2308 = ~a2306 & a1888;
assign a2310 = ~a2308 & ~a870;
assign a2312 = a2310 & a1008;
assign a2314 = a2312 & ~a1036;
assign a2316 = ~a2314 & ~a2300;
assign a2318 = a2316 & a2296;
assign a2320 = ~a2318 & a1022;
assign a2322 = a1490 & ~a838;
assign a2324 = a2322 & a924;
assign a2326 = a2324 & a952;
assign a2328 = a2326 & ~a890;
assign a2330 = ~a1720 & ~a1716;
assign a2332 = ~a2330 & a952;
assign a2334 = ~a2332 & ~a2328;
assign a2336 = ~a2334 & ~a974;
assign a2338 = a2324 & ~a952;
assign a2340 = a2322 & ~a924;
assign a2342 = a2340 & a952;
assign a2344 = a1524 & ~a838;
assign a2346 = ~a2344 & ~a2342;
assign a2348 = a2346 & ~a2338;
assign a2350 = ~a2348 & ~a890;
assign a2352 = ~a2350 & ~a2336;
assign a2354 = ~a2352 & a870;
assign a2356 = a2354 & l146;
assign a2358 = ~a2232 & ~a2110;
assign a2360 = ~a2358 & ~a1008;
assign a2362 = ~a2360 & ~a2356;
assign a2364 = ~a2362 & ~l142;
assign a2366 = a1700 & a890;
assign a2368 = ~a2366 & ~a1710;
assign a2370 = ~a2368 & a974;
assign a2372 = ~a2370 & a2098;
assign a2374 = ~a2372 & ~a870;
assign a2376 = a2374 & ~l146;
assign a2378 = a2376 & ~a1008;
assign a2380 = ~a2378 & ~a2364;
assign a2382 = ~a2380 & ~l144;
assign a2384 = ~a2382 & ~a2320;
assign a2386 = a2384 & ~a2250;
assign a2388 = a2386 & a2060;
assign a2390 = a2210 & a1036;
assign a2392 = a2390 & a1050;
assign a2394 = a1746 & a1008;
assign a2396 = a2394 & ~l144;
assign a2398 = ~a2396 & ~a2392;
assign a2400 = a2140 & a1050;
assign a2402 = a2400 & ~l140;
assign a2404 = ~a2402 & ~a2224;
assign a2406 = a2404 & a2398;
assign a2408 = ~a2406 & a1022;
assign a2410 = a1588 & ~l142;
assign a2412 = a2410 & ~l144;
assign a2414 = a2066 & ~l144;
assign a2416 = ~a2414 & ~a2086;
assign a2418 = a2416 & ~a2412;
assign a2420 = ~a2418 & ~l140;
assign a2422 = ~a2108 & ~l146;
assign a2424 = a2422 & a1008;
assign a2426 = a2424 & ~l142;
assign a2428 = a2426 & ~l144;
assign a2430 = ~a2428 & ~a2420;
assign a2432 = a2430 & ~a2408;
assign a2434 = a2128 & a1050;
assign a2436 = a2434 & l142;
assign a2438 = ~a2436 & ~a2400;
assign a2440 = ~a2438 & l140;
assign a2442 = a2180 & a1036;
assign a2444 = a2442 & ~a1050;
assign a2446 = a2444 & l140;
assign a2448 = a2390 & ~a1050;
assign a2450 = ~a2448 & ~a2446;
assign a2452 = a2450 & a1904;
assign a2454 = a2452 & ~a2440;
assign a2456 = ~a2454 & a1022;
assign a2458 = a1594 & ~l142;
assign a2460 = ~a2458 & ~a2410;
assign a2462 = ~a2460 & l144;
assign a2464 = ~a1548 & ~l142;
assign a2466 = a2464 & ~l144;
assign a2468 = ~a2466 & a2052;
assign a2470 = a2468 & ~a2462;
assign a2472 = ~a2470 & ~l140;
assign a2474 = a2422 & ~a1008;
assign a2476 = a2474 & ~l142;
assign a2478 = a2476 & ~l144;
assign a2480 = a2230 & ~l146;
assign a2482 = a2480 & ~a1008;
assign a2484 = a2482 & ~l142;
assign a2486 = a2484 & ~l144;
assign a2488 = a1752 & a1008;
assign a2490 = a2488 & ~a1036;
assign a2492 = a2490 & ~l144;
assign a2494 = ~a2492 & ~a2396;
assign a2496 = a2494 & ~a2486;
assign a2498 = ~a2496 & ~a1022;
assign a2500 = ~a2498 & ~a2478;
assign a2502 = a2500 & ~a2472;
assign a2504 = a2502 & ~a2456;
assign a2506 = a2504 & a2432;
assign a2508 = ~a2506 & ~i48;
assign a2510 = a2292 & a1050;
assign a2512 = a2312 & a1036;
assign a2514 = ~a2512 & ~a1818;
assign a2516 = a2514 & ~a2510;
assign a2518 = ~a2516 & a1022;
assign a2520 = a1568 & ~l142;
assign a2522 = a2520 & ~l144;
assign a2524 = a1642 & ~l142;
assign a2526 = ~a2524 & ~a1970;
assign a2528 = a2526 & ~a2522;
assign a2530 = ~a2528 & ~l140;
assign a2532 = a2354 & ~l146;
assign a2534 = a2532 & ~l142;
assign a2536 = a2376 & a1008;
assign a2538 = ~a2536 & ~a2534;
assign a2540 = ~a2538 & ~l144;
assign a2542 = ~a2540 & ~a2530;
assign a2544 = a2542 & ~a2518;
assign a2546 = a2544 & ~a2508;
assign a2548 = a2546 & a2388;
assign a2550 = ~a2548 & ~i46;
assign a2552 = a2152 & ~a952;
assign a2554 = a2552 & a890;
assign a2556 = a2554 & ~a974;
assign a2558 = a1790 & a952;
assign a2560 = a2558 & ~a890;
assign a2562 = a2560 & a974;
assign a2564 = ~a2562 & ~a2556;
assign a2566 = a2564 & a1812;
assign a2568 = ~a2566 & ~a870;
assign a2570 = a2568 & a1008;
assign a2572 = ~a2270 & a974;
assign a2574 = a2284 & ~a2262;
assign a2576 = ~a2574 & a890;
assign a2578 = ~a2576 & ~a2572;
assign a2580 = ~a2578 & a870;
assign a2582 = a2580 & a1036;
assign a2584 = ~a2582 & ~a2570;
assign a2586 = ~a2584 & a1022;
assign a2588 = ~a2334 & a974;
assign a2590 = a2348 & ~a2326;
assign a2592 = ~a2590 & a890;
assign a2594 = ~a2592 & ~a2588;
assign a2596 = ~a2594 & a870;
assign a2598 = a2596 & ~l142;
assign a2600 = a2340 & ~a952;
assign a2602 = a2600 & ~a890;
assign a2604 = a2602 & a974;
assign a2606 = a1706 & a952;
assign a2608 = a2606 & a890;
assign a2610 = a2608 & ~a974;
assign a2612 = ~a2610 & ~a2604;
assign a2614 = a2612 & a2352;
assign a2616 = ~a2614 & ~a870;
assign a2618 = a2616 & ~l146;
assign a2620 = ~a2618 & ~a2598;
assign a2622 = ~a2620 & ~l144;
assign a2624 = ~a2622 & ~a2586;
assign a2626 = ~a1624 & a974;
assign a2628 = a1634 & ~a1620;
assign a2630 = ~a2628 & a890;
assign a2632 = ~a2630 & ~a2626;
assign a2634 = ~a2632 & a870;
assign a2636 = a2634 & a1050;
assign a2638 = a1436 & ~a952;
assign a2640 = a2638 & a890;
assign a2642 = a2640 & ~a974;
assign a2644 = a1618 & a952;
assign a2646 = a2644 & ~a890;
assign a2648 = a2646 & a974;
assign a2650 = ~a2648 & ~a2642;
assign a2652 = a2650 & a1638;
assign a2654 = ~a2652 & ~a870;
assign a2656 = a2654 & ~l142;
assign a2658 = ~a2656 & ~a2636;
assign a2660 = ~a2658 & ~l140;
assign a2662 = ~a1796 & a974;
assign a2664 = a1808 & ~a1792;
assign a2666 = ~a2664 & a890;
assign a2668 = ~a2666 & ~a2662;
assign a2670 = ~a2668 & a870;
assign a2672 = a2670 & ~l146;
assign a2674 = a2672 & a1008;
assign a2676 = a2274 & ~a952;
assign a2678 = a2676 & ~a890;
assign a2680 = a2678 & a974;
assign a2682 = a1950 & a952;
assign a2684 = a2682 & a890;
assign a2686 = a2684 & ~a974;
assign a2688 = ~a2686 & ~a2680;
assign a2690 = a2688 & a2288;
assign a2692 = ~a2690 & ~a870;
assign a2694 = a2692 & a1036;
assign a2696 = a2694 & a1050;
assign a2698 = ~a2696 & ~a2674;
assign a2700 = a2698 & ~a2660;
assign a2702 = a2700 & a2624;
assign a2704 = a2702 & ~a2550;
assign a2706 = a2126 & ~a1036;
assign a2708 = a2706 & a1050;
assign a2710 = a2708 & l142;
assign a2712 = ~a2138 & ~a1036;
assign a2714 = a2712 & a1050;
assign a2716 = ~a2714 & ~a2710;
assign a2718 = ~a2716 & ~l140;
assign a2720 = ~a1744 & l146;
assign a2722 = a2720 & a1008;
assign a2724 = a1750 & l146;
assign a2726 = a2724 & a1008;
assign a2728 = a2726 & ~a1036;
assign a2730 = ~a2728 & ~a2722;
assign a2732 = ~a2730 & ~l144;
assign a2734 = a1896 & ~a1008;
assign a2736 = a2734 & a1036;
assign a2738 = a1868 & ~a1008;
assign a2740 = a2738 & a1036;
assign a2742 = a2740 & ~a1050;
assign a2744 = ~a2742 & ~a2736;
assign a2746 = a2744 & ~a2732;
assign a2748 = a2746 & ~a2718;
assign a2750 = ~a2748 & a1022;
assign a2752 = a2458 & ~l144;
assign a2754 = ~a2752 & ~a2412;
assign a2756 = ~a2754 & l140;
assign a2758 = a2442 & a1050;
assign a2760 = a2758 & l140;
assign a2762 = ~a2760 & ~a2392;
assign a2764 = ~a2762 & ~a1022;
assign a2766 = ~a2764 & ~a2756;
assign a2768 = a2012 & ~a1050;
assign a2770 = a2768 & ~l142;
assign a2772 = a2770 & l144;
assign a2774 = a2046 & ~a1050;
assign a2776 = a2774 & ~l142;
assign a2778 = ~a2776 & ~a2772;
assign a2780 = ~a2778 & ~l140;
assign a2782 = a2426 & l144;
assign a2784 = ~a2782 & ~a2780;
assign a2786 = a2480 & a1008;
assign a2788 = a2786 & ~l142;
assign a2790 = a2788 & l144;
assign a2792 = a2790 & ~a1022;
assign a2794 = ~a2070 & ~a2064;
assign a2796 = ~a2794 & l142;
assign a2798 = a2796 & ~l144;
assign a2800 = a2798 & ~l140;
assign a2802 = ~a2800 & ~a2792;
assign a2804 = a2802 & a2784;
assign a2806 = a2804 & a2766;
assign a2808 = a2806 & ~a2750;
assign a2810 = ~a2808 & ~i48;
assign a2812 = a2708 & ~l142;
assign a2814 = ~a2812 & a2716;
assign a2816 = ~a2814 & l140;
assign a2818 = a2290 & ~a1036;
assign a2820 = a2818 & a1050;
assign a2822 = ~a2820 & ~a2816;
assign a2824 = ~a2822 & a1022;
assign a2826 = a2462 & l140;
assign a2828 = a1602 & ~l142;
assign a2830 = a2828 & l144;
assign a2832 = ~a2830 & ~a2524;
assign a2834 = ~a2832 & l140;
assign a2836 = ~a2834 & ~a2826;
assign a2838 = a2836 & ~a2824;
assign a2840 = a2444 & ~l140;
assign a2842 = a2726 & a1036;
assign a2844 = a2842 & ~l144;
assign a2846 = ~a2844 & ~a2840;
assign a2848 = a2846 & a2450;
assign a2850 = a2848 & ~a2732;
assign a2852 = ~a2850 & ~a1022;
assign a2854 = a1816 & ~a1008;
assign a2856 = ~a2738 & ~a2734;
assign a2858 = ~a2856 & ~a1036;
assign a2860 = ~a2858 & ~a2854;
assign a2862 = ~a2860 & a1022;
assign a2864 = ~a2862 & ~a2852;
assign a2866 = ~a1572 & l142;
assign a2868 = a2866 & ~l144;
assign a2870 = ~a2774 & ~a2768;
assign a2872 = ~a2870 & l142;
assign a2874 = a1968 & ~a1050;
assign a2876 = ~a2874 & ~a2872;
assign a2878 = a2876 & ~a2868;
assign a2880 = ~a2878 & ~l140;
assign a2882 = ~a2534 & ~a2476;
assign a2884 = ~a2882 & l144;
assign a2886 = a2484 & l144;
assign a2888 = a2512 & ~a1022;
assign a2890 = a2374 & l146;
assign a2892 = a2890 & a1008;
assign a2894 = a2892 & ~l144;
assign a2896 = ~a2894 & ~a2888;
assign a2898 = a2896 & ~a2886;
assign a2900 = a2898 & ~a2884;
assign a2902 = a2900 & ~a2880;
assign a2904 = a2902 & a2864;
assign a2906 = a2904 & a2838;
assign a2908 = a2906 & ~a2810;
assign a2910 = ~a2908 & ~i46;
assign a2912 = ~a2770 & ~a1604;
assign a2914 = ~a2912 & ~l144;
assign a2916 = a2876 & a2778;
assign a2918 = a2916 & ~a2914;
assign a2920 = ~a2918 & l140;
assign a2922 = ~a2598 & ~a2364;
assign a2924 = ~a2922 & l144;
assign a2926 = ~a2924 & ~a2920;
assign a2928 = a2184 & ~l140;
assign a2930 = a2740 & a1050;
assign a2932 = ~a2930 & ~a2928;
assign a2934 = ~a2570 & a2216;
assign a2936 = a2934 & a2932;
assign a2938 = a2744 & a2316;
assign a2940 = a2938 & a2860;
assign a2942 = a2940 & a2936;
assign a2944 = ~a2942 & ~a1022;
assign a2946 = ~a2944 & a2926;
assign a2948 = ~a2062 & a1646;
assign a2950 = ~a2948 & l140;
assign a2952 = a2068 & a1008;
assign a2954 = a2952 & l142;
assign a2956 = ~a2954 & ~a2796;
assign a2958 = a2956 & ~a2866;
assign a2960 = ~a2958 & l144;
assign a2962 = a2654 & l142;
assign a2964 = ~a2962 & ~a2960;
assign a2966 = ~a2964 & ~l140;
assign a2968 = a2694 & ~a1050;
assign a2970 = a2672 & ~a1008;
assign a2972 = a2636 & l140;
assign a2974 = ~a2972 & ~a2970;
assign a2976 = a2974 & ~a2968;
assign a2978 = a2616 & l146;
assign a2980 = ~a2890 & ~a2724;
assign a2982 = a2980 & ~a2720;
assign a2984 = ~a2982 & ~a1008;
assign a2986 = ~a2984 & ~a2978;
assign a2988 = ~a2986 & ~l144;
assign a2990 = ~a2988 & a2976;
assign a2992 = a2580 & ~a1036;
assign a2994 = ~a2818 & ~a2706;
assign a2996 = a2994 & ~a2712;
assign a2998 = ~a2996 & ~a1050;
assign a3000 = ~a2998 & ~a2992;
assign a3002 = ~a3000 & a1022;
assign a3004 = ~a2236 & ~a2114;
assign a3006 = ~a3004 & l144;
assign a3008 = ~a3006 & ~a3002;
assign a3010 = a3008 & a2990;
assign a3012 = a3010 & ~a2966;
assign a3014 = a3012 & ~a2950;
assign a3016 = a3014 & a2946;
assign a3018 = a3016 & ~a2910;
assign a3020 = a3018 & a2704;
assign a3022 = ~a3020 & ~i44;
assign a3024 = a2676 & a890;
assign a3026 = ~a3024 & ~a2684;
assign a3028 = ~a3026 & a974;
assign a3030 = ~a3028 & a2578;
assign a3032 = ~a3030 & ~a870;
assign a3034 = a3032 & a1036;
assign a3036 = a1990 & ~a1950;
assign a3038 = ~a3036 & ~a890;
assign a3040 = ~a2676 & ~a1956;
assign a3042 = a1978 & ~a890;
assign a3044 = ~a3042 & ~a1974;
assign a3046 = a3044 & a3040;
assign a3048 = ~a3046 & ~a974;
assign a3050 = ~a3048 & ~a3038;
assign a3052 = ~a3050 & a870;
assign a3054 = a3052 & a1022;
assign a3056 = ~a2638 & ~a1502;
assign a3058 = a3056 & a1460;
assign a3060 = ~a3058 & ~a890;
assign a3062 = ~a2644 & ~a1496;
assign a3064 = a1438 & ~a890;
assign a3066 = ~a3064 & ~a1426;
assign a3068 = a3066 & a3062;
assign a3070 = ~a3068 & ~a974;
assign a3072 = ~a3070 & ~a3060;
assign a3074 = ~a3072 & a870;
assign a3076 = a3074 & a1050;
assign a3078 = ~a3076 & ~a3054;
assign a3080 = a3078 & ~a3034;
assign a3082 = a2558 & a890;
assign a3084 = ~a3082 & ~a2554;
assign a3086 = ~a3084 & a974;
assign a3088 = ~a3086 & a2668;
assign a3090 = ~a3088 & ~a870;
assign a3092 = a3090 & a1008;
assign a3094 = a2600 & a890;
assign a3096 = ~a3094 & ~a2608;
assign a3098 = ~a3096 & a974;
assign a3100 = ~a3098 & a2594;
assign a3102 = ~a3100 & ~a870;
assign a3104 = a3102 & ~l144;
assign a3106 = ~a3104 & ~a3092;
assign a3108 = ~a2552 & ~a2190;
assign a3110 = a3108 & a2168;
assign a3112 = ~a3110 & ~a890;
assign a3114 = a2154 & ~a890;
assign a3116 = ~a3114 & ~a2148;
assign a3118 = ~a2558 & ~a2196;
assign a3120 = a3118 & a3116;
assign a3122 = ~a3120 & ~a974;
assign a3124 = ~a3122 & ~a3112;
assign a3126 = ~a3124 & a870;
assign a3128 = a3126 & ~l146;
assign a3130 = ~a1706 & a1676;
assign a3132 = ~a3130 & ~a890;
assign a3134 = ~a2600 & ~a1700;
assign a3136 = a1664 & ~a890;
assign a3138 = ~a3136 & ~a1658;
assign a3140 = a3138 & a3134;
assign a3142 = ~a3140 & ~a974;
assign a3144 = ~a3142 & ~a3132;
assign a3146 = ~a3144 & a870;
assign a3148 = a3146 & ~l142;
assign a3150 = ~a3148 & ~a3128;
assign a3152 = a2644 & a890;
assign a3154 = ~a3152 & ~a2640;
assign a3156 = ~a3154 & a974;
assign a3158 = ~a3156 & a2632;
assign a3160 = ~a3158 & ~a870;
assign a3162 = a3160 & ~l140;
assign a3164 = ~a3162 & a3150;
assign a3166 = a3164 & a3106;
assign a3168 = a3166 & a3080;
assign a3170 = a3168 & ~a3022;
assign a3172 = ~a3170 & i54;
assign a3174 = ~a1592 & a1586;
assign a3176 = ~a3174 & ~a1050;
assign a3178 = a3176 & ~l142;
assign a3180 = a3178 & ~l144;
assign a3182 = a2010 & ~a1036;
assign a3184 = a3182 & a1050;
assign a3186 = a3184 & ~l142;
assign a3188 = a3186 & l144;
assign a3190 = ~a2044 & ~a1036;
assign a3192 = a3190 & a1050;
assign a3194 = a3192 & ~l142;
assign a3196 = ~a3194 & ~a3188;
assign a3198 = a3196 & ~a3180;
assign a3200 = ~a3198 & ~l140;
assign a3202 = a2072 & ~l144;
assign a3204 = ~a3202 & ~a2414;
assign a3206 = ~a3204 & l140;
assign a3208 = a2424 & l142;
assign a3210 = a3208 & ~l144;
assign a3212 = ~a3210 & ~a3206;
assign a3214 = a3212 & ~a3200;
assign a3216 = ~a1894 & l146;
assign a3218 = a3216 & a1008;
assign a3220 = a3218 & a1036;
assign a3222 = a1866 & l146;
assign a3224 = a3222 & a1008;
assign a3226 = a3224 & a1036;
assign a3228 = a3226 & ~a1050;
assign a3230 = ~a3228 & ~a3220;
assign a3232 = ~a2490 & ~a2394;
assign a3234 = ~a3232 & l144;
assign a3236 = a2178 & ~a1008;
assign a3238 = a3236 & a1036;
assign a3240 = a3238 & a1050;
assign a3242 = a3240 & l140;
assign a3244 = ~a2208 & ~a1008;
assign a3246 = a3244 & a1036;
assign a3248 = a3246 & a1050;
assign a3250 = ~a3248 & ~a3242;
assign a3252 = a3250 & ~a3234;
assign a3254 = a3252 & a3230;
assign a3256 = ~a3254 & a1022;
assign a3258 = a2786 & l142;
assign a3260 = a3258 & ~l144;
assign a3262 = a2436 & ~l140;
assign a3264 = ~a3262 & ~a2402;
assign a3266 = a3264 & ~a3260;
assign a3268 = ~a3266 & ~a1022;
assign a3270 = ~a3268 & ~a3256;
assign a3272 = a3270 & a3214;
assign a3274 = ~a3272 & ~i48;
assign a3276 = ~a3246 & ~a3238;
assign a3278 = ~a3276 & ~a1050;
assign a3280 = a2310 & ~a1008;
assign a3282 = a3280 & a1036;
assign a3284 = ~a3282 & ~a3278;
assign a3286 = a1814 & l146;
assign a3288 = a3286 & a1008;
assign a3290 = ~a3224 & ~a3218;
assign a3292 = ~a3290 & ~a1036;
assign a3294 = ~a3292 & ~a3288;
assign a3296 = a3294 & a3284;
assign a3298 = ~a3296 & a1022;
assign a3300 = ~a3234 & ~a2510;
assign a3302 = a2434 & ~l142;
assign a3304 = a3302 & l140;
assign a3306 = a2488 & a1036;
assign a3308 = a3306 & l144;
assign a3310 = ~a3308 & ~a3304;
assign a3312 = a3310 & ~a2440;
assign a3314 = a3312 & a3300;
assign a3316 = ~a3314 & ~a1022;
assign a3318 = ~a3316 & ~a3298;
assign a3320 = a1600 & ~a1050;
assign a3322 = a3320 & ~l142;
assign a3324 = ~a3322 & ~a3178;
assign a3326 = ~a3324 & l144;
assign a3328 = a1640 & ~a1050;
assign a3330 = a3328 & ~l142;
assign a3332 = ~a3330 & ~a3326;
assign a3334 = ~a3332 & ~l140;
assign a3336 = ~a2532 & ~a2482;
assign a3338 = a3336 & ~a2474;
assign a3340 = ~a3338 & l142;
assign a3342 = a3340 & ~l144;
assign a3344 = a2536 & l144;
assign a3346 = ~a3344 & ~a3342;
assign a3348 = ~a3192 & ~a3184;
assign a3350 = ~a3348 & l142;
assign a3352 = a1966 & ~a1036;
assign a3354 = a3352 & a1050;
assign a3356 = ~a3354 & ~a3350;
assign a3358 = ~a3356 & ~l140;
assign a3360 = a1574 & ~l144;
assign a3362 = a3360 & l140;
assign a3364 = ~a3362 & ~a3358;
assign a3366 = a3364 & a3346;
assign a3368 = a3366 & ~a3334;
assign a3370 = a3368 & a3318;
assign a3372 = a3370 & ~a3274;
assign a3374 = ~a3372 & ~i46;
assign a3376 = a3294 & ~a2146;
assign a3378 = a3226 & a1050;
assign a3380 = a2252 & ~l140;
assign a3382 = ~a3380 & ~a3378;
assign a3384 = a3382 & a3230;
assign a3386 = a3384 & a2296;
assign a3388 = a3386 & a3376;
assign a3390 = ~a3388 & ~a1022;
assign a3392 = ~a2596 & ~a2234;
assign a3394 = a3392 & ~a2112;
assign a3396 = a3394 & a2362;
assign a3398 = ~a3396 & l142;
assign a3400 = a3398 & ~l144;
assign a3402 = a3196 & ~a2656;
assign a3404 = a3402 & a3356;
assign a3406 = a3186 & ~l144;
assign a3408 = a2952 & ~l142;
assign a3410 = a3408 & l144;
assign a3412 = ~a3410 & ~a3406;
assign a3414 = a3412 & ~a2076;
assign a3416 = a3414 & ~a1576;
assign a3418 = a3416 & a3404;
assign a3420 = ~a3418 & l140;
assign a3422 = ~a3420 & ~a3400;
assign a3424 = a2634 & ~a1050;
assign a3426 = ~a3328 & ~a3320;
assign a3428 = a3426 & ~a3176;
assign a3430 = ~a3428 & l142;
assign a3432 = ~a3430 & ~a3424;
assign a3434 = ~a3432 & ~l140;
assign a3436 = a2568 & ~a1008;
assign a3438 = ~a3280 & ~a3236;
assign a3440 = a3438 & ~a3244;
assign a3442 = ~a3440 & ~a1036;
assign a3444 = ~a3442 & ~a3436;
assign a3446 = ~a3444 & a1022;
assign a3448 = ~a2618 & ~a2378;
assign a3450 = a3448 & ~a1876;
assign a3452 = a3450 & a1758;
assign a3454 = ~a3452 & l144;
assign a3456 = a2692 & ~a1036;
assign a3458 = a3456 & a1050;
assign a3460 = a2670 & l146;
assign a3462 = a3460 & a1008;
assign a3464 = a2582 & ~a1022;
assign a3466 = ~a3464 & ~a3462;
assign a3468 = a3466 & ~a3458;
assign a3470 = a3468 & ~a3454;
assign a3472 = a3470 & ~a3446;
assign a3474 = a3472 & ~a3434;
assign a3476 = a3474 & a3422;
assign a3478 = a3476 & ~a3390;
assign a3480 = a3478 & ~a3374;
assign a3482 = ~a3480 & ~i44;
assign a3484 = ~a3258 & a2730;
assign a3486 = a3484 & ~a3208;
assign a3488 = ~a3102 & ~a2892;
assign a3490 = a3488 & ~a2842;
assign a3492 = a3490 & a2986;
assign a3494 = a3492 & ~a3340;
assign a3496 = a3494 & a3486;
assign a3498 = a3496 & ~a3398;
assign a3500 = ~a3498 & l144;
assign a3502 = ~a3240 & ~a2812;
assign a3504 = ~a3502 & ~l140;
assign a3506 = a3504 & ~a1022;
assign a3508 = ~a3460 & ~a3222;
assign a3510 = ~a3286 & ~a3090;
assign a3512 = a3510 & ~a3216;
assign a3514 = a3512 & a3508;
assign a3516 = ~a3514 & ~a1008;
assign a3518 = a3160 & l140;
assign a3520 = a3032 & ~a1036;
assign a3522 = ~a3520 & ~a3518;
assign a3524 = a3146 & l142;
assign a3526 = a3126 & l146;
assign a3528 = ~a3526 & ~a3524;
assign a3530 = a3052 & ~a1022;
assign a3532 = a3074 & ~a1050;
assign a3534 = ~a3532 & ~a3530;
assign a3536 = a3534 & a3528;
assign a3538 = a3536 & a3522;
assign a3540 = ~a3352 & ~a3182;
assign a3542 = ~a3456 & ~a3190;
assign a3544 = a3542 & a3540;
assign a3546 = ~a3544 & ~a1050;
assign a3548 = ~a3546 & a3538;
assign a3550 = a3548 & ~a3516;
assign a3552 = a3550 & ~a3506;
assign a3554 = a3552 & ~a3500;
assign a3556 = ~a3322 & ~a2954;
assign a3558 = ~a3556 & ~l144;
assign a3560 = ~a3558 & ~a3180;
assign a3562 = a3560 & a2964;
assign a3564 = ~a2868 & ~a2798;
assign a3566 = a3564 & a3432;
assign a3568 = a3566 & a3332;
assign a3570 = a3568 & a3562;
assign a3572 = ~a3570 & l140;
assign a3574 = a3000 & ~a2718;
assign a3576 = a3444 & a3250;
assign a3578 = a3576 & a3284;
assign a3580 = a3578 & a3574;
assign a3582 = a3580 & a2822;
assign a3584 = ~a3582 & ~a1022;
assign a3586 = ~a3584 & ~a3572;
assign a3588 = a3586 & a3554;
assign a3590 = a3588 & ~a3482;
assign a3592 = a3590 & ~a3172;
assign a3594 = ~a3592 & i52;
assign a3596 = a3594 & ~l160;
assign a3598 = ~a3596 & a1406;
assign a3600 = a3598 & i70;
assign a3602 = a1402 & ~a1096;
assign a3604 = a1394 & ~a1300;
assign a3606 = ~a3604 & ~a3602;
assign a3608 = a1390 & ~a1374;
assign a3610 = a1398 & ~a1226;
assign a3612 = ~a3610 & ~a3608;
assign a3614 = a3612 & a3606;
assign a3616 = a1406 & ~a1138;
assign a3618 = a1406 & i54;
assign a3620 = ~a3618 & ~a3616;
assign a3622 = a3620 & a3614;
assign a3624 = ~a3622 & i64;
assign a3626 = ~a3624 & l172;
assign a3628 = a3622 & ~l172;
assign a3630 = ~a3628 & ~a3626;
assign a3632 = a3630 & i62;
assign a3634 = a3624 & l172;
assign a3636 = ~a3622 & ~l172;
assign a3638 = a3636 & l174;
assign a3640 = ~a3638 & ~a3634;
assign a3642 = ~a3640 & a3632;
assign a3644 = ~a3642 & ~a3628;
assign a3646 = a3636 & ~l174;
assign a3648 = ~a3646 & a3644;
assign a3650 = ~a3626 & i66;
assign a3652 = ~a3650 & a3648;
assign a3654 = ~a3622 & l176;
assign a3656 = a1390 & i56;
assign a3658 = ~i60 & ~i58;
assign a3660 = ~a3658 & i56;
assign a3662 = ~a3660 & i58;
assign a3664 = ~a3660 & i60;
assign a3666 = a3664 & a1394;
assign a3668 = ~a3664 & a1398;
assign a3670 = ~a3668 & ~a3666;
assign a3672 = ~a3670 & a3662;
assign a3674 = a3664 & a1402;
assign a3676 = ~a3664 & a1406;
assign a3678 = ~a3676 & ~a3674;
assign a3680 = ~a3678 & ~a3662;
assign a3682 = ~a3680 & ~a3672;
assign a3684 = ~a3682 & ~i56;
assign a3686 = ~a3684 & ~a3656;
assign a3688 = ~a3686 & a3614;
assign a3690 = ~a3688 & a1406;
assign a3692 = a3688 & ~i56;
assign a3694 = ~a3692 & ~a3690;
assign a3696 = ~a3694 & ~a3608;
assign a3698 = ~a3696 & ~a3616;
assign a3700 = a3688 & a3664;
assign a3702 = ~a3700 & a1406;
assign a3704 = a3702 & a3606;
assign a3706 = ~a3704 & ~a3616;
assign a3708 = a3688 & a3662;
assign a3710 = ~a3610 & ~a3604;
assign a3712 = a3710 & ~a3708;
assign a3714 = ~a3712 & ~a3616;
assign a3716 = ~a3714 & ~a3706;
assign a3718 = a3716 & a3698;
assign a3720 = a3718 & a810;
assign a3722 = a3714 & a3706;
assign a3724 = a3722 & a1306;
assign a3726 = a3714 & ~a3706;
assign a3728 = a3726 & a1230;
assign a3730 = ~a3714 & ~a3698;
assign a3732 = a3730 & a3706;
assign a3734 = a1040 & ~a810;
assign a3736 = ~a1040 & a810;
assign a3738 = ~a3736 & ~a3734;
assign a3740 = a3738 & a3732;
assign a3742 = a3716 & ~a3698;
assign a3744 = a3742 & ~a810;
assign a3746 = ~a3744 & ~a3740;
assign a3748 = a3746 & ~a3728;
assign a3750 = a3748 & ~a3724;
assign a3754 = a3752 & l178;
assign a3756 = ~a3754 & a3654;
assign a3758 = ~a3752 & ~l178;
assign a3760 = ~a3758 & a3756;
assign a3762 = a3716 & ~a838;
assign a3764 = a3762 & a3698;
assign a3766 = ~a1040 & ~a992;
assign a3768 = ~a3766 & a3722;
assign a3770 = a3726 & a838;
assign a3772 = a3766 & a3732;
assign a3774 = a3762 & ~a3698;
assign a3776 = ~a3774 & ~a3772;
assign a3778 = a3776 & ~a3770;
assign a3780 = a3778 & ~a3768;
assign a3784 = a3782 & l180;
assign a3786 = ~a3784 & a3760;
assign a3788 = ~a3782 & ~l180;
assign a3790 = ~a3788 & a3786;
assign a3792 = ~a3706 & a870;
assign a3794 = ~a3698 & a870;
assign a3796 = ~a3794 & a3706;
assign a3800 = ~a3798 & l182;
assign a3802 = ~a3800 & a3790;
assign a3804 = a3798 & ~l182;
assign a3806 = ~a3804 & a3802;
assign a3808 = a3806 & a792;
assign a3810 = a3808 & ~a3652;
assign a3812 = ~a3810 & ~a3632;
assign a3814 = ~i76 & ~i72;
assign a3816 = ~a3814 & i74;
assign a3818 = ~a3816 & i72;
assign a3820 = ~a3706 & ~a3622;
assign a3822 = a3820 & ~a3714;
assign a3824 = a3822 & a3698;
assign a3826 = ~a3824 & a1390;
assign a3828 = a3826 & i74;
assign a3830 = ~a3816 & i76;
assign a3832 = a3706 & ~a3622;
assign a3834 = a3832 & a3714;
assign a3836 = ~a3834 & a1394;
assign a3838 = a3836 & a3818;
assign a3840 = a3820 & a3714;
assign a3842 = ~a3840 & a1398;
assign a3844 = a3842 & ~a3818;
assign a3846 = ~a3844 & ~a3838;
assign a3848 = ~a3846 & a3830;
assign a3850 = a3832 & a3730;
assign a3852 = ~a3850 & a1402;
assign a3854 = a3852 & a3818;
assign a3856 = a3822 & ~a3698;
assign a3858 = ~a3856 & a1406;
assign a3860 = a3858 & ~a3818;
assign a3862 = ~a3860 & ~a3854;
assign a3864 = ~a3862 & ~a3830;
assign a3866 = ~a3864 & ~a3848;
assign a3868 = ~a3866 & ~i74;
assign a3870 = ~a3868 & ~a3828;
assign a3872 = ~a3870 & a3818;
assign a3874 = a3870 & ~a3858;
assign a3876 = ~a3874 & ~a3872;
assign a3878 = a3876 & a3706;
assign a3880 = ~a3848 & a3714;
assign a3882 = ~a3880 & ~a3878;
assign a3884 = a3848 & ~a3714;
assign a3886 = ~a3884 & ~a3882;
assign a3888 = ~a3828 & a3598;
assign a3890 = a3888 & a3698;
assign a3892 = ~a3890 & ~a3886;
assign a3894 = ~a3888 & ~a3698;
assign a3896 = ~a3894 & ~a3892;
assign a3898 = ~a3896 & ~a3812;
assign a3900 = ~a3898 & a3600;
assign a3902 = ~a3900 & a804;
assign a3904 = ~a3170 & ~i54;
assign a3906 = a3904 & i52;
assign a3908 = ~a2704 & i44;
assign a3910 = a3908 & i54;
assign a3912 = a3480 & a3018;
assign a3914 = ~a3912 & i44;
assign a3916 = ~a2486 & a1880;
assign a3918 = ~a3260 & ~a2790;
assign a3920 = a3918 & a3382;
assign a3922 = a3920 & a3916;
assign a3924 = a2846 & ~a2238;
assign a3926 = a3924 & a3310;
assign a3928 = ~a3504 & a2932;
assign a3930 = a3928 & a3926;
assign a3932 = a3930 & a3922;
assign a3934 = ~a3932 & a1022;
assign a3936 = ~a3302 & ~a2758;
assign a3938 = ~a3936 & ~l140;
assign a3940 = a2226 & a1050;
assign a3942 = a3306 & ~l144;
assign a3944 = ~a3942 & ~a3940;
assign a3946 = a3944 & ~a3938;
assign a3948 = ~a3946 & ~a1022;
assign a3950 = ~a3408 & ~a2082;
assign a3952 = a3950 & ~a2828;
assign a3954 = ~a3952 & ~l144;
assign a3956 = a3954 & l140;
assign a3958 = ~a3956 & ~a3948;
assign a3960 = a1550 & ~l142;
assign a3962 = a3960 & ~l144;
assign a3964 = ~a3962 & ~a2018;
assign a3966 = a3964 & ~a2914;
assign a3968 = a3412 & ~a2830;
assign a3970 = a3968 & ~a3558;
assign a3972 = a3970 & a3966;
assign a3974 = ~a3972 & ~l140;
assign a3976 = ~a3974 & a3958;
assign a3978 = a3976 & ~a3934;
assign a3980 = a3954 & ~l140;
assign a3982 = a2788 & ~l144;
assign a3984 = ~a3982 & a3946;
assign a3986 = ~a3984 & a1022;
assign a3988 = ~a3986 & ~a3980;
assign a3990 = i56 & i54;
assign a3992 = ~a3990 & ~a3988;
assign a3994 = ~a3992 & a3978;
assign a3996 = ~a3994 & i74;
assign a3998 = ~a3996 & ~a3914;
assign a4000 = a3998 & ~a3910;
assign a4002 = a4000 & ~a3906;
assign a4004 = i76 & ~i72;
assign a4006 = ~a2504 & i48;
assign a4008 = ~a2432 & i48;
assign a4010 = a4008 & i54;
assign a4012 = a3664 & i58;
assign a4014 = a4012 & a4010;
assign a4016 = ~a4014 & ~a4006;
assign a4018 = a3372 & a2908;
assign a4020 = ~a4018 & i46;
assign a4022 = ~a4020 & a4016;
assign a4024 = ~a2546 & i46;
assign a4026 = ~i60 & ~i56;
assign a4028 = a4026 & i58;
assign a4030 = a4028 & i54;
assign a4032 = ~a4030 & a4024;
assign a4034 = ~a4032 & a4022;
assign a4036 = ~a4034 & a4004;
assign a4038 = ~a3908 & ~i76;
assign a4040 = ~a4008 & i76;
assign a4042 = ~a4040 & ~a4038;
assign a4044 = a4042 & ~i54;
assign a4046 = a2808 & a2248;
assign a4048 = a4046 & a3272;
assign a4050 = ~a4048 & i48;
assign a4052 = ~a4012 & a4010;
assign a4054 = a3990 & ~a3988;
assign a4056 = ~a2760 & ~a2492;
assign a4058 = ~a3262 & ~a2228;
assign a4060 = a4058 & a4056;
assign a4062 = ~a4060 & a1022;
assign a4064 = ~a3202 & ~a2084;
assign a4066 = a4064 & ~a2752;
assign a4068 = ~a4066 & ~l140;
assign a4070 = a3982 & ~a1022;
assign a4072 = ~a4070 & ~a4068;
assign a4074 = a4072 & ~a4062;
assign a4076 = a4074 & ~a4054;
assign a4078 = a4076 & ~a4052;
assign a4080 = a4078 & ~a4050;
assign a4082 = ~a4080 & i76;
assign a4084 = a4030 & a4024;
assign a4086 = ~a2388 & i46;
assign a4088 = ~a4086 & ~a4084;
assign a4090 = ~a4088 & ~i76;
assign a4092 = ~a4090 & ~a4082;
assign a4094 = a4092 & ~a4044;
assign a4096 = ~a4094 & i72;
assign a4098 = ~a4096 & ~a4036;
assign a4100 = ~a4098 & ~i74;
assign a4102 = ~a4100 & a4002;
assign a4104 = ~a4102 & ~l160;
assign a4106 = ~a4104 & a3598;
assign a4108 = a4106 & i78;
assign a4110 = ~i84 & ~i80;
assign a4112 = ~a4110 & i82;
assign a4114 = ~a4112 & i80;
assign a4116 = a3826 & ~i74;
assign a4118 = a4116 & i82;
assign a4120 = ~a4112 & i84;
assign a4122 = ~a3876 & a3848;
assign a4124 = ~a4122 & ~a3828;
assign a4126 = a4124 & a3836;
assign a4128 = a4126 & a4114;
assign a4130 = a3876 & a3848;
assign a4132 = ~a4130 & a3842;
assign a4134 = a4132 & a4124;
assign a4136 = a4134 & ~a4114;
assign a4138 = ~a4136 & ~a4128;
assign a4140 = ~a4138 & a4120;
assign a4142 = ~a4140 & ~a4118;
assign a4144 = a3888 & ~a3848;
assign a4146 = a4144 & a3876;
assign a4148 = a4146 & a3852;
assign a4150 = ~a4120 & a4114;
assign a4152 = a4150 & a4148;
assign a4154 = ~a4152 & a4142;
assign a4156 = ~a4154 & a4114;
assign a4158 = ~a4134 & ~a4126;
assign a4160 = a4158 & ~a4148;
assign a4162 = a4160 & a4116;
assign a4164 = ~a4148 & a4134;
assign a4166 = ~a4164 & ~a4162;
assign a4168 = a4166 & a4154;
assign a4170 = ~a4168 & ~a4156;
assign a4172 = a4170 & a3706;
assign a4174 = ~a4158 & ~a4148;
assign a4176 = a4174 & a4154;
assign a4178 = ~a4176 & ~a4140;
assign a4180 = a4178 & a3714;
assign a4182 = ~a4180 & ~a4172;
assign a4184 = ~a4178 & ~a3714;
assign a4186 = ~a4184 & ~a4182;
assign a4188 = a4160 & a4154;
assign a4190 = ~a4188 & ~a4118;
assign a4192 = a4190 & a3698;
assign a4194 = ~a4192 & ~a4186;
assign a4196 = ~a4190 & ~a3698;
assign a4198 = ~a4196 & ~a4194;
assign a4200 = ~a4198 & ~a3812;
assign a4202 = ~a4200 & a4108;
assign a4204 = a4202 & a3902;
assign a4206 = a4204 & i68;
assign a4208 = a3900 & a804;
assign a4210 = a4208 & i86;
assign a4212 = ~a4210 & ~a4206;
assign a4214 = a1406 & a804;
assign a4216 = ~l188 & l102;
assign a4218 = ~a756 & ~l102;
assign a4220 = ~a4218 & ~a4216;
assign a4222 = ~a4220 & ~a4214;
assign a4226 = ~l190 & l102;
assign a4228 = a758 & ~l102;
assign a4230 = ~a4228 & ~a4226;
assign a4232 = a4230 & i88;
assign a4236 = a4204 & ~i68;
assign a4238 = a4208 & ~i86;
assign a4240 = ~a4238 & ~a4236;
assign a4242 = ~a3812 & a796;
assign a4244 = a4242 & a4240;
assign a4246 = ~a4244 & ~a762;
assign a4250 = a4212 & a802;
assign a4252 = ~a4250 & ~a762;
assign a4254 = ~a952 & l118;
assign a4256 = a3766 & a1390;
assign a4258 = a1394 & ~a838;
assign a4260 = a1406 & ~a870;
assign a4262 = ~a4260 & ~a1402;
assign a4264 = a4262 & ~a838;
assign a4266 = ~a4262 & a838;
assign a4268 = ~a4266 & ~a4264;
assign a4270 = ~a4268 & ~a1398;
assign a4272 = ~a3766 & a1398;
assign a4274 = ~a4272 & ~a4270;
assign a4276 = ~a4274 & ~a1394;
assign a4278 = ~a4276 & ~a4258;
assign a4280 = ~a4278 & ~a1390;
assign a4282 = ~a4280 & ~a4256;
assign a4284 = ~a4282 & ~l118;
assign a4288 = ~a974 & l118;
assign a4290 = a1406 & ~a1402;
assign a4292 = ~a4290 & ~a1398;
assign a4294 = ~a4292 & ~a1394;
assign a4296 = ~a4294 & ~a1390;
assign a4298 = a4296 & ~a870;
assign a4300 = ~a4296 & a870;
assign a4302 = ~a4300 & ~a4298;
assign a4304 = ~a4302 & ~l118;
assign a4308 = ~a924 & l118;
assign a4310 = ~a3738 & a1390;
assign a4312 = a1394 & a810;
assign a4314 = a1402 & a1230;
assign a4316 = a3738 & a1406;
assign a4318 = ~a1406 & ~a810;
assign a4320 = ~a4318 & ~a4316;
assign a4322 = ~a4320 & ~a1402;
assign a4324 = ~a4322 & ~a4314;
assign a4326 = ~a4324 & ~a1398;
assign a4328 = a1398 & a1306;
assign a4330 = ~a4328 & ~a4326;
assign a4332 = ~a4330 & ~a1394;
assign a4334 = ~a4332 & ~a4312;
assign a4336 = ~a4334 & ~a1390;
assign a4338 = ~a4336 & ~a4310;
assign a4340 = ~a4338 & ~l118;
assign a4344 = a4204 & a4198;
assign a4346 = a4208 & a3896;
assign a4348 = ~a4346 & ~a4344;
assign a4350 = a4348 & a804;
assign a4352 = a3798 & a3782;
assign a4354 = ~l382 & l102;
assign a4356 = a766 & a720;
assign a4358 = a768 & a744;
assign a4360 = ~a4358 & ~a4356;
assign a4362 = ~a4360 & a526;
assign a4364 = ~a4362 & ~a758;
assign a4366 = a4364 & a528;
assign a4368 = a4366 & ~l102;
assign a4370 = ~a4368 & ~a4354;
assign a4372 = a4370 & ~a3622;
assign a4374 = a4372 & ~l384;
assign a4376 = a4374 & a3752;
assign a4378 = a4376 & a4352;
assign a4380 = a4378 & ~a4350;
assign a4382 = ~l184 & l102;
assign a4384 = ~a528 & ~l102;
assign a4386 = ~a4384 & ~a4382;
assign a4388 = ~a4386 & ~a3812;
assign a4392 = a4236 & a4198;
assign a4394 = a4238 & a3896;
assign a4396 = ~a4394 & ~a4392;
assign a4398 = ~a4396 & ~a3622;
assign a4400 = ~a4398 & a796;
assign a4402 = a4400 & ~a4234;
assign a4406 = ~a3798 & a3782;
assign a4408 = a4406 & a3752;
assign a4410 = ~a824 & ~a802;
assign a4412 = ~a924 & ~a794;
assign a4414 = ~a810 & a794;
assign a4416 = ~a4414 & ~a4412;
assign a4418 = ~a4416 & a802;
assign a4420 = ~a4418 & ~a4410;
assign a4422 = ~a850 & ~a802;
assign a4424 = ~a952 & ~a794;
assign a4426 = ~a838 & a794;
assign a4428 = ~a4426 & ~a4424;
assign a4430 = ~a4428 & a802;
assign a4432 = ~a4430 & ~a4422;
assign a4434 = a4432 & a4420;
assign a4436 = a4434 & ~a4408;
assign a4438 = a4420 & ~a3752;
assign a4440 = ~a4420 & a3752;
assign a4442 = ~a890 & ~a802;
assign a4444 = ~a974 & ~a794;
assign a4446 = ~a870 & a794;
assign a4448 = ~a4446 & ~a4444;
assign a4450 = ~a4448 & a802;
assign a4452 = ~a4450 & ~a4442;
assign a4454 = ~a4452 & ~a3798;
assign a4456 = ~a4432 & a3782;
assign a4458 = ~a4456 & ~a4454;
assign a4460 = a4432 & ~a3782;
assign a4462 = ~a4460 & ~a4458;
assign a4464 = ~a4462 & ~a4440;
assign a4466 = ~a4464 & ~a4438;
assign a4468 = ~a4434 & a4408;
assign a4470 = ~a4468 & a4466;
assign a4472 = ~a4470 & ~a4436;
assign a4474 = a4472 & a4404;
assign a4476 = ~a4474 & ~a4378;
assign a4478 = a4476 & ~a1008;
assign a4482 = ~a3798 & ~a3782;
assign a4484 = a4482 & a4376;
assign a4486 = a4484 & ~a4350;
assign a4488 = a3782 & a3752;
assign a4490 = ~a4452 & ~a4432;
assign a4492 = ~a4490 & a4420;
assign a4494 = a4492 & ~a4488;
assign a4496 = ~a4492 & a4488;
assign a4498 = ~a4496 & a4466;
assign a4500 = ~a4498 & ~a4494;
assign a4502 = a4500 & a4404;
assign a4504 = ~a4502 & ~a4484;
assign a4506 = a4504 & ~a1022;
assign a4510 = a3798 & ~a3782;
assign a4512 = a4510 & a4376;
assign a4514 = a4512 & ~a4350;
assign a4516 = ~a4510 & a3752;
assign a4518 = ~a4516 & a4420;
assign a4520 = ~a4518 & ~a4466;
assign a4522 = ~a4510 & a4440;
assign a4524 = ~a4522 & ~a4520;
assign a4526 = ~a4524 & a4404;
assign a4528 = ~a4526 & ~a4512;
assign a4530 = a4528 & ~a1036;
assign a4534 = a4374 & ~a3752;
assign a4536 = a4534 & a4406;
assign a4538 = a4536 & ~a4350;
assign a4540 = a4452 & ~a4420;
assign a4542 = a4540 & a4432;
assign a4544 = ~a4462 & ~a4438;
assign a4546 = ~a4544 & ~a4440;
assign a4548 = ~a4546 & ~a4542;
assign a4550 = a4548 & a4404;
assign a4552 = ~a4550 & ~a4536;
assign a4554 = a4552 & ~a1050;
assign a4558 = a4534 & a4352;
assign a4560 = a4558 & ~a4350;
assign a4562 = ~a4406 & ~a3752;
assign a4564 = ~a4432 & ~a4420;
assign a4566 = ~a4564 & a4562;
assign a4568 = ~a4566 & ~a4466;
assign a4570 = a4564 & ~a4562;
assign a4572 = ~a4570 & ~a4568;
assign a4574 = ~a4572 & a4404;
assign a4576 = ~a4574 & ~a4558;
assign a4578 = a4576 & l140;
assign a4580 = ~a4578 & ~a4560;
assign a4582 = a4534 & a4482;
assign a4584 = a4582 & ~a4350;
assign a4586 = ~a3782 & ~a3752;
assign a4588 = a4490 & ~a4420;
assign a4590 = ~a4588 & a4586;
assign a4592 = ~a4590 & ~a4466;
assign a4594 = a4588 & ~a4586;
assign a4596 = ~a4594 & ~a4592;
assign a4598 = ~a4596 & a4404;
assign a4600 = ~a4598 & ~a4582;
assign a4602 = a4600 & l142;
assign a4604 = ~a4602 & ~a4584;
assign a4606 = a4510 & ~a3752;
assign a4608 = a4606 & a4374;
assign a4610 = a4608 & ~a4350;
assign a4612 = ~a4466 & a4404;
assign a4614 = a4612 & ~a4606;
assign a4616 = ~a4614 & ~a4608;
assign a4618 = a4616 & l144;
assign a4620 = ~a4618 & ~a4610;
assign a4622 = a4408 & a4374;
assign a4624 = a4622 & ~a4350;
assign a4626 = a4452 & a4434;
assign a4628 = ~a4626 & a4612;
assign a4630 = ~a4628 & ~a4622;
assign a4632 = a4630 & l146;
assign a4634 = ~a4632 & ~a4624;
assign a4636 = a4212 & ~a824;
assign a4638 = a4190 & a4178;
assign a4640 = a4638 & a3738;
assign a4642 = ~a4178 & ~a4170;
assign a4644 = a4642 & a1306;
assign a4646 = ~a4644 & ~a4640;
assign a4648 = ~a4178 & a4170;
assign a4650 = a4648 & a1230;
assign a4652 = ~a4190 & a4170;
assign a4654 = a4652 & a810;
assign a4656 = ~a4654 & ~a4650;
assign a4658 = a4656 & a4646;
assign a4660 = ~a4658 & a4206;
assign a4662 = a4122 & a1306;
assign a4664 = a4146 & ~a810;
assign a4666 = ~a4664 & ~a4662;
assign a4668 = a4144 & ~a3876;
assign a4670 = a4668 & a3738;
assign a4672 = a4130 & a1230;
assign a4674 = a3828 & a810;
assign a4676 = ~a4674 & ~a4672;
assign a4678 = a4676 & ~a4670;
assign a4680 = a4678 & a4666;
assign a4682 = ~a4680 & a4210;
assign a4684 = ~a4682 & ~a4660;
assign a4688 = a4212 & ~a850;
assign a4690 = a4638 & a3766;
assign a4692 = a4648 & a838;
assign a4694 = ~a4692 & ~a4690;
assign a4696 = a4652 & ~a838;
assign a4698 = a4642 & ~a3766;
assign a4700 = ~a4698 & ~a4696;
assign a4702 = a4700 & a4694;
assign a4704 = ~a4702 & a4206;
assign a4706 = a4130 & a838;
assign a4708 = a4668 & a3766;
assign a4710 = ~a4708 & ~a4706;
assign a4712 = a4122 & ~a3766;
assign a4714 = a3876 & ~a3848;
assign a4716 = a4714 & ~a838;
assign a4718 = ~a4716 & ~a4712;
assign a4720 = a4718 & a4710;
assign a4722 = ~a4720 & a4210;
assign a4724 = ~a4722 & ~a4704;
assign a4728 = a4212 & ~a890;
assign a4730 = ~a4170 & ~a870;
assign a4732 = ~a4638 & ~a870;
assign a4734 = a4190 & ~a4170;
assign a4736 = ~a4734 & ~a4732;
assign a4738 = ~a4736 & ~a4730;
assign a4740 = a4738 & a4206;
assign a4742 = a3876 & a870;
assign a4744 = ~a3876 & ~a870;
assign a4746 = ~a4744 & ~a4742;
assign a4748 = a4746 & a3598;
assign a4750 = a4748 & a4210;
assign a4752 = ~a4750 & ~a4740;
assign a4756 = a4248 & ~a924;
assign a4758 = ~a4606 & ~a4516;
assign a4760 = a4758 & a4244;
assign a4762 = ~a4658 & a4236;
assign a4764 = ~a4680 & a4238;
assign a4766 = ~a824 & a762;
assign a4768 = ~a4766 & ~a4764;
assign a4770 = a4768 & ~a4762;
assign a4772 = a4770 & ~a4760;
assign a4776 = a4248 & ~a952;
assign a4778 = ~a4482 & ~a4352;
assign a4780 = ~a4778 & a4244;
assign a4782 = ~a4702 & a4236;
assign a4784 = ~a4720 & a4238;
assign a4786 = ~a850 & a762;
assign a4788 = ~a4786 & ~a4784;
assign a4790 = a4788 & ~a4782;
assign a4792 = a4790 & ~a4780;
assign a4796 = a4248 & ~a974;
assign a4798 = a4244 & ~a3798;
assign a4800 = a4738 & a4236;
assign a4802 = a4748 & a4238;
assign a4804 = ~a890 & a762;
assign a4806 = ~a4804 & ~a4802;
assign a4808 = a4806 & ~a4800;
assign a4810 = a4808 & ~a4798;
assign a4814 = l360 & l118;
assign a4816 = a3736 & l162;
assign a4818 = ~a3736 & ~l162;
assign a4820 = ~a4818 & ~a4816;
assign a4822 = ~a4820 & a1390;
assign a4824 = a810 & l162;
assign a4826 = ~a810 & ~l162;
assign a4828 = ~a4826 & ~a4824;
assign a4830 = ~a4828 & a1394;
assign a4832 = ~a1064 & l162;
assign a4834 = a1064 & ~l162;
assign a4836 = ~a4834 & ~a4832;
assign a4838 = ~a4836 & a1402;
assign a4840 = ~a3734 & l162;
assign a4842 = a3734 & ~l162;
assign a4844 = ~a4842 & ~a4840;
assign a4846 = ~a4844 & a1406;
assign a4848 = ~a1406 & l162;
assign a4850 = ~a4848 & ~a4846;
assign a4852 = ~a4850 & ~a1402;
assign a4854 = ~a4852 & ~a4838;
assign a4856 = ~a4854 & ~a1398;
assign a4858 = ~a1304 & l162;
assign a4860 = a1304 & ~l162;
assign a4862 = ~a4860 & ~a4858;
assign a4864 = ~a4862 & a1398;
assign a4866 = ~a4864 & ~a4856;
assign a4868 = ~a4866 & ~a1394;
assign a4870 = ~a4868 & ~a4830;
assign a4872 = ~a4870 & ~a1390;
assign a4874 = ~a4872 & ~a4822;
assign a4876 = ~a4874 & ~l118;
assign a4878 = ~a4876 & ~a4814;
assign a4880 = ~a4828 & a3718;
assign a4882 = ~a4862 & a3722;
assign a4884 = ~a4836 & a3726;
assign a4886 = ~a4844 & a3732;
assign a4888 = a3742 & l162;
assign a4890 = ~a4888 & ~a4886;
assign a4892 = a4890 & ~a4884;
assign a4894 = a4892 & ~a4882;
assign a4896 = a4894 & ~a4880;
assign a4898 = ~l186 & l102;
assign a4900 = ~a4364 & a528;
assign a4902 = a4900 & ~l102;
assign a4904 = ~a4902 & ~a4898;
assign a4906 = a4896 & l164;
assign a4908 = ~a4896 & ~l164;
assign a4910 = ~a4908 & ~a4906;
assign a4912 = ~l170 & l102;
assign a4914 = a4900 & a536;
assign a4916 = a4914 & ~l102;
assign a4918 = ~a4916 & ~a4912;
assign a4920 = a4918 & ~a3752;
assign a4922 = ~l166 & l102;
assign a4924 = a4900 & a562;
assign a4926 = a4924 & ~l102;
assign a4928 = ~a4926 & ~a4922;
assign a4930 = a4928 & a3798;
assign a4932 = ~l168 & l102;
assign a4934 = a4900 & a546;
assign a4936 = a4934 & ~l102;
assign a4938 = ~a4936 & ~a4932;
assign a4940 = a4938 & ~a3782;
assign a4942 = ~a4940 & ~a4930;
assign a4944 = ~a4938 & a3782;
assign a4946 = ~a4918 & a3752;
assign a4948 = ~a4946 & ~a4944;
assign a4950 = a4948 & ~a4942;
assign a4952 = ~a4950 & ~a4920;
assign a4954 = a4952 & a4910;
assign a4956 = ~a4952 & ~a4910;
assign a4958 = ~a4956 & ~a4954;
assign a4960 = a4958 & ~a4904;
assign a4962 = ~a4960 & ~a4402;
assign a4964 = a4962 & a4390;
assign a4966 = a4964 & ~a4896;
assign a4968 = ~a4964 & l164;
assign a4970 = ~a4968 & ~a4966;
assign a4972 = a4964 & a3798;
assign a4974 = ~a4964 & ~a4928;
assign a4978 = a4964 & ~a3782;
assign a4980 = ~a4964 & ~a4938;
assign a4984 = ~a4964 & ~a4918;
assign a4986 = a4964 & ~a3752;
assign a4990 = ~a3808 & l176;
assign a4992 = ~a4990 & ~l296;
assign a4994 = ~a4390 & ~a4386;
assign a4998 = ~a4928 & ~a3798;
assign a5000 = a4948 & ~a4920;
assign a5002 = a5000 & ~a4998;
assign a5004 = a5002 & a4942;
assign a5006 = ~a4202 & a3902;
assign a5008 = ~a5006 & a5004;
assign a5010 = ~a5008 & ~a4958;
assign a5012 = a5010 & a4404;
assign a5014 = ~a5012 & ~a4904;
assign a5018 = ~l192 & l102;
assign a5020 = a758 & ~l102;
assign a5022 = ~a5020 & ~a5018;
assign a5026 = ~l194 & l102;
assign a5028 = a758 & ~l102;
assign a5030 = ~a5028 & ~a5026;
assign a5034 = ~l196 & l102;
assign a5036 = a758 & ~l102;
assign a5038 = ~a5036 & ~a5034;
assign a5042 = ~l198 & l102;
assign a5044 = a758 & ~l102;
assign a5046 = ~a5044 & ~a5042;
assign a5050 = ~a4234 & ~l200;
assign a5054 = ~l212 & l210;
assign a5056 = ~l214 & l102;
assign a5058 = ~a528 & ~l102;
assign a5062 = ~a5060 & ~l216;
assign a5064 = ~a5060 & ~l218;
assign a5068 = ~a5066 & ~a4390;
assign a5070 = ~l220 & ~l218;
assign a5072 = a5070 & a5068;
assign a5074 = a5072 & a5062;
assign a5076 = ~a5074 & l222;
assign a5080 = ~a5078 & l208;
assign a5082 = ~a5054 & l222;
assign a5084 = a5082 & ~l220;
assign a5086 = ~a5068 & ~l216;
assign a5088 = a5086 & a5084;
assign a5090 = a5088 & a3798;
assign a5092 = a5082 & ~a5070;
assign a5094 = a5092 & l224;
assign a5096 = ~l226 & l102;
assign a5098 = ~a562 & ~l102;
assign a5102 = a5084 & ~a5062;
assign a5104 = a5102 & a5100;
assign a5106 = ~a5104 & ~a5094;
assign a5108 = a5106 & ~a5090;
assign a5110 = a5108 & ~a5080;
assign a5112 = ~a5076 & ~l210;
assign a5116 = ~l228 & l102;
assign a5118 = a758 & ~l102;
assign a5120 = ~a5118 & ~a5116;
assign a5122 = ~l230 & l102;
assign a5124 = ~a4362 & ~l102;
assign a5126 = ~a5124 & ~a5122;
assign a5128 = ~a5126 & a5120;
assign a5130 = ~a3622 & a804;
assign a5132 = a4198 & a4108;
assign a5134 = a3896 & a3600;
assign a5136 = ~a5134 & ~a5132;
assign a5138 = ~a5136 & a5130;
assign a5140 = ~a5138 & a802;
assign a5142 = a5140 & a794;
assign a5144 = ~a5142 & a5066;
assign a5148 = a790 & ~a788;
assign a5150 = a5148 & a4248;
assign a5152 = a5150 & a786;
assign a5158 = ~l242 & l102;
assign a5160 = ~a726 & ~a516;
assign a5162 = a5160 & ~l102;
assign a5164 = ~a5162 & ~a5158;
assign a5166 = a4108 & ~a3600;
assign a5168 = a5166 & ~l244;
assign a5170 = a3600 & ~l244;
assign a5172 = ~l246 & l102;
assign a5174 = ~a726 & a516;
assign a5176 = a5174 & i40;
assign a5178 = a726 & i42;
assign a5180 = ~a5178 & ~a5176;
assign a5182 = ~a5180 & ~l102;
assign a5184 = ~a5182 & ~a5172;
assign a5186 = a5184 & ~a5170;
assign a5188 = a5186 & ~a5168;
assign a5190 = ~l248 & l102;
assign a5192 = a726 & ~i42;
assign a5194 = a5174 & ~i40;
assign a5196 = ~a5194 & ~a5192;
assign a5198 = ~a5196 & ~l102;
assign a5200 = ~a5198 & ~a5190;
assign a5202 = a5200 & ~a762;
assign a5204 = a5202 & ~a5188;
assign a5208 = ~a5126 & l216;
assign a5210 = ~a5208 & ~l240;
assign a5214 = a5188 & ~a5164;
assign a5218 = ~l252 & l102;
assign a5220 = a5196 & ~a758;
assign a5222 = ~a5220 & ~l102;
assign a5224 = ~a5222 & ~a5218;
assign a5226 = a5224 & a5168;
assign a5228 = a5226 & i68;
assign a5230 = a5224 & a5170;
assign a5232 = a5230 & i86;
assign a5236 = ~l250 & l102;
assign a5238 = ~a5160 & ~l102;
assign a5240 = ~a5238 & ~a5236;
assign a5242 = a5230 & ~i86;
assign a5244 = a5226 & ~i68;
assign a5246 = ~a5244 & ~a5242;
assign a5248 = ~a5246 & a5240;
assign a5250 = ~l254 & l102;
assign a5252 = a720 & a516;
assign a5254 = ~a5252 & a528;
assign a5256 = a5254 & ~a1000;
assign a5258 = ~a5256 & ~l102;
assign a5260 = ~a5258 & ~a5250;
assign a5264 = a5262 & ~a4234;
assign a5266 = ~l256 & l102;
assign a5268 = a5252 & i40;
assign a5270 = a5268 & ~a4358;
assign a5272 = a1000 & i42;
assign a5274 = ~a5272 & ~a5270;
assign a5276 = ~a5274 & a528;
assign a5278 = ~a5276 & ~l102;
assign a5280 = ~a5278 & ~a5266;
assign a5284 = ~l258 & l102;
assign a5286 = ~a5220 & ~l102;
assign a5288 = ~a5286 & ~a5284;
assign a5290 = ~l270 & ~l268;
assign a5292 = a5290 & ~l266;
assign a5294 = a5292 & ~l264;
assign a5296 = a5294 & ~l262;
assign a5298 = a5296 & ~l260;
assign a5300 = a5298 & a5288;
assign a5304 = a3632 & a792;
assign a5308 = ~a5306 & a794;
assign a5310 = a5136 & a802;
assign a5314 = a5134 & a4250;
assign a5316 = ~a5314 & i68;
assign a5318 = a5316 & a5132;
assign a5320 = a5134 & i86;
assign a5322 = ~a5320 & ~a5318;
assign a5324 = a5322 & a802;
assign a5326 = ~a5324 & ~a762;
assign a5330 = ~a5078 & l278;
assign a5332 = a5088 & ~a3782;
assign a5334 = a5092 & l280;
assign a5336 = ~l282 & l102;
assign a5338 = a546 & ~l102;
assign a5340 = ~a5338 & ~a5336;
assign a5342 = ~a5340 & a5102;
assign a5344 = ~a5342 & ~a5334;
assign a5346 = a5344 & ~a5332;
assign a5348 = a5346 & ~a5330;
assign a5350 = ~a5078 & l290;
assign a5352 = a5088 & ~a3752;
assign a5354 = a5092 & l292;
assign a5356 = ~l294 & l102;
assign a5358 = a536 & ~l102;
assign a5360 = ~a5358 & ~a5356;
assign a5362 = ~a5360 & a5102;
assign a5364 = ~a5362 & ~a5354;
assign a5366 = a5364 & ~a5352;
assign a5368 = a5366 & ~a5350;
assign a5370 = ~l322 & l102;
assign a5372 = ~a5160 & i90;
assign a5374 = ~a5372 & ~l102;
assign a5378 = ~a4108 & ~a3600;
assign a5380 = ~l326 & ~l324;
assign a5382 = ~l330 & ~l328;
assign a5384 = a5382 & a5380;
assign a5388 = ~l332 & l102;
assign a5390 = a5160 & ~l102;
assign a5394 = ~a5392 & ~l330;
assign a5396 = a5394 & ~a5386;
assign a5400 = ~l336 & l102;
assign a5402 = a526 & ~i96;
assign a5404 = a5402 & i94;
assign a5406 = a5404 & a528;
assign a5408 = a5406 & ~l102;
assign a5410 = ~a5408 & ~a5400;
assign a5412 = ~l334 & l102;
assign a5414 = ~a5404 & ~l102;
assign a5416 = ~a5414 & ~a5412;
assign a5418 = ~a5416 & ~l338;
assign a5420 = a5418 & ~i98;
assign a5422 = ~a3622 & a788;
assign a5424 = ~l340 & l102;
assign a5426 = a526 & i96;
assign a5428 = a5426 & ~l102;
assign a5430 = ~a5428 & ~a5424;
assign a5432 = a5430 & ~l174;
assign a5434 = a5432 & ~i64;
assign a5436 = a5434 & a5422;
assign a5438 = a5436 & a5420;
assign a5440 = a5438 & ~a5306;
assign a5442 = ~a5440 & a5410;
assign a5444 = ~l342 & l102;
assign a5446 = a526 & i94;
assign a5448 = ~a5446 & a5402;
assign a5450 = a5448 & a528;
assign a5452 = a5450 & ~l102;
assign a5454 = ~a5452 & ~a5444;
assign a5456 = a5454 & ~a5442;
assign a5458 = a5456 & l338;
assign a5460 = ~a5458 & a5382;
assign a5464 = a5462 & ~l324;
assign a5466 = ~a5464 & ~l354;
assign a5468 = a5456 & a5416;
assign a5470 = ~l344 & l102;
assign a5472 = ~a5450 & ~l102;
assign a5474 = ~a5472 & ~a5470;
assign a5476 = ~a5474 & ~a5468;
assign a5480 = ~l346 & l102;
assign a5482 = a528 & ~l102;
assign a5484 = ~a5482 & ~a5480;
assign a5486 = ~a5484 & ~a5430;
assign a5488 = a5478 & ~a5306;
assign a5492 = ~a5434 & a5422;
assign a5494 = ~a5454 & ~l118;
assign a5500 = ~l350 & l102;
assign a5502 = ~a1002 & a526;
assign a5504 = a5502 & ~l102;
assign a5506 = ~a5504 & ~a5500;
assign a5508 = a786 & ~l120;
assign a5512 = ~a5464 & ~l356;
assign a5514 = a4248 & l360;
assign a5516 = ~a4896 & ~a4606;
assign a5518 = a4896 & a4606;
assign a5520 = ~a5518 & ~a5516;
assign a5522 = ~a5520 & a4244;
assign a5524 = ~a4844 & a4638;
assign a5526 = ~a4862 & a4642;
assign a5528 = ~a5526 & ~a5524;
assign a5530 = ~a4836 & a4648;
assign a5532 = ~a4828 & a4652;
assign a5534 = ~a5532 & ~a5530;
assign a5536 = a5534 & a5528;
assign a5538 = ~a5536 & a4236;
assign a5540 = ~a4862 & a4122;
assign a5542 = ~a4844 & a4668;
assign a5544 = ~a5542 & ~a5540;
assign a5546 = a4146 & l162;
assign a5548 = ~a4836 & a4130;
assign a5550 = ~a4828 & a3828;
assign a5552 = ~a5550 & ~a5548;
assign a5554 = a5552 & ~a5546;
assign a5556 = a5554 & a5544;
assign a5558 = ~a5556 & a4238;
assign a5560 = a762 & l362;
assign a5562 = ~a5560 & ~a5558;
assign a5564 = a5562 & ~a5538;
assign a5566 = a5564 & ~a5522;
assign a5568 = a5566 & ~a5514;
assign a5570 = a4212 & l362;
assign a5572 = ~a5536 & a4206;
assign a5574 = ~a5556 & a4210;
assign a5576 = ~a5574 & ~a5572;
assign a5578 = a5576 & ~a5570;
assign a5580 = ~l378 & l102;
assign a5582 = ~a770 & ~l102;
assign a5584 = ~a5582 & ~a5580;
assign a5586 = ~l380 & l102;
assign a5588 = a770 & ~a758;
assign a5590 = ~a5588 & ~l102;
assign a5592 = ~a5590 & ~a5586;
assign a5596 = ~a5280 & ~a5260;
assign a5598 = a4240 & ~a4234;
assign a5600 = a5598 & a5596;
assign a5604 = ~a4404 & ~l388;
assign a5608 = ~l386 & l102;
assign a5610 = ~a4366 & ~l102;
assign a5614 = ~l392 & l102;
assign a5616 = a4366 & ~l102;
assign a5618 = ~a5616 & ~a5614;
assign a5620 = ~l394 & l102;
assign a5622 = a4366 & ~l102;
assign a5624 = ~a5622 & ~a5620;
assign a5626 = a5624 & ~a4404;
assign a5632 = ~l398 & l102;
assign a5634 = a4366 & ~l102;
assign a5636 = ~a5634 & ~a5632;
assign a5638 = a5636 & ~l384;
assign a5642 = ~a5612 & ~l384;
assign a5644 = ~a4904 & ~a4390;
assign a5646 = a5644 & a5004;
assign a5648 = a5646 & a4910;
assign a5650 = a5648 & a5130;
assign p0 = a5650;

assert property (~p0);

endmodule
