module m6s12 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58;

output p0;

wire a1274,na1300,c1,a1302,na1406,na1486,na1506,na1530,na1550,na1570,na1670,na1728,na1740,na1764,na1770,
na1800,na1810,na1820,na1830,na1840,na1850,na1860,na1870,na1880,na1890,na1900,na1924,na1928,na1946,na1956,
na1966,na2014,a2018,na2024,a2042,na2060,na2066,na2078,na2090,na2102,a2112,na2118,na2136,na2154,na2168,
na2186,na2206,a2224,na2234,na2240,na2252,na2264,na2278,na2296,na2308,na2326,na2338,na2356,na2374,na2380,
na2418,na2424,na2438,na2454,na2470,a2490,na2498,na2464,nl1064,na2510,na2614,a2634,na2698,a2484,na2722,
na2734,na2746,na2758,na2770,na2782,na2794,na2806,na2818,na2830,na2842,na2854,na2866,na2878,na2890,na2902,
na2914,na2934,na2946,na2958,na2970,na2982,na2992,na3014,na3044,na3056,na2692,na3050,na3076,na3098,na3110,
na3130,na3038,na3142,na3124,na3136,na3154,na3104,na3148,na3188,na3208,na3232,na3258,na3276,na3296,na3322,
na3344,na3364,na3384,na3406,na3424,na3442,na3460,na3480,na3502,na3522,na3542,na3560,na3578,na3596,na3616,
na3634,na3652,na3670,na3688,na3720,na3742,na3766,na3092,na3794,na3814,na3844,na3878,na3760,na3890,na3910,
na3872,na3924,na3904,na3918,na3884,a3936,a3954,a3966,na3984,a3996,a4008,a4020,a4032,na3838,na4026,
na4014,na4002,na3990,na3978,na3960,a3948,na3930,na3808,na4050,na4068,na4080,na4094,na4106,na3788,na4100,
na4088,a4074,na4140,na4158,na4190,na4208,na4238,na4134,na4256,na4286,na4232,na4304,na4334,na4280,na4352,
na4366,na4396,na4328,na4414,na4444,na4390,na4474,na4438,na4504,na4468,na4510,na4540,na4498,na4546,na4576,
na4534,na4606,na4570,na4624,na4654,na4600,na4672,na4702,na4648,na4720,na4750,na4696,na4768,na4798,na4744,
na4816,na4836,na4866,na4792,na4884,a4902,na4932,na4860,a4950,na4976,na4926,na4994,na5018,na4970,na5036,
na5060,na5012,na5078,na5102,na5054,na5126,na5096,na5150,na5120,na5168,na5192,na5144,na5210,na5186,na5228,
na5204,na5246,na5222,na5264,na5240,na5282,na5258,na5300,na5276,na5318,na5294,na5336,na5312,na5362,na5330,
na5366,na5390,na5356,na5394,na5418,na5384,na5422,na5446,na5412,na5450,na5474,na5440,na5480,na5504,na5468,
na5508,na5532,na5498,na5536,na5560,na5526,na5564,na5588,na5554,na5592,na5616,na5582,na5620,na5644,na5610,
na5648,na5672,na5638,na5676,na5700,na5666,na5704,na5728,na5694,na5732,na5750,na5722,na5768,na5744,na5786,
na5762,na5804,na5780,na5822,na5798,na5840,na5816,na5858,na5834,na5876,na5852,na5894,na5870,na5912,na5888,
na5930,na5906,na5948,na5924,na5966,na5942,na5984,na5960,na6002,na5978,na6020,na5996,na6038,na6014,na6058,
na6032,na6074,na6052,na6068,na6170,na6194,na6214,na6236,na6256,na6276,na6296,na6316,na6350,na6370,na6390,
na6410,na6430,na6450,na6470,na6490,na6516,na6524,na6310,na6528,na6540,na6534,na6554,na6566,na6578,na6510,
nl814,na6572,z0,na6560,na6548,na6484,na6464,na6444,na6424,na6404,na6384,na6364,na6344,na6290,na6270,
na6250,na6230,na6208,na6188,na6606,na6626,na6632,na6600,na6646,na6666,na6620,na6660,na6640,na6678,na6672,
na6684,na6702,na5162,a6708,na6696,na6704,na5072,na5030,na4988,a4944,a4896,na4878,na4830,na4810,na4762,
na4714,na4666,na4618,na4408,na4346,na4298,na4250,na4202,na6724,na6870,na4184,na6864,na6718,na4152,na6888,
na6908,na6926,na6944,na6970,na4062,na6964,na6938,na6920,na6902,na6882,na4044,na3736,na3714,na3682,na3664,
na3646,na3628,na3610,na3590,na3572,na3554,na3536,na3516,na3496,na3474,na3454,na3436,na3418,na3400,na3378,
na3358,na3338,na3316,na3290,na3270,na3252,na3226,na3202,na3182,na3070,na3008,a2986,na2976,na2964,na2952,
na2940,na2928,na2908,na2896,na2884,na2872,na2860,na2848,na2836,na2824,na2812,na2800,na2788,na2776,na2764,
na2752,na2740,na2728,na2716,a2628,na2608,na2504,z1,na2448,na2432,na6990,na7008,na7026,na2412,na7020,
na7002,na6984,na2368,na2350,na2332,na2320,na7032,na2290,na2270,na2258,na2246,a2218,na7036,na7052,na7058,
na7046,na7070,na7074,a7064,na2180,na2162,na2148,na2096,na2084,na2072,na2054,na2008,na7086,na7106,na7118,
na7140,na7134,na7112,na7100,na7080,na1940,na1758,na1564,na1544,na1524,na1500,na1480,a1168,a1170,a1172,
a1174,a1176,a1178,a1180,a1182,a1184,a1186,a1188,a1190,a1192,a1194,a1196,a1198,a1200,a1202,
a1204,a1206,a1208,a1210,a1212,a1214,a1216,a1218,a1220,a1222,a1224,a1226,a1228,a1230,a1232,
a1234,a1236,a1238,a1240,a1242,a1244,a1246,a1248,a1250,a1252,a1254,a1256,a1258,a1260,a1262,
a1264,a1266,a1268,a1270,a1272,a1276,a1278,a1280,a1282,a1284,a1286,a1288,a1290,a1292,a1294,
a1296,a1298,a1300,a1304,a1306,a1308,a1310,a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,
a1328,a1330,a1332,a1334,a1336,a1338,a1340,a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,
a1358,a1360,a1362,a1364,a1366,a1368,a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,
a1388,a1390,a1392,a1394,a1396,a1398,a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,
a1418,a1420,a1422,a1424,a1426,a1428,a1430,a1432,a1434,a1436,a1438,a1440,a1442,a1444,a1446,
a1448,a1450,a1452,a1454,a1456,a1458,a1460,a1462,a1464,a1466,a1468,a1470,a1472,a1474,a1476,
a1478,a1480,a1482,a1484,a1486,a1488,a1490,a1492,a1494,a1496,a1498,a1500,a1502,a1504,a1506,
a1508,a1510,a1512,a1514,a1516,a1518,a1520,a1522,a1524,a1526,a1528,a1530,a1532,a1534,a1536,
a1538,a1540,a1542,a1544,a1546,a1548,a1550,a1552,a1554,a1556,a1558,a1560,a1562,a1564,a1566,
a1568,a1570,a1572,a1574,a1576,a1578,a1580,a1582,a1584,a1586,a1588,a1590,a1592,a1594,a1596,
a1598,a1600,a1602,a1604,a1606,a1608,a1610,a1612,a1614,a1616,a1618,a1620,a1622,a1624,a1626,
a1628,a1630,a1632,a1634,a1636,a1638,a1640,a1642,a1644,a1646,a1648,a1650,a1652,a1654,a1656,
a1658,a1660,a1662,a1664,a1666,a1668,a1670,a1672,a1674,a1676,a1678,a1680,a1682,a1684,a1686,
a1688,a1690,a1692,a1694,a1696,a1698,a1700,a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,
a1718,a1720,a1722,a1724,a1726,a1728,a1730,a1732,a1734,a1736,a1738,a1740,a1742,a1744,a1746,
a1748,a1750,a1752,a1754,a1756,a1758,a1760,a1762,a1764,a1766,a1768,a1770,a1772,a1774,a1776,
a1778,a1780,a1782,a1784,a1786,a1788,a1790,a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,
a1808,a1810,a1812,a1814,a1816,a1818,a1820,a1822,a1824,a1826,a1828,a1830,a1832,a1834,a1836,
a1838,a1840,a1842,a1844,a1846,a1848,a1850,a1852,a1854,a1856,a1858,a1860,a1862,a1864,a1866,
a1868,a1870,a1872,a1874,a1876,a1878,a1880,a1882,a1884,a1886,a1888,a1890,a1892,a1894,a1896,
a1898,a1900,a1902,a1904,a1906,a1908,a1910,a1912,a1914,a1916,a1918,a1920,a1922,a1924,a1926,
a1928,a1930,a1932,a1934,a1936,a1938,a1940,a1942,a1944,a1946,a1948,a1950,a1952,a1954,a1956,
a1958,a1960,a1962,a1964,a1966,a1968,a1970,a1972,a1974,a1976,a1978,a1980,a1982,a1984,a1986,
a1988,a1990,a1992,a1994,a1996,a1998,a2000,a2002,a2004,a2006,a2008,a2010,a2012,a2014,a2016,
a2020,a2022,a2024,a2026,a2028,a2030,a2032,a2034,a2036,a2038,a2040,a2044,a2046,a2048,a2050,
a2052,a2054,a2056,a2058,a2060,a2062,a2064,a2066,a2068,a2070,a2072,a2074,a2076,a2078,a2080,
a2082,a2084,a2086,a2088,a2090,a2092,a2094,a2096,a2098,a2100,a2102,a2104,a2106,a2108,a2110,
a2114,a2116,a2118,a2120,a2122,a2124,a2126,a2128,a2130,a2132,a2134,a2136,a2138,a2140,a2142,
a2144,a2146,a2148,a2150,a2152,a2154,a2156,a2158,a2160,a2162,a2164,a2166,a2168,a2170,a2172,
a2174,a2176,a2178,a2180,a2182,a2184,a2186,a2188,a2190,a2192,a2194,a2196,a2198,a2200,a2202,
a2204,a2206,a2208,a2210,a2212,a2214,a2216,a2220,a2222,a2226,a2228,a2230,a2232,a2234,a2236,
a2238,a2240,a2242,a2244,a2246,a2248,a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,
a2268,a2270,a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,
a2298,a2300,a2302,a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,
a2328,a2330,a2332,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,
a2358,a2360,a2362,a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,
a2388,a2390,a2392,a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,
a2418,a2420,a2422,a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,
a2448,a2450,a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,
a2478,a2480,a2482,a2486,a2488,a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,a2508,a2510,
a2512,a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,a2540,
a2542,a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,
a2572,a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,
a2602,a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2630,a2632,
a2636,a2638,a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,a2662,a2664,
a2666,a2668,a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,a2692,a2694,
a2696,a2698,a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,a2718,a2720,a2722,a2724,
a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,a2752,a2754,
a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,a2782,a2784,
a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,a2810,a2812,a2814,
a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,a2840,a2842,a2844,
a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,a2870,a2872,a2874,
a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,a2900,a2902,a2904,
a2906,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2930,a2932,a2934,
a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,a2960,a2962,a2964,
a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2988,a2990,a2992,a2994,a2996,
a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,a3022,a3024,a3026,
a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,a3048,a3050,a3052,a3054,a3056,
a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,a3078,a3080,a3082,a3084,a3086,
a3088,a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,a3112,a3114,a3116,
a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,a3142,a3144,a3146,
a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,a3172,a3174,a3176,
a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3200,a3202,a3204,a3206,
a3208,a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,a3228,a3230,a3232,a3234,a3236,
a3238,a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,a3262,a3264,a3266,
a3268,a3270,a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,a3288,a3290,a3292,a3294,a3296,
a3298,a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,a3324,a3326,
a3328,a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,a3354,a3356,
a3358,a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3382,a3384,a3386,
a3388,a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,a3408,a3410,a3412,a3414,a3416,
a3418,a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,a3438,a3440,a3442,a3444,a3446,
a3448,a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,a3468,a3470,a3472,a3474,a3476,
a3478,a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,a3498,a3500,a3502,a3504,a3506,
a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,a3528,a3530,a3532,a3534,a3536,
a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,a3558,a3560,a3562,a3564,a3566,
a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,a3588,a3590,a3592,a3594,a3596,
a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,a3618,a3620,a3622,a3624,a3626,
a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3648,a3650,a3652,a3654,a3656,
a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,a3678,a3680,a3682,a3684,a3686,
a3688,a3690,a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,a3712,a3714,a3716,
a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,a3738,a3740,a3742,a3744,a3746,
a3748,a3750,a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,a3768,a3770,a3772,a3774,a3776,
a3778,a3780,a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,a3798,a3800,a3802,a3804,a3806,
a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,a3828,a3830,a3832,a3834,a3836,
a3838,a3840,a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,a3858,a3860,a3862,a3864,a3866,
a3868,a3870,a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,a3888,a3890,a3892,a3894,a3896,
a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,a3918,a3920,a3922,a3924,a3926,
a3928,a3930,a3932,a3934,a3938,a3940,a3942,a3944,a3946,a3950,a3952,a3956,a3958,a3960,a3962,
a3964,a3968,a3970,a3972,a3974,a3976,a3978,a3980,a3982,a3984,a3986,a3988,a3990,a3992,a3994,
a3998,a4000,a4002,a4004,a4006,a4010,a4012,a4014,a4016,a4018,a4022,a4024,a4026,a4028,a4030,
a4034,a4036,a4038,a4040,a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,
a4064,a4066,a4068,a4070,a4072,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,
a4096,a4098,a4100,a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4124,
a4126,a4128,a4130,a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,a4152,a4154,
a4156,a4158,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,a4184,
a4186,a4188,a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,a4214,
a4216,a4218,a4220,a4222,a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,a4244,
a4246,a4248,a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,a4274,
a4276,a4278,a4280,a4282,a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,
a4306,a4308,a4310,a4312,a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,a4334,
a4336,a4338,a4340,a4342,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,
a4366,a4368,a4370,a4372,a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,a4394,
a4396,a4398,a4400,a4402,a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,
a4426,a4428,a4430,a4432,a4434,a4436,a4438,a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,
a4456,a4458,a4460,a4462,a4464,a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4482,a4484,
a4486,a4488,a4490,a4492,a4494,a4496,a4498,a4500,a4502,a4504,a4506,a4508,a4510,a4512,a4514,
a4516,a4518,a4520,a4522,a4524,a4526,a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,
a4546,a4548,a4550,a4552,a4554,a4556,a4558,a4560,a4562,a4564,a4566,a4568,a4570,a4572,a4574,
a4576,a4578,a4580,a4582,a4584,a4586,a4588,a4590,a4592,a4594,a4596,a4598,a4600,a4602,a4604,
a4606,a4608,a4610,a4612,a4614,a4616,a4618,a4620,a4622,a4624,a4626,a4628,a4630,a4632,a4634,
a4636,a4638,a4640,a4642,a4644,a4646,a4648,a4650,a4652,a4654,a4656,a4658,a4660,a4662,a4664,
a4666,a4668,a4670,a4672,a4674,a4676,a4678,a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,
a4696,a4698,a4700,a4702,a4704,a4706,a4708,a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,
a4726,a4728,a4730,a4732,a4734,a4736,a4738,a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,
a4756,a4758,a4760,a4762,a4764,a4766,a4768,a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4784,
a4786,a4788,a4790,a4792,a4794,a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,a4812,a4814,
a4816,a4818,a4820,a4822,a4824,a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,a4844,
a4846,a4848,a4850,a4852,a4854,a4856,a4858,a4860,a4862,a4864,a4866,a4868,a4870,a4872,a4874,
a4876,a4878,a4880,a4882,a4884,a4886,a4888,a4890,a4892,a4894,a4898,a4900,a4904,a4906,a4908,
a4910,a4912,a4914,a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,a4938,
a4940,a4942,a4946,a4948,a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,a4968,a4970,a4972,
a4974,a4976,a4978,a4980,a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,a4998,a5000,a5002,
a5004,a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,a5028,a5030,a5032,
a5034,a5036,a5038,a5040,a5042,a5044,a5046,a5048,a5050,a5052,a5054,a5056,a5058,a5060,a5062,
a5064,a5066,a5068,a5070,a5072,a5074,a5076,a5078,a5080,a5082,a5084,a5086,a5088,a5090,a5092,
a5094,a5096,a5098,a5100,a5102,a5104,a5106,a5108,a5110,a5112,a5114,a5116,a5118,a5120,a5122,
a5124,a5126,a5128,a5130,a5132,a5134,a5136,a5138,a5140,a5142,a5144,a5146,a5148,a5150,a5152,
a5154,a5156,a5158,a5160,a5162,a5164,a5166,a5168,a5170,a5172,a5174,a5176,a5178,a5180,a5182,
a5184,a5186,a5188,a5190,a5192,a5194,a5196,a5198,a5200,a5202,a5204,a5206,a5208,a5210,a5212,
a5214,a5216,a5218,a5220,a5222,a5224,a5226,a5228,a5230,a5232,a5234,a5236,a5238,a5240,a5242,
a5244,a5246,a5248,a5250,a5252,a5254,a5256,a5258,a5260,a5262,a5264,a5266,a5268,a5270,a5272,
a5274,a5276,a5278,a5280,a5282,a5284,a5286,a5288,a5290,a5292,a5294,a5296,a5298,a5300,a5302,
a5304,a5306,a5308,a5310,a5312,a5314,a5316,a5318,a5320,a5322,a5324,a5326,a5328,a5330,a5332,
a5334,a5336,a5338,a5340,a5342,a5344,a5346,a5348,a5350,a5352,a5354,a5356,a5358,a5360,a5362,
a5364,a5366,a5368,a5370,a5372,a5374,a5376,a5378,a5380,a5382,a5384,a5386,a5388,a5390,a5392,
a5394,a5396,a5398,a5400,a5402,a5404,a5406,a5408,a5410,a5412,a5414,a5416,a5418,a5420,a5422,
a5424,a5426,a5428,a5430,a5432,a5434,a5436,a5438,a5440,a5442,a5444,a5446,a5448,a5450,a5452,
a5454,a5456,a5458,a5460,a5462,a5464,a5466,a5468,a5470,a5472,a5474,a5476,a5478,a5480,a5482,
a5484,a5486,a5488,a5490,a5492,a5494,a5496,a5498,a5500,a5502,a5504,a5506,a5508,a5510,a5512,
a5514,a5516,a5518,a5520,a5522,a5524,a5526,a5528,a5530,a5532,a5534,a5536,a5538,a5540,a5542,
a5544,a5546,a5548,a5550,a5552,a5554,a5556,a5558,a5560,a5562,a5564,a5566,a5568,a5570,a5572,
a5574,a5576,a5578,a5580,a5582,a5584,a5586,a5588,a5590,a5592,a5594,a5596,a5598,a5600,a5602,
a5604,a5606,a5608,a5610,a5612,a5614,a5616,a5618,a5620,a5622,a5624,a5626,a5628,a5630,a5632,
a5634,a5636,a5638,a5640,a5642,a5644,a5646,a5648,a5650,a5652,a5654,a5656,a5658,a5660,a5662,
a5664,a5666,a5668,a5670,a5672,a5674,a5676,a5678,a5680,a5682,a5684,a5686,a5688,a5690,a5692,
a5694,a5696,a5698,a5700,a5702,a5704,a5706,a5708,a5710,a5712,a5714,a5716,a5718,a5720,a5722,
a5724,a5726,a5728,a5730,a5732,a5734,a5736,a5738,a5740,a5742,a5744,a5746,a5748,a5750,a5752,
a5754,a5756,a5758,a5760,a5762,a5764,a5766,a5768,a5770,a5772,a5774,a5776,a5778,a5780,a5782,
a5784,a5786,a5788,a5790,a5792,a5794,a5796,a5798,a5800,a5802,a5804,a5806,a5808,a5810,a5812,
a5814,a5816,a5818,a5820,a5822,a5824,a5826,a5828,a5830,a5832,a5834,a5836,a5838,a5840,a5842,
a5844,a5846,a5848,a5850,a5852,a5854,a5856,a5858,a5860,a5862,a5864,a5866,a5868,a5870,a5872,
a5874,a5876,a5878,a5880,a5882,a5884,a5886,a5888,a5890,a5892,a5894,a5896,a5898,a5900,a5902,
a5904,a5906,a5908,a5910,a5912,a5914,a5916,a5918,a5920,a5922,a5924,a5926,a5928,a5930,a5932,
a5934,a5936,a5938,a5940,a5942,a5944,a5946,a5948,a5950,a5952,a5954,a5956,a5958,a5960,a5962,
a5964,a5966,a5968,a5970,a5972,a5974,a5976,a5978,a5980,a5982,a5984,a5986,a5988,a5990,a5992,
a5994,a5996,a5998,a6000,a6002,a6004,a6006,a6008,a6010,a6012,a6014,a6016,a6018,a6020,a6022,
a6024,a6026,a6028,a6030,a6032,a6034,a6036,a6038,a6040,a6042,a6044,a6046,a6048,a6050,a6052,
a6054,a6056,a6058,a6060,a6062,a6064,a6066,a6068,a6070,a6072,a6074,a6076,a6078,a6080,a6082,
a6084,a6086,a6088,a6090,a6092,a6094,a6096,a6098,a6100,a6102,a6104,a6106,a6108,a6110,a6112,
a6114,a6116,a6118,a6120,a6122,a6124,a6126,a6128,a6130,a6132,a6134,a6136,a6138,a6140,a6142,
a6144,a6146,a6148,a6150,a6152,a6154,a6156,a6158,a6160,a6162,a6164,a6166,a6168,a6170,a6172,
a6174,a6176,a6178,a6180,a6182,a6184,a6186,a6188,a6190,a6192,a6194,a6196,a6198,a6200,a6202,
a6204,a6206,a6208,a6210,a6212,a6214,a6216,a6218,a6220,a6222,a6224,a6226,a6228,a6230,a6232,
a6234,a6236,a6238,a6240,a6242,a6244,a6246,a6248,a6250,a6252,a6254,a6256,a6258,a6260,a6262,
a6264,a6266,a6268,a6270,a6272,a6274,a6276,a6278,a6280,a6282,a6284,a6286,a6288,a6290,a6292,
a6294,a6296,a6298,a6300,a6302,a6304,a6306,a6308,a6310,a6312,a6314,a6316,a6318,a6320,a6322,
a6324,a6326,a6328,a6330,a6332,a6334,a6336,a6338,a6340,a6342,a6344,a6346,a6348,a6350,a6352,
a6354,a6356,a6358,a6360,a6362,a6364,a6366,a6368,a6370,a6372,a6374,a6376,a6378,a6380,a6382,
a6384,a6386,a6388,a6390,a6392,a6394,a6396,a6398,a6400,a6402,a6404,a6406,a6408,a6410,a6412,
a6414,a6416,a6418,a6420,a6422,a6424,a6426,a6428,a6430,a6432,a6434,a6436,a6438,a6440,a6442,
a6444,a6446,a6448,a6450,a6452,a6454,a6456,a6458,a6460,a6462,a6464,a6466,a6468,a6470,a6472,
a6474,a6476,a6478,a6480,a6482,a6484,a6486,a6488,a6490,a6492,a6494,a6496,a6498,a6500,a6502,
a6504,a6506,a6508,a6510,a6512,a6514,a6516,a6518,a6520,a6522,a6524,a6526,a6528,a6530,a6532,
a6534,a6536,a6538,a6540,a6542,a6544,a6546,a6548,a6550,a6552,a6554,a6556,a6558,a6560,a6562,
a6564,a6566,a6568,a6570,a6572,a6574,a6576,a6578,a6580,a6582,a6584,a6586,a6588,a6590,a6592,
a6594,a6596,a6598,a6600,a6602,a6604,a6606,a6608,a6610,a6612,a6614,a6616,a6618,a6620,a6622,
a6624,a6626,a6628,a6630,a6632,a6634,a6636,a6638,a6640,a6642,a6644,a6646,a6648,a6650,a6652,
a6654,a6656,a6658,a6660,a6662,a6664,a6666,a6668,a6670,a6672,a6674,a6676,a6678,a6680,a6682,
a6684,a6686,a6688,a6690,a6692,a6694,a6696,a6698,a6700,a6702,a6704,a6706,a6710,a6712,a6714,
a6716,a6718,a6720,a6722,a6724,a6726,a6728,a6730,a6732,a6734,a6736,a6738,a6740,a6742,a6744,
a6746,a6748,a6750,a6752,a6754,a6756,a6758,a6760,a6762,a6764,a6766,a6768,a6770,a6772,a6774,
a6776,a6778,a6780,a6782,a6784,a6786,a6788,a6790,a6792,a6794,a6796,a6798,a6800,a6802,a6804,
a6806,a6808,a6810,a6812,a6814,a6816,a6818,a6820,a6822,a6824,a6826,a6828,a6830,a6832,a6834,
a6836,a6838,a6840,a6842,a6844,a6846,a6848,a6850,a6852,a6854,a6856,a6858,a6860,a6862,a6864,
a6866,a6868,a6870,a6872,a6874,a6876,a6878,a6880,a6882,a6884,a6886,a6888,a6890,a6892,a6894,
a6896,a6898,a6900,a6902,a6904,a6906,a6908,a6910,a6912,a6914,a6916,a6918,a6920,a6922,a6924,
a6926,a6928,a6930,a6932,a6934,a6936,a6938,a6940,a6942,a6944,a6946,a6948,a6950,a6952,a6954,
a6956,a6958,a6960,a6962,a6964,a6966,a6968,a6970,a6972,a6974,a6976,a6978,a6980,a6982,a6984,
a6986,a6988,a6990,a6992,a6994,a6996,a6998,a7000,a7002,a7004,a7006,a7008,a7010,a7012,a7014,
a7016,a7018,a7020,a7022,a7024,a7026,a7028,a7030,a7032,a7034,a7036,a7038,a7040,a7042,a7044,
a7046,a7048,a7050,a7052,a7054,a7056,a7058,a7060,a7062,a7066,a7068,a7070,a7072,a7074,a7076,
a7078,a7080,a7082,a7084,a7086,a7088,a7090,a7092,a7094,a7096,a7098,a7100,a7102,a7104,a7106,
a7108,a7110,a7112,a7114,a7116,a7118,a7120,a7122,a7124,a7126,a7128,a7130,a7132,a7134,a7136,
a7138,a7140,p0;

reg l60,l62,l64,l66,l68,l70,l72,l74,l76,l78,l80,l82,l84,l86,l88,
l90,l92,l94,l96,l98,l100,l102,l104,l106,l108,l110,l112,l114,l116,l118,
l120,l122,l124,l126,l128,l130,l132,l134,l136,l138,l140,l142,l144,l146,l148,
l150,l152,l154,l156,l158,l160,l162,l164,l166,l168,l170,l172,l174,l176,l178,
l180,l182,l184,l186,l188,l190,l192,l194,l196,l198,l200,l202,l204,l206,l208,
l210,l212,l214,l216,l218,l220,l222,l224,l226,l228,l230,l232,l234,l236,l238,
l240,l242,l244,l246,l248,l250,l252,l254,l256,l258,l260,l262,l264,l266,l268,
l270,l272,l274,l276,l278,l280,l282,l284,l286,l288,l290,l292,l294,l296,l298,
l300,l302,l304,l306,l308,l310,l312,l314,l316,l318,l320,l322,l324,l326,l328,
l330,l332,l334,l336,l338,l340,l342,l344,l346,l348,l350,l352,l354,l356,l358,
l360,l362,l364,l366,l368,l370,l372,l374,l376,l378,l380,l382,l384,l386,l388,
l390,l392,l394,l396,l398,l400,l402,l404,l406,l408,l410,l412,l414,l416,l418,
l420,l422,l424,l426,l428,l430,l432,l434,l436,l438,l440,l442,l444,l446,l448,
l450,l452,l454,l456,l458,l460,l462,l464,l466,l468,l470,l472,l474,l476,l478,
l480,l482,l484,l486,l488,l490,l492,l494,l496,l498,l500,l502,l504,l506,l508,
l510,l512,l514,l516,l518,l520,l522,l524,l526,l528,l530,l532,l534,l536,l538,
l540,l542,l544,l546,l548,l550,l552,l554,l556,l558,l560,l562,l564,l566,l568,
l570,l572,l574,l576,l578,l580,l582,l584,l586,l588,l590,l592,l594,l596,l598,
l600,l602,l604,l606,l608,l610,l612,l614,l616,l618,l620,l622,l624,l626,l628,
l630,l632,l634,l636,l638,l640,l642,l644,l646,l648,l650,l652,l654,l656,l658,
l660,l662,l664,l666,l668,l670,l672,l674,l676,l678,l680,l682,l684,l686,l688,
l690,l692,l694,l696,l698,l700,l702,l704,l706,l708,l710,l712,l714,l716,l718,
l720,l722,l724,l726,l728,l730,l732,l734,l736,l738,l740,l742,l744,l746,l748,
l750,l752,l754,l756,l758,l760,l762,l764,l766,l768,l770,l772,l774,l776,l778,
l780,l782,l784,l786,l788,l790,l792,l794,l796,l798,l800,l802,l804,l806,l808,
l810,l812,l814,l816,l818,l820,l822,l824,l826,l828,l830,l832,l834,l836,l838,
l840,l842,l844,l846,l848,l850,l852,l854,l856,l858,l860,l862,l864,l866,l868,
l870,l872,l874,l876,l878,l880,l882,l884,l886,l888,l890,l892,l894,l896,l898,
l900,l902,l904,l906,l908,l910,l912,l914,l916,l918,l920,l922,l924,l926,l928,
l930,l932,l934,l936,l938,l940,l942,l944,l946,l948,l950,l952,l954,l956,l958,
l960,l962,l964,l966,l968,l970,l972,l974,l976,l978,l980,l982,l984,l986,l988,
l990,l992,l994,l996,l998,l1000,l1002,l1004,l1006,l1008,l1010,l1012,l1014,l1016,l1018,
l1020,l1022,l1024,l1026,l1028,l1030,l1032,l1034,l1036,l1038,l1040,l1042,l1044,l1046,l1048,
l1050,l1052,l1054,l1056,l1058,l1060,l1062,l1064,l1066,l1068,l1070,l1072,l1074,l1076,l1078,
l1080,l1082,l1084,l1086,l1088,l1090,l1092,l1094,l1096,l1098,l1100,l1102,l1104,l1106,l1108,
l1110,l1112,l1114,l1116,l1118,l1120,l1122,l1124,l1126,l1128,l1130,l1132,l1134,l1136,l1138,
l1140,l1142,l1144,l1146,l1148,l1150,l1152,l1154,l1156,l1158,l1160,l1162,l1164,l1166;

initial
begin
   l60 = 0;
   l62 = 0;
   l64 = 0;
   l66 = 0;
   l68 = 0;
   l70 = 0;
   l72 = 0;
   l74 = 0;
   l76 = 0;
   l78 = 0;
   l80 = 0;
   l82 = 0;
   l84 = 0;
   l86 = 0;
   l88 = 0;
   l90 = 0;
   l92 = 0;
   l94 = 0;
   l96 = 0;
   l98 = 0;
   l100 = 0;
   l102 = 0;
   l104 = 0;
   l106 = 0;
   l108 = 0;
   l110 = 0;
   l112 = 0;
   l114 = 0;
   l116 = 0;
   l118 = 0;
   l120 = 0;
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
   l392 = 0;
   l394 = 0;
   l396 = 0;
   l398 = 0;
   l400 = 0;
   l402 = 0;
   l404 = 0;
   l406 = 0;
   l408 = 0;
   l410 = 0;
   l412 = 0;
   l414 = 0;
   l416 = 0;
   l418 = 0;
   l420 = 0;
   l422 = 0;
   l424 = 0;
   l426 = 0;
   l428 = 0;
   l430 = 0;
   l432 = 0;
   l434 = 0;
   l436 = 0;
   l438 = 0;
   l440 = 0;
   l442 = 0;
   l444 = 0;
   l446 = 0;
   l448 = 0;
   l450 = 0;
   l452 = 0;
   l454 = 0;
   l456 = 0;
   l458 = 0;
   l460 = 0;
   l462 = 0;
   l464 = 0;
   l466 = 0;
   l468 = 0;
   l470 = 0;
   l472 = 0;
   l474 = 0;
   l476 = 0;
   l478 = 0;
   l480 = 0;
   l482 = 0;
   l484 = 0;
   l486 = 0;
   l488 = 0;
   l490 = 0;
   l492 = 0;
   l494 = 0;
   l496 = 0;
   l498 = 0;
   l500 = 0;
   l502 = 0;
   l504 = 0;
   l506 = 0;
   l508 = 0;
   l510 = 0;
   l512 = 0;
   l514 = 0;
   l516 = 0;
   l518 = 0;
   l520 = 0;
   l522 = 0;
   l524 = 0;
   l526 = 0;
   l528 = 0;
   l530 = 0;
   l532 = 0;
   l534 = 0;
   l536 = 0;
   l538 = 0;
   l540 = 0;
   l542 = 0;
   l544 = 0;
   l546 = 0;
   l548 = 0;
   l550 = 0;
   l552 = 0;
   l554 = 0;
   l556 = 0;
   l558 = 0;
   l560 = 0;
   l562 = 0;
   l564 = 0;
   l566 = 0;
   l568 = 0;
   l570 = 0;
   l572 = 0;
   l574 = 0;
   l576 = 0;
   l578 = 0;
   l580 = 0;
   l582 = 0;
   l584 = 0;
   l586 = 0;
   l588 = 0;
   l590 = 0;
   l592 = 0;
   l594 = 0;
   l596 = 0;
   l598 = 0;
   l600 = 0;
   l602 = 0;
   l604 = 0;
   l606 = 0;
   l608 = 0;
   l610 = 0;
   l612 = 0;
   l614 = 0;
   l616 = 0;
   l618 = 0;
   l620 = 0;
   l622 = 0;
   l624 = 0;
   l626 = 0;
   l628 = 0;
   l630 = 0;
   l632 = 0;
   l634 = 0;
   l636 = 0;
   l638 = 0;
   l640 = 0;
   l642 = 0;
   l644 = 0;
   l646 = 0;
   l648 = 0;
   l650 = 0;
   l652 = 0;
   l654 = 0;
   l656 = 0;
   l658 = 0;
   l660 = 0;
   l662 = 0;
   l664 = 0;
   l666 = 0;
   l668 = 0;
   l670 = 0;
   l672 = 0;
   l674 = 0;
   l676 = 0;
   l678 = 0;
   l680 = 0;
   l682 = 0;
   l684 = 0;
   l686 = 0;
   l688 = 0;
   l690 = 0;
   l692 = 0;
   l694 = 0;
   l696 = 0;
   l698 = 0;
   l700 = 0;
   l702 = 0;
   l704 = 0;
   l706 = 0;
   l708 = 0;
   l710 = 0;
   l712 = 0;
   l714 = 0;
   l716 = 0;
   l718 = 0;
   l720 = 0;
   l722 = 0;
   l724 = 0;
   l726 = 0;
   l728 = 0;
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
   l802 = 0;
   l804 = 0;
   l806 = 0;
   l808 = 0;
   l810 = 0;
   l812 = 0;
   l814 = 0;
   l816 = 0;
   l818 = 0;
   l820 = 0;
   l822 = 0;
   l824 = 0;
   l826 = 0;
   l828 = 0;
   l830 = 0;
   l832 = 0;
   l834 = 0;
   l836 = 0;
   l838 = 0;
   l840 = 0;
   l842 = 0;
   l844 = 0;
   l846 = 0;
   l848 = 0;
   l850 = 0;
   l852 = 0;
   l854 = 0;
   l856 = 0;
   l858 = 0;
   l860 = 0;
   l862 = 0;
   l864 = 0;
   l866 = 0;
   l868 = 0;
   l870 = 0;
   l872 = 0;
   l874 = 0;
   l876 = 0;
   l878 = 0;
   l880 = 0;
   l882 = 0;
   l884 = 0;
   l886 = 0;
   l888 = 0;
   l890 = 0;
   l892 = 0;
   l894 = 0;
   l896 = 0;
   l898 = 0;
   l900 = 0;
   l902 = 0;
   l904 = 0;
   l906 = 0;
   l908 = 0;
   l910 = 0;
   l912 = 0;
   l914 = 0;
   l916 = 0;
   l918 = 0;
   l920 = 0;
   l922 = 0;
   l924 = 0;
   l926 = 0;
   l928 = 0;
   l930 = 0;
   l932 = 0;
   l934 = 0;
   l936 = 0;
   l938 = 0;
   l940 = 0;
   l942 = 0;
   l944 = 0;
   l946 = 0;
   l948 = 0;
   l950 = 0;
   l952 = 0;
   l954 = 0;
   l956 = 0;
   l958 = 0;
   l960 = 0;
   l962 = 0;
   l964 = 0;
   l966 = 0;
   l968 = 0;
   l970 = 0;
   l972 = 0;
   l974 = 0;
   l976 = 0;
   l978 = 0;
   l980 = 0;
   l982 = 0;
   l984 = 0;
   l986 = 0;
   l988 = 0;
   l990 = 0;
   l992 = 0;
   l994 = 0;
   l996 = 0;
   l998 = 0;
   l1000 = 0;
   l1002 = 0;
   l1004 = 0;
   l1006 = 0;
   l1008 = 0;
   l1010 = 0;
   l1012 = 0;
   l1014 = 0;
   l1016 = 0;
   l1018 = 0;
   l1020 = 0;
   l1022 = 0;
   l1024 = 0;
   l1026 = 0;
   l1028 = 0;
   l1030 = 0;
   l1032 = 0;
   l1034 = 0;
   l1036 = 0;
   l1038 = 0;
   l1040 = 0;
   l1042 = 0;
   l1044 = 0;
   l1046 = 0;
   l1048 = 0;
   l1050 = 0;
   l1052 = 0;
   l1054 = 0;
   l1056 = 0;
   l1058 = 0;
   l1060 = 0;
   l1062 = 0;
   l1064 = 0;
   l1066 = 0;
   l1068 = 0;
   l1070 = 0;
   l1072 = 0;
   l1074 = 0;
   l1076 = 0;
   l1078 = 0;
   l1080 = 0;
   l1082 = 0;
   l1084 = 0;
   l1086 = 0;
   l1088 = 0;
   l1090 = 0;
   l1092 = 0;
   l1094 = 0;
   l1096 = 0;
   l1098 = 0;
   l1100 = 0;
   l1102 = 0;
   l1104 = 0;
   l1106 = 0;
   l1108 = 0;
   l1110 = 0;
   l1112 = 0;
   l1114 = 0;
   l1116 = 0;
   l1118 = 0;
   l1120 = 0;
   l1122 = 0;
   l1124 = 0;
   l1126 = 0;
   l1128 = 0;
   l1130 = 0;
   l1132 = 0;
   l1134 = 0;
   l1136 = 0;
   l1138 = 0;
   l1140 = 0;
   l1142 = 0;
   l1144 = 0;
   l1146 = 0;
   l1148 = 0;
   l1150 = 0;
   l1152 = 0;
   l1154 = 0;
   l1156 = 0;
   l1158 = 0;
   l1160 = 0;
   l1162 = 0;
   l1164 = 0;
   l1166 = 0;
end

always @(posedge a1274)
   l60 <= a1274;

always @(posedge na1300)
   l62 <= na1300;

always @(posedge c1)
   l64 <= c1;

always @(posedge a1302)
   l66 <= a1302;

always @(posedge na1406)
   l68 <= na1406;

always @(posedge na1486)
   l70 <= na1486;

always @(posedge na1506)
   l72 <= na1506;

always @(posedge na1530)
   l74 <= na1530;

always @(posedge na1550)
   l76 <= na1550;

always @(posedge na1570)
   l78 <= na1570;

always @(posedge na1670)
   l80 <= na1670;

always @(posedge na1728)
   l82 <= na1728;

always @(posedge na1740)
   l84 <= na1740;

always @(posedge na1764)
   l86 <= na1764;

always @(posedge na1770)
   l88 <= na1770;

always @(posedge na1800)
   l90 <= na1800;

always @(posedge na1810)
   l92 <= na1810;

always @(posedge na1820)
   l94 <= na1820;

always @(posedge na1830)
   l96 <= na1830;

always @(posedge na1840)
   l98 <= na1840;

always @(posedge na1850)
   l100 <= na1850;

always @(posedge na1860)
   l102 <= na1860;

always @(posedge na1870)
   l104 <= na1870;

always @(posedge na1880)
   l106 <= na1880;

always @(posedge na1890)
   l108 <= na1890;

always @(posedge na1900)
   l110 <= na1900;

always @(posedge na1924)
   l112 <= na1924;

always @(posedge na1928)
   l114 <= na1928;

always @(posedge na1946)
   l116 <= na1946;

always @(posedge na1956)
   l118 <= na1956;

always @(posedge na1966)
   l120 <= na1966;

always @(posedge na2014)
   l122 <= na2014;

always @(posedge a2018)
   l124 <= a2018;

always @(posedge na2024)
   l126 <= na2024;

always @(posedge a2042)
   l128 <= a2042;

always @(posedge na2060)
   l130 <= na2060;

always @(posedge na2066)
   l132 <= na2066;

always @(posedge na2078)
   l134 <= na2078;

always @(posedge na2090)
   l136 <= na2090;

always @(posedge na2102)
   l138 <= na2102;

always @(posedge a2112)
   l140 <= a2112;

always @(posedge na2118)
   l142 <= na2118;

always @(posedge na2136)
   l144 <= na2136;

always @(posedge na2154)
   l146 <= na2154;

always @(posedge na2168)
   l148 <= na2168;

always @(posedge na2186)
   l150 <= na2186;

always @(posedge na2206)
   l152 <= na2206;

always @(posedge a2224)
   l154 <= a2224;

always @(posedge na2234)
   l156 <= na2234;

always @(posedge na2240)
   l158 <= na2240;

always @(posedge na2252)
   l160 <= na2252;

always @(posedge na2264)
   l162 <= na2264;

always @(posedge na2278)
   l164 <= na2278;

always @(posedge na2296)
   l166 <= na2296;

always @(posedge na2308)
   l168 <= na2308;

always @(posedge na2326)
   l170 <= na2326;

always @(posedge na2338)
   l172 <= na2338;

always @(posedge na2356)
   l174 <= na2356;

always @(posedge na2374)
   l176 <= na2374;

always @(posedge na2380)
   l178 <= na2380;

always @(posedge na2418)
   l180 <= na2418;

always @(posedge na2424)
   l182 <= na2424;

always @(posedge na2438)
   l184 <= na2438;

always @(posedge na2454)
   l186 <= na2454;

always @(posedge na2470)
   l188 <= na2470;

always @(posedge a2490)
   l190 <= a2490;

always @(posedge na2498)
   l192 <= na2498;

always @(posedge na2464)
   l194 <= na2464;

always @(posedge nl1064)
   l196 <= nl1064;

always @(posedge na2510)
   l198 <= na2510;

always @(posedge na2614)
   l200 <= na2614;

always @(posedge a2634)
   l202 <= a2634;

always @(posedge na2698)
   l204 <= na2698;

always @(posedge a2484)
   l206 <= a2484;

always @(posedge na2722)
   l208 <= na2722;

always @(posedge na2734)
   l210 <= na2734;

always @(posedge na2746)
   l212 <= na2746;

always @(posedge na2758)
   l214 <= na2758;

always @(posedge na2770)
   l216 <= na2770;

always @(posedge na2782)
   l218 <= na2782;

always @(posedge na2794)
   l220 <= na2794;

always @(posedge na2806)
   l222 <= na2806;

always @(posedge na2818)
   l224 <= na2818;

always @(posedge na2830)
   l226 <= na2830;

always @(posedge na2842)
   l228 <= na2842;

always @(posedge na2854)
   l230 <= na2854;

always @(posedge na2866)
   l232 <= na2866;

always @(posedge na2878)
   l234 <= na2878;

always @(posedge na2890)
   l236 <= na2890;

always @(posedge na2902)
   l238 <= na2902;

always @(posedge na2914)
   l240 <= na2914;

always @(posedge na2934)
   l242 <= na2934;

always @(posedge na2946)
   l244 <= na2946;

always @(posedge na2958)
   l246 <= na2958;

always @(posedge na2970)
   l248 <= na2970;

always @(posedge na2982)
   l250 <= na2982;

always @(posedge na2992)
   l252 <= na2992;

always @(posedge na3014)
   l254 <= na3014;

always @(posedge na3044)
   l256 <= na3044;

always @(posedge na3056)
   l258 <= na3056;

always @(posedge na2692)
   l260 <= na2692;

always @(posedge na3050)
   l262 <= na3050;

always @(posedge na3076)
   l264 <= na3076;

always @(posedge na3098)
   l266 <= na3098;

always @(posedge na3110)
   l268 <= na3110;

always @(posedge na3130)
   l270 <= na3130;

always @(posedge na3038)
   l272 <= na3038;

always @(posedge na3142)
   l274 <= na3142;

always @(posedge na3124)
   l276 <= na3124;

always @(posedge na3136)
   l278 <= na3136;

always @(posedge na3154)
   l280 <= na3154;

always @(posedge na3104)
   l282 <= na3104;

always @(posedge na3148)
   l284 <= na3148;

always @(posedge na3188)
   l286 <= na3188;

always @(posedge na3208)
   l288 <= na3208;

always @(posedge na3232)
   l290 <= na3232;

always @(posedge na3258)
   l292 <= na3258;

always @(posedge na3276)
   l294 <= na3276;

always @(posedge na3296)
   l296 <= na3296;

always @(posedge na3322)
   l298 <= na3322;

always @(posedge na3344)
   l300 <= na3344;

always @(posedge na3364)
   l302 <= na3364;

always @(posedge na3384)
   l304 <= na3384;

always @(posedge na3406)
   l306 <= na3406;

always @(posedge na3424)
   l308 <= na3424;

always @(posedge na3442)
   l310 <= na3442;

always @(posedge na3460)
   l312 <= na3460;

always @(posedge na3480)
   l314 <= na3480;

always @(posedge na3502)
   l316 <= na3502;

always @(posedge na3522)
   l318 <= na3522;

always @(posedge na3542)
   l320 <= na3542;

always @(posedge na3560)
   l322 <= na3560;

always @(posedge na3578)
   l324 <= na3578;

always @(posedge na3596)
   l326 <= na3596;

always @(posedge na3616)
   l328 <= na3616;

always @(posedge na3634)
   l330 <= na3634;

always @(posedge na3652)
   l332 <= na3652;

always @(posedge na3670)
   l334 <= na3670;

always @(posedge na3688)
   l336 <= na3688;

always @(posedge na3720)
   l338 <= na3720;

always @(posedge na3742)
   l340 <= na3742;

always @(posedge na3766)
   l342 <= na3766;

always @(posedge na3092)
   l344 <= na3092;

always @(posedge na3794)
   l346 <= na3794;

always @(posedge na3814)
   l348 <= na3814;

always @(posedge na3844)
   l350 <= na3844;

always @(posedge na3878)
   l352 <= na3878;

always @(posedge na3760)
   l354 <= na3760;

always @(posedge na3890)
   l356 <= na3890;

always @(posedge na3910)
   l358 <= na3910;

always @(posedge na3872)
   l360 <= na3872;

always @(posedge na3924)
   l362 <= na3924;

always @(posedge na3904)
   l364 <= na3904;

always @(posedge na3918)
   l366 <= na3918;

always @(posedge na3884)
   l368 <= na3884;

always @(posedge a3936)
   l370 <= a3936;

always @(posedge a3954)
   l372 <= a3954;

always @(posedge a3966)
   l374 <= a3966;

always @(posedge na3984)
   l376 <= na3984;

always @(posedge a3996)
   l378 <= a3996;

always @(posedge a4008)
   l380 <= a4008;

always @(posedge a4020)
   l382 <= a4020;

always @(posedge a4032)
   l384 <= a4032;

always @(posedge na3838)
   l386 <= na3838;

always @(posedge na4026)
   l388 <= na4026;

always @(posedge na4014)
   l390 <= na4014;

always @(posedge na4002)
   l392 <= na4002;

always @(posedge na3990)
   l394 <= na3990;

always @(posedge na3978)
   l396 <= na3978;

always @(posedge na3960)
   l398 <= na3960;

always @(posedge a3948)
   l400 <= a3948;

always @(posedge na3930)
   l402 <= na3930;

always @(posedge na3808)
   l404 <= na3808;

always @(posedge na4050)
   l406 <= na4050;

always @(posedge na4068)
   l408 <= na4068;

always @(posedge na4080)
   l410 <= na4080;

always @(posedge na4094)
   l412 <= na4094;

always @(posedge na4106)
   l414 <= na4106;

always @(posedge na3788)
   l416 <= na3788;

always @(posedge na4100)
   l418 <= na4100;

always @(posedge na4088)
   l420 <= na4088;

always @(posedge a4074)
   l422 <= a4074;

always @(posedge na4140)
   l424 <= na4140;

always @(posedge na4158)
   l426 <= na4158;

always @(posedge na4190)
   l428 <= na4190;

always @(posedge na4208)
   l430 <= na4208;

always @(posedge na4238)
   l432 <= na4238;

always @(posedge na4134)
   l434 <= na4134;

always @(posedge na4256)
   l436 <= na4256;

always @(posedge na4286)
   l438 <= na4286;

always @(posedge na4232)
   l440 <= na4232;

always @(posedge na4304)
   l442 <= na4304;

always @(posedge na4334)
   l444 <= na4334;

always @(posedge na4280)
   l446 <= na4280;

always @(posedge na4352)
   l448 <= na4352;

always @(posedge na4366)
   l450 <= na4366;

always @(posedge na4396)
   l452 <= na4396;

always @(posedge na4328)
   l454 <= na4328;

always @(posedge na4414)
   l456 <= na4414;

always @(posedge na4444)
   l458 <= na4444;

always @(posedge na4390)
   l460 <= na4390;

always @(posedge na4474)
   l462 <= na4474;

always @(posedge na4438)
   l464 <= na4438;

always @(posedge na4504)
   l466 <= na4504;

always @(posedge na4468)
   l468 <= na4468;

always @(posedge na4510)
   l470 <= na4510;

always @(posedge na4540)
   l472 <= na4540;

always @(posedge na4498)
   l474 <= na4498;

always @(posedge na4546)
   l476 <= na4546;

always @(posedge na4576)
   l478 <= na4576;

always @(posedge na4534)
   l480 <= na4534;

always @(posedge na4606)
   l482 <= na4606;

always @(posedge na4570)
   l484 <= na4570;

always @(posedge na4624)
   l486 <= na4624;

always @(posedge na4654)
   l488 <= na4654;

always @(posedge na4600)
   l490 <= na4600;

always @(posedge na4672)
   l492 <= na4672;

always @(posedge na4702)
   l494 <= na4702;

always @(posedge na4648)
   l496 <= na4648;

always @(posedge na4720)
   l498 <= na4720;

always @(posedge na4750)
   l500 <= na4750;

always @(posedge na4696)
   l502 <= na4696;

always @(posedge na4768)
   l504 <= na4768;

always @(posedge na4798)
   l506 <= na4798;

always @(posedge na4744)
   l508 <= na4744;

always @(posedge na4816)
   l510 <= na4816;

always @(posedge na4836)
   l512 <= na4836;

always @(posedge na4866)
   l514 <= na4866;

always @(posedge na4792)
   l516 <= na4792;

always @(posedge na4884)
   l518 <= na4884;

always @(posedge a4902)
   l520 <= a4902;

always @(posedge na4932)
   l522 <= na4932;

always @(posedge na4860)
   l524 <= na4860;

always @(posedge a4950)
   l526 <= a4950;

always @(posedge na4976)
   l528 <= na4976;

always @(posedge na4926)
   l530 <= na4926;

always @(posedge na4994)
   l532 <= na4994;

always @(posedge na5018)
   l534 <= na5018;

always @(posedge na4970)
   l536 <= na4970;

always @(posedge na5036)
   l538 <= na5036;

always @(posedge na5060)
   l540 <= na5060;

always @(posedge na5012)
   l542 <= na5012;

always @(posedge na5078)
   l544 <= na5078;

always @(posedge na5102)
   l546 <= na5102;

always @(posedge na5054)
   l548 <= na5054;

always @(posedge na5126)
   l550 <= na5126;

always @(posedge na5096)
   l552 <= na5096;

always @(posedge na5150)
   l554 <= na5150;

always @(posedge na5120)
   l556 <= na5120;

always @(posedge na5168)
   l558 <= na5168;

always @(posedge na5192)
   l560 <= na5192;

always @(posedge na5144)
   l562 <= na5144;

always @(posedge na5210)
   l564 <= na5210;

always @(posedge na5186)
   l566 <= na5186;

always @(posedge na5228)
   l568 <= na5228;

always @(posedge na5204)
   l570 <= na5204;

always @(posedge na5246)
   l572 <= na5246;

always @(posedge na5222)
   l574 <= na5222;

always @(posedge na5264)
   l576 <= na5264;

always @(posedge na5240)
   l578 <= na5240;

always @(posedge na5282)
   l580 <= na5282;

always @(posedge na5258)
   l582 <= na5258;

always @(posedge na5300)
   l584 <= na5300;

always @(posedge na5276)
   l586 <= na5276;

always @(posedge na5318)
   l588 <= na5318;

always @(posedge na5294)
   l590 <= na5294;

always @(posedge na5336)
   l592 <= na5336;

always @(posedge na5312)
   l594 <= na5312;

always @(posedge na5362)
   l596 <= na5362;

always @(posedge na5330)
   l598 <= na5330;

always @(posedge na5366)
   l600 <= na5366;

always @(posedge na5390)
   l602 <= na5390;

always @(posedge na5356)
   l604 <= na5356;

always @(posedge na5394)
   l606 <= na5394;

always @(posedge na5418)
   l608 <= na5418;

always @(posedge na5384)
   l610 <= na5384;

always @(posedge na5422)
   l612 <= na5422;

always @(posedge na5446)
   l614 <= na5446;

always @(posedge na5412)
   l616 <= na5412;

always @(posedge na5450)
   l618 <= na5450;

always @(posedge na5474)
   l620 <= na5474;

always @(posedge na5440)
   l622 <= na5440;

always @(posedge na5480)
   l624 <= na5480;

always @(posedge na5504)
   l626 <= na5504;

always @(posedge na5468)
   l628 <= na5468;

always @(posedge na5508)
   l630 <= na5508;

always @(posedge na5532)
   l632 <= na5532;

always @(posedge na5498)
   l634 <= na5498;

always @(posedge na5536)
   l636 <= na5536;

always @(posedge na5560)
   l638 <= na5560;

always @(posedge na5526)
   l640 <= na5526;

always @(posedge na5564)
   l642 <= na5564;

always @(posedge na5588)
   l644 <= na5588;

always @(posedge na5554)
   l646 <= na5554;

always @(posedge na5592)
   l648 <= na5592;

always @(posedge na5616)
   l650 <= na5616;

always @(posedge na5582)
   l652 <= na5582;

always @(posedge na5620)
   l654 <= na5620;

always @(posedge na5644)
   l656 <= na5644;

always @(posedge na5610)
   l658 <= na5610;

always @(posedge na5648)
   l660 <= na5648;

always @(posedge na5672)
   l662 <= na5672;

always @(posedge na5638)
   l664 <= na5638;

always @(posedge na5676)
   l666 <= na5676;

always @(posedge na5700)
   l668 <= na5700;

always @(posedge na5666)
   l670 <= na5666;

always @(posedge na5704)
   l672 <= na5704;

always @(posedge na5728)
   l674 <= na5728;

always @(posedge na5694)
   l676 <= na5694;

always @(posedge na5732)
   l678 <= na5732;

always @(posedge na5750)
   l680 <= na5750;

always @(posedge na5722)
   l682 <= na5722;

always @(posedge na5768)
   l684 <= na5768;

always @(posedge na5744)
   l686 <= na5744;

always @(posedge na5786)
   l688 <= na5786;

always @(posedge na5762)
   l690 <= na5762;

always @(posedge na5804)
   l692 <= na5804;

always @(posedge na5780)
   l694 <= na5780;

always @(posedge na5822)
   l696 <= na5822;

always @(posedge na5798)
   l698 <= na5798;

always @(posedge na5840)
   l700 <= na5840;

always @(posedge na5816)
   l702 <= na5816;

always @(posedge na5858)
   l704 <= na5858;

always @(posedge na5834)
   l706 <= na5834;

always @(posedge na5876)
   l708 <= na5876;

always @(posedge na5852)
   l710 <= na5852;

always @(posedge na5894)
   l712 <= na5894;

always @(posedge na5870)
   l714 <= na5870;

always @(posedge na5912)
   l716 <= na5912;

always @(posedge na5888)
   l718 <= na5888;

always @(posedge na5930)
   l720 <= na5930;

always @(posedge na5906)
   l722 <= na5906;

always @(posedge na5948)
   l724 <= na5948;

always @(posedge na5924)
   l726 <= na5924;

always @(posedge na5966)
   l728 <= na5966;

always @(posedge na5942)
   l730 <= na5942;

always @(posedge na5984)
   l732 <= na5984;

always @(posedge na5960)
   l734 <= na5960;

always @(posedge na6002)
   l736 <= na6002;

always @(posedge na5978)
   l738 <= na5978;

always @(posedge na6020)
   l740 <= na6020;

always @(posedge na5996)
   l742 <= na5996;

always @(posedge na6038)
   l744 <= na6038;

always @(posedge na6014)
   l746 <= na6014;

always @(posedge na6058)
   l748 <= na6058;

always @(posedge na6032)
   l750 <= na6032;

always @(posedge na6074)
   l752 <= na6074;

always @(posedge na6052)
   l754 <= na6052;

always @(posedge na6068)
   l756 <= na6068;

always @(posedge na6170)
   l758 <= na6170;

always @(posedge na6194)
   l760 <= na6194;

always @(posedge na6214)
   l762 <= na6214;

always @(posedge na6236)
   l764 <= na6236;

always @(posedge na6256)
   l766 <= na6256;

always @(posedge na6276)
   l768 <= na6276;

always @(posedge na6296)
   l770 <= na6296;

always @(posedge na6316)
   l772 <= na6316;

always @(posedge na6350)
   l774 <= na6350;

always @(posedge na6370)
   l776 <= na6370;

always @(posedge na6390)
   l778 <= na6390;

always @(posedge na6410)
   l780 <= na6410;

always @(posedge na6430)
   l782 <= na6430;

always @(posedge na6450)
   l784 <= na6450;

always @(posedge na6470)
   l786 <= na6470;

always @(posedge na6490)
   l788 <= na6490;

always @(posedge na6516)
   l790 <= na6516;

always @(posedge na6524)
   l792 <= na6524;

always @(posedge na6310)
   l794 <= na6310;

always @(posedge na6528)
   l796 <= na6528;

always @(posedge na6540)
   l798 <= na6540;

always @(posedge na6534)
   l800 <= na6534;

always @(posedge na6554)
   l802 <= na6554;

always @(posedge na6566)
   l804 <= na6566;

always @(posedge na6578)
   l806 <= na6578;

always @(posedge na6510)
   l808 <= na6510;

always @(posedge nl814)
   l810 <= nl814;

always @(posedge na6572)
   l812 <= na6572;

always @(posedge z0)
   l814 <= z0;

always @(posedge na6560)
   l816 <= na6560;

always @(posedge na6548)
   l818 <= na6548;

always @(posedge na6484)
   l820 <= na6484;

always @(posedge na6464)
   l822 <= na6464;

always @(posedge na6444)
   l824 <= na6444;

always @(posedge na6424)
   l826 <= na6424;

always @(posedge na6404)
   l828 <= na6404;

always @(posedge na6384)
   l830 <= na6384;

always @(posedge na6364)
   l832 <= na6364;

always @(posedge na6344)
   l834 <= na6344;

always @(posedge na6290)
   l836 <= na6290;

always @(posedge na6270)
   l838 <= na6270;

always @(posedge na6250)
   l840 <= na6250;

always @(posedge na6230)
   l842 <= na6230;

always @(posedge na6208)
   l844 <= na6208;

always @(posedge na6188)
   l846 <= na6188;

always @(posedge na6606)
   l848 <= na6606;

always @(posedge na6626)
   l850 <= na6626;

always @(posedge na6632)
   l852 <= na6632;

always @(posedge na6600)
   l854 <= na6600;

always @(posedge na6646)
   l856 <= na6646;

always @(posedge na6666)
   l858 <= na6666;

always @(posedge na6620)
   l860 <= na6620;

always @(posedge na6660)
   l862 <= na6660;

always @(posedge na6640)
   l864 <= na6640;

always @(posedge na6678)
   l866 <= na6678;

always @(posedge na6672)
   l868 <= na6672;

always @(posedge na6684)
   l870 <= na6684;

always @(posedge na6702)
   l872 <= na6702;

always @(posedge na5162)
   l874 <= na5162;

always @(posedge a6708)
   l876 <= a6708;

always @(posedge na6696)
   l878 <= na6696;

always @(posedge na6704)
   l880 <= na6704;

always @(posedge na5072)
   l882 <= na5072;

always @(posedge na5030)
   l884 <= na5030;

always @(posedge na4988)
   l886 <= na4988;

always @(posedge a4944)
   l888 <= a4944;

always @(posedge a4896)
   l890 <= a4896;

always @(posedge na4878)
   l892 <= na4878;

always @(posedge na4830)
   l894 <= na4830;

always @(posedge na4810)
   l896 <= na4810;

always @(posedge na4762)
   l898 <= na4762;

always @(posedge na4714)
   l900 <= na4714;

always @(posedge na4666)
   l902 <= na4666;

always @(posedge na4618)
   l904 <= na4618;

always @(posedge na4408)
   l906 <= na4408;

always @(posedge na4346)
   l908 <= na4346;

always @(posedge na4298)
   l910 <= na4298;

always @(posedge na4250)
   l912 <= na4250;

always @(posedge na4202)
   l914 <= na4202;

always @(posedge na6724)
   l916 <= na6724;

always @(posedge na6870)
   l918 <= na6870;

always @(posedge na4184)
   l920 <= na4184;

always @(posedge na6864)
   l922 <= na6864;

always @(posedge na6718)
   l924 <= na6718;

always @(posedge na4152)
   l926 <= na4152;

always @(posedge na6888)
   l928 <= na6888;

always @(posedge na6908)
   l930 <= na6908;

always @(posedge na6926)
   l932 <= na6926;

always @(posedge na6944)
   l934 <= na6944;

always @(posedge na6970)
   l936 <= na6970;

always @(posedge na4062)
   l938 <= na4062;

always @(posedge na6964)
   l940 <= na6964;

always @(posedge na6938)
   l942 <= na6938;

always @(posedge na6920)
   l944 <= na6920;

always @(posedge na6902)
   l946 <= na6902;

always @(posedge na6882)
   l948 <= na6882;

always @(posedge na4044)
   l950 <= na4044;

always @(posedge na3736)
   l952 <= na3736;

always @(posedge na3714)
   l954 <= na3714;

always @(posedge na3682)
   l956 <= na3682;

always @(posedge na3664)
   l958 <= na3664;

always @(posedge na3646)
   l960 <= na3646;

always @(posedge na3628)
   l962 <= na3628;

always @(posedge na3610)
   l964 <= na3610;

always @(posedge na3590)
   l966 <= na3590;

always @(posedge na3572)
   l968 <= na3572;

always @(posedge na3554)
   l970 <= na3554;

always @(posedge na3536)
   l972 <= na3536;

always @(posedge na3516)
   l974 <= na3516;

always @(posedge na3496)
   l976 <= na3496;

always @(posedge na3474)
   l978 <= na3474;

always @(posedge na3454)
   l980 <= na3454;

always @(posedge na3436)
   l982 <= na3436;

always @(posedge na3418)
   l984 <= na3418;

always @(posedge na3400)
   l986 <= na3400;

always @(posedge na3378)
   l988 <= na3378;

always @(posedge na3358)
   l990 <= na3358;

always @(posedge na3338)
   l992 <= na3338;

always @(posedge na3316)
   l994 <= na3316;

always @(posedge na3290)
   l996 <= na3290;

always @(posedge na3270)
   l998 <= na3270;

always @(posedge na3252)
   l1000 <= na3252;

always @(posedge na3226)
   l1002 <= na3226;

always @(posedge na3202)
   l1004 <= na3202;

always @(posedge na3182)
   l1006 <= na3182;

always @(posedge na3070)
   l1008 <= na3070;

always @(posedge na3008)
   l1010 <= na3008;

always @(posedge a2986)
   l1012 <= a2986;

always @(posedge na2976)
   l1014 <= na2976;

always @(posedge na2964)
   l1016 <= na2964;

always @(posedge na2952)
   l1018 <= na2952;

always @(posedge na2940)
   l1020 <= na2940;

always @(posedge na2928)
   l1022 <= na2928;

always @(posedge na2908)
   l1024 <= na2908;

always @(posedge na2896)
   l1026 <= na2896;

always @(posedge na2884)
   l1028 <= na2884;

always @(posedge na2872)
   l1030 <= na2872;

always @(posedge na2860)
   l1032 <= na2860;

always @(posedge na2848)
   l1034 <= na2848;

always @(posedge na2836)
   l1036 <= na2836;

always @(posedge na2824)
   l1038 <= na2824;

always @(posedge na2812)
   l1040 <= na2812;

always @(posedge na2800)
   l1042 <= na2800;

always @(posedge na2788)
   l1044 <= na2788;

always @(posedge na2776)
   l1046 <= na2776;

always @(posedge na2764)
   l1048 <= na2764;

always @(posedge na2752)
   l1050 <= na2752;

always @(posedge na2740)
   l1052 <= na2740;

always @(posedge na2728)
   l1054 <= na2728;

always @(posedge na2716)
   l1056 <= na2716;

always @(posedge a2628)
   l1058 <= a2628;

always @(posedge na2608)
   l1060 <= na2608;

always @(posedge na2504)
   l1062 <= na2504;

always @(posedge l1066)
   l1064 <= l1066;

always @(posedge l1068)
   l1066 <= l1068;

always @(posedge z1)
   l1068 <= z1;

always @(posedge na2448)
   l1070 <= na2448;

always @(posedge na2432)
   l1072 <= na2432;

always @(posedge na6990)
   l1074 <= na6990;

always @(posedge na7008)
   l1076 <= na7008;

always @(posedge na7026)
   l1078 <= na7026;

always @(posedge na2412)
   l1080 <= na2412;

always @(posedge na7020)
   l1082 <= na7020;

always @(posedge na7002)
   l1084 <= na7002;

always @(posedge na6984)
   l1086 <= na6984;

always @(posedge na2368)
   l1088 <= na2368;

always @(posedge na2350)
   l1090 <= na2350;

always @(posedge na2332)
   l1092 <= na2332;

always @(posedge na2320)
   l1094 <= na2320;

always @(posedge na7032)
   l1096 <= na7032;

always @(posedge na2290)
   l1098 <= na2290;

always @(posedge na2270)
   l1100 <= na2270;

always @(posedge na2258)
   l1102 <= na2258;

always @(posedge na2246)
   l1104 <= na2246;

always @(posedge a2218)
   l1106 <= a2218;

always @(posedge na7036)
   l1108 <= na7036;

always @(posedge na7052)
   l1110 <= na7052;

always @(posedge na7058)
   l1112 <= na7058;

always @(posedge na7046)
   l1114 <= na7046;

always @(posedge na7070)
   l1116 <= na7070;

always @(posedge na7074)
   l1118 <= na7074;

always @(posedge a7064)
   l1120 <= a7064;

always @(posedge na2180)
   l1122 <= na2180;

always @(posedge na2162)
   l1124 <= na2162;

always @(posedge na2148)
   l1126 <= na2148;

always @(posedge na2096)
   l1128 <= na2096;

always @(posedge na2084)
   l1130 <= na2084;

always @(posedge na2072)
   l1132 <= na2072;

always @(posedge na2054)
   l1134 <= na2054;

always @(posedge na2008)
   l1136 <= na2008;

always @(posedge na7086)
   l1138 <= na7086;

always @(posedge na7106)
   l1140 <= na7106;

always @(posedge na7118)
   l1142 <= na7118;

always @(posedge na7140)
   l1144 <= na7140;

always @(posedge na7134)
   l1146 <= na7134;

always @(posedge na7112)
   l1148 <= na7112;

always @(posedge na7100)
   l1150 <= na7100;

always @(posedge na7080)
   l1152 <= na7080;

always @(posedge na1940)
   l1154 <= na1940;

always @(posedge na1758)
   l1156 <= na1758;

always @(posedge na1564)
   l1158 <= na1564;

always @(posedge na1544)
   l1160 <= na1544;

always @(posedge na1524)
   l1162 <= na1524;

always @(posedge na1500)
   l1164 <= na1500;

always @(posedge na1480)
   l1166 <= na1480;


assign a1274 = ~a1272 & ~a1270;
assign na1300 = ~a1300;
assign c1 = 1;
assign a1302 = l66 & ~l64;
assign na1406 = ~a1406;
assign na1486 = ~a1486;
assign na1506 = ~a1506;
assign na1530 = ~a1530;
assign na1550 = ~a1550;
assign na1570 = ~a1570;
assign na1670 = ~a1670;
assign na1728 = ~a1728;
assign na1740 = ~a1740;
assign na1764 = ~a1764;
assign na1770 = ~a1770;
assign na1800 = ~a1800;
assign na1810 = ~a1810;
assign na1820 = ~a1820;
assign na1830 = ~a1830;
assign na1840 = ~a1840;
assign na1850 = ~a1850;
assign na1860 = ~a1860;
assign na1870 = ~a1870;
assign na1880 = ~a1880;
assign na1890 = ~a1890;
assign na1900 = ~a1900;
assign na1924 = ~a1924;
assign na1928 = ~a1928;
assign na1946 = ~a1946;
assign na1956 = ~a1956;
assign na1966 = ~a1966;
assign na2014 = ~a2014;
assign a2018 = ~a2016 & ~a1736;
assign na2024 = ~a2024;
assign a2042 = ~a2040 & ~a2030;
assign na2060 = ~a2060;
assign na2066 = ~a2066;
assign na2078 = ~a2078;
assign na2090 = ~a2090;
assign na2102 = ~a2102;
assign a2112 = ~a2110 & ~a2106;
assign na2118 = ~a2118;
assign na2136 = ~a2136;
assign na2154 = ~a2154;
assign na2168 = ~a2168;
assign na2186 = ~a2186;
assign na2206 = ~a2206;
assign a2224 = ~a2222 & ~a2220;
assign na2234 = ~a2234;
assign na2240 = ~a2240;
assign na2252 = ~a2252;
assign na2264 = ~a2264;
assign na2278 = ~a2278;
assign na2296 = ~a2296;
assign na2308 = ~a2308;
assign na2326 = ~a2326;
assign na2338 = ~a2338;
assign na2356 = ~a2356;
assign na2374 = ~a2374;
assign na2380 = ~a2380;
assign na2418 = ~a2418;
assign na2424 = ~a2424;
assign na2438 = ~a2438;
assign na2454 = ~a2454;
assign na2470 = ~a2470;
assign a2490 = ~a2488 & ~a2486;
assign na2498 = ~a2498;
assign na2464 = ~a2464;
assign nl1064 = ~l1064;
assign na2510 = ~a2510;
assign na2614 = ~a2614;
assign a2634 = ~a2632 & ~a2630;
assign na2698 = ~a2698;
assign a2484 = ~a2482 & ~a2480;
assign na2722 = ~a2722;
assign na2734 = ~a2734;
assign na2746 = ~a2746;
assign na2758 = ~a2758;
assign na2770 = ~a2770;
assign na2782 = ~a2782;
assign na2794 = ~a2794;
assign na2806 = ~a2806;
assign na2818 = ~a2818;
assign na2830 = ~a2830;
assign na2842 = ~a2842;
assign na2854 = ~a2854;
assign na2866 = ~a2866;
assign na2878 = ~a2878;
assign na2890 = ~a2890;
assign na2902 = ~a2902;
assign na2914 = ~a2914;
assign na2934 = ~a2934;
assign na2946 = ~a2946;
assign na2958 = ~a2958;
assign na2970 = ~a2970;
assign na2982 = ~a2982;
assign na2992 = ~a2992;
assign na3014 = ~a3014;
assign na3044 = ~a3044;
assign na3056 = ~a3056;
assign na2692 = ~a2692;
assign na3050 = ~a3050;
assign na3076 = ~a3076;
assign na3098 = ~a3098;
assign na3110 = ~a3110;
assign na3130 = ~a3130;
assign na3038 = ~a3038;
assign na3142 = ~a3142;
assign na3124 = ~a3124;
assign na3136 = ~a3136;
assign na3154 = ~a3154;
assign na3104 = ~a3104;
assign na3148 = ~a3148;
assign na3188 = ~a3188;
assign na3208 = ~a3208;
assign na3232 = ~a3232;
assign na3258 = ~a3258;
assign na3276 = ~a3276;
assign na3296 = ~a3296;
assign na3322 = ~a3322;
assign na3344 = ~a3344;
assign na3364 = ~a3364;
assign na3384 = ~a3384;
assign na3406 = ~a3406;
assign na3424 = ~a3424;
assign na3442 = ~a3442;
assign na3460 = ~a3460;
assign na3480 = ~a3480;
assign na3502 = ~a3502;
assign na3522 = ~a3522;
assign na3542 = ~a3542;
assign na3560 = ~a3560;
assign na3578 = ~a3578;
assign na3596 = ~a3596;
assign na3616 = ~a3616;
assign na3634 = ~a3634;
assign na3652 = ~a3652;
assign na3670 = ~a3670;
assign na3688 = ~a3688;
assign na3720 = ~a3720;
assign na3742 = ~a3742;
assign na3766 = ~a3766;
assign na3092 = ~a3092;
assign na3794 = ~a3794;
assign na3814 = ~a3814;
assign na3844 = ~a3844;
assign na3878 = ~a3878;
assign na3760 = ~a3760;
assign na3890 = ~a3890;
assign na3910 = ~a3910;
assign na3872 = ~a3872;
assign na3924 = ~a3924;
assign na3904 = ~a3904;
assign na3918 = ~a3918;
assign na3884 = ~a3884;
assign a3936 = ~a3934 & ~a3932;
assign a3954 = ~a3952 & ~a3950;
assign a3966 = ~a3964 & ~a3962;
assign na3984 = ~a3984;
assign a3996 = ~a3994 & ~a3992;
assign a4008 = ~a4006 & ~a4004;
assign a4020 = ~a4018 & ~a4016;
assign a4032 = ~a4030 & ~a4028;
assign na3838 = ~a3838;
assign na4026 = ~a4026;
assign na4014 = ~a4014;
assign na4002 = ~a4002;
assign na3990 = ~a3990;
assign na3978 = ~a3978;
assign na3960 = ~a3960;
assign a3948 = ~a3946 & ~a3944;
assign na3930 = ~a3930;
assign na3808 = ~a3808;
assign na4050 = ~a4050;
assign na4068 = ~a4068;
assign na4080 = ~a4080;
assign na4094 = ~a4094;
assign na4106 = ~a4106;
assign na3788 = ~a3788;
assign na4100 = ~a4100;
assign na4088 = ~a4088;
assign a4074 = ~a4072 & ~a4070;
assign na4140 = ~a4140;
assign na4158 = ~a4158;
assign na4190 = ~a4190;
assign na4208 = ~a4208;
assign na4238 = ~a4238;
assign na4134 = ~a4134;
assign na4256 = ~a4256;
assign na4286 = ~a4286;
assign na4232 = ~a4232;
assign na4304 = ~a4304;
assign na4334 = ~a4334;
assign na4280 = ~a4280;
assign na4352 = ~a4352;
assign na4366 = ~a4366;
assign na4396 = ~a4396;
assign na4328 = ~a4328;
assign na4414 = ~a4414;
assign na4444 = ~a4444;
assign na4390 = ~a4390;
assign na4474 = ~a4474;
assign na4438 = ~a4438;
assign na4504 = ~a4504;
assign na4468 = ~a4468;
assign na4510 = ~a4510;
assign na4540 = ~a4540;
assign na4498 = ~a4498;
assign na4546 = ~a4546;
assign na4576 = ~a4576;
assign na4534 = ~a4534;
assign na4606 = ~a4606;
assign na4570 = ~a4570;
assign na4624 = ~a4624;
assign na4654 = ~a4654;
assign na4600 = ~a4600;
assign na4672 = ~a4672;
assign na4702 = ~a4702;
assign na4648 = ~a4648;
assign na4720 = ~a4720;
assign na4750 = ~a4750;
assign na4696 = ~a4696;
assign na4768 = ~a4768;
assign na4798 = ~a4798;
assign na4744 = ~a4744;
assign na4816 = ~a4816;
assign na4836 = ~a4836;
assign na4866 = ~a4866;
assign na4792 = ~a4792;
assign na4884 = ~a4884;
assign a4902 = ~a4900 & ~a4898;
assign na4932 = ~a4932;
assign na4860 = ~a4860;
assign a4950 = ~a4948 & ~a4946;
assign na4976 = ~a4976;
assign na4926 = ~a4926;
assign na4994 = ~a4994;
assign na5018 = ~a5018;
assign na4970 = ~a4970;
assign na5036 = ~a5036;
assign na5060 = ~a5060;
assign na5012 = ~a5012;
assign na5078 = ~a5078;
assign na5102 = ~a5102;
assign na5054 = ~a5054;
assign na5126 = ~a5126;
assign na5096 = ~a5096;
assign na5150 = ~a5150;
assign na5120 = ~a5120;
assign na5168 = ~a5168;
assign na5192 = ~a5192;
assign na5144 = ~a5144;
assign na5210 = ~a5210;
assign na5186 = ~a5186;
assign na5228 = ~a5228;
assign na5204 = ~a5204;
assign na5246 = ~a5246;
assign na5222 = ~a5222;
assign na5264 = ~a5264;
assign na5240 = ~a5240;
assign na5282 = ~a5282;
assign na5258 = ~a5258;
assign na5300 = ~a5300;
assign na5276 = ~a5276;
assign na5318 = ~a5318;
assign na5294 = ~a5294;
assign na5336 = ~a5336;
assign na5312 = ~a5312;
assign na5362 = ~a5362;
assign na5330 = ~a5330;
assign na5366 = ~a5366;
assign na5390 = ~a5390;
assign na5356 = ~a5356;
assign na5394 = ~a5394;
assign na5418 = ~a5418;
assign na5384 = ~a5384;
assign na5422 = ~a5422;
assign na5446 = ~a5446;
assign na5412 = ~a5412;
assign na5450 = ~a5450;
assign na5474 = ~a5474;
assign na5440 = ~a5440;
assign na5480 = ~a5480;
assign na5504 = ~a5504;
assign na5468 = ~a5468;
assign na5508 = ~a5508;
assign na5532 = ~a5532;
assign na5498 = ~a5498;
assign na5536 = ~a5536;
assign na5560 = ~a5560;
assign na5526 = ~a5526;
assign na5564 = ~a5564;
assign na5588 = ~a5588;
assign na5554 = ~a5554;
assign na5592 = ~a5592;
assign na5616 = ~a5616;
assign na5582 = ~a5582;
assign na5620 = ~a5620;
assign na5644 = ~a5644;
assign na5610 = ~a5610;
assign na5648 = ~a5648;
assign na5672 = ~a5672;
assign na5638 = ~a5638;
assign na5676 = ~a5676;
assign na5700 = ~a5700;
assign na5666 = ~a5666;
assign na5704 = ~a5704;
assign na5728 = ~a5728;
assign na5694 = ~a5694;
assign na5732 = ~a5732;
assign na5750 = ~a5750;
assign na5722 = ~a5722;
assign na5768 = ~a5768;
assign na5744 = ~a5744;
assign na5786 = ~a5786;
assign na5762 = ~a5762;
assign na5804 = ~a5804;
assign na5780 = ~a5780;
assign na5822 = ~a5822;
assign na5798 = ~a5798;
assign na5840 = ~a5840;
assign na5816 = ~a5816;
assign na5858 = ~a5858;
assign na5834 = ~a5834;
assign na5876 = ~a5876;
assign na5852 = ~a5852;
assign na5894 = ~a5894;
assign na5870 = ~a5870;
assign na5912 = ~a5912;
assign na5888 = ~a5888;
assign na5930 = ~a5930;
assign na5906 = ~a5906;
assign na5948 = ~a5948;
assign na5924 = ~a5924;
assign na5966 = ~a5966;
assign na5942 = ~a5942;
assign na5984 = ~a5984;
assign na5960 = ~a5960;
assign na6002 = ~a6002;
assign na5978 = ~a5978;
assign na6020 = ~a6020;
assign na5996 = ~a5996;
assign na6038 = ~a6038;
assign na6014 = ~a6014;
assign na6058 = ~a6058;
assign na6032 = ~a6032;
assign na6074 = ~a6074;
assign na6052 = ~a6052;
assign na6068 = ~a6068;
assign na6170 = ~a6170;
assign na6194 = ~a6194;
assign na6214 = ~a6214;
assign na6236 = ~a6236;
assign na6256 = ~a6256;
assign na6276 = ~a6276;
assign na6296 = ~a6296;
assign na6316 = ~a6316;
assign na6350 = ~a6350;
assign na6370 = ~a6370;
assign na6390 = ~a6390;
assign na6410 = ~a6410;
assign na6430 = ~a6430;
assign na6450 = ~a6450;
assign na6470 = ~a6470;
assign na6490 = ~a6490;
assign na6516 = ~a6516;
assign na6524 = ~a6524;
assign na6310 = ~a6310;
assign na6528 = ~a6528;
assign na6540 = ~a6540;
assign na6534 = ~a6534;
assign na6554 = ~a6554;
assign na6566 = ~a6566;
assign na6578 = ~a6578;
assign na6510 = ~a6510;
assign nl814 = ~l814;
assign na6572 = ~a6572;
assign z0 = l810;
assign na6560 = ~a6560;
assign na6548 = ~a6548;
assign na6484 = ~a6484;
assign na6464 = ~a6464;
assign na6444 = ~a6444;
assign na6424 = ~a6424;
assign na6404 = ~a6404;
assign na6384 = ~a6384;
assign na6364 = ~a6364;
assign na6344 = ~a6344;
assign na6290 = ~a6290;
assign na6270 = ~a6270;
assign na6250 = ~a6250;
assign na6230 = ~a6230;
assign na6208 = ~a6208;
assign na6188 = ~a6188;
assign na6606 = ~a6606;
assign na6626 = ~a6626;
assign na6632 = ~a6632;
assign na6600 = ~a6600;
assign na6646 = ~a6646;
assign na6666 = ~a6666;
assign na6620 = ~a6620;
assign na6660 = ~a6660;
assign na6640 = ~a6640;
assign na6678 = ~a6678;
assign na6672 = ~a6672;
assign na6684 = ~a6684;
assign na6702 = ~a6702;
assign na5162 = ~a5162;
assign a6708 = ~a6706 & ~a6704;
assign na6696 = ~a6696;
assign na6704 = ~a6704;
assign na5072 = ~a5072;
assign na5030 = ~a5030;
assign na4988 = ~a4988;
assign a4944 = ~a4942 & ~a4940;
assign a4896 = ~a4894 & ~a4892;
assign na4878 = ~a4878;
assign na4830 = ~a4830;
assign na4810 = ~a4810;
assign na4762 = ~a4762;
assign na4714 = ~a4714;
assign na4666 = ~a4666;
assign na4618 = ~a4618;
assign na4408 = ~a4408;
assign na4346 = ~a4346;
assign na4298 = ~a4298;
assign na4250 = ~a4250;
assign na4202 = ~a4202;
assign na6724 = ~a6724;
assign na6870 = ~a6870;
assign na4184 = ~a4184;
assign na6864 = ~a6864;
assign na6718 = ~a6718;
assign na4152 = ~a4152;
assign na6888 = ~a6888;
assign na6908 = ~a6908;
assign na6926 = ~a6926;
assign na6944 = ~a6944;
assign na6970 = ~a6970;
assign na4062 = ~a4062;
assign na6964 = ~a6964;
assign na6938 = ~a6938;
assign na6920 = ~a6920;
assign na6902 = ~a6902;
assign na6882 = ~a6882;
assign na4044 = ~a4044;
assign na3736 = ~a3736;
assign na3714 = ~a3714;
assign na3682 = ~a3682;
assign na3664 = ~a3664;
assign na3646 = ~a3646;
assign na3628 = ~a3628;
assign na3610 = ~a3610;
assign na3590 = ~a3590;
assign na3572 = ~a3572;
assign na3554 = ~a3554;
assign na3536 = ~a3536;
assign na3516 = ~a3516;
assign na3496 = ~a3496;
assign na3474 = ~a3474;
assign na3454 = ~a3454;
assign na3436 = ~a3436;
assign na3418 = ~a3418;
assign na3400 = ~a3400;
assign na3378 = ~a3378;
assign na3358 = ~a3358;
assign na3338 = ~a3338;
assign na3316 = ~a3316;
assign na3290 = ~a3290;
assign na3270 = ~a3270;
assign na3252 = ~a3252;
assign na3226 = ~a3226;
assign na3202 = ~a3202;
assign na3182 = ~a3182;
assign na3070 = ~a3070;
assign na3008 = ~a3008;
assign a2986 = ~a2984 & ~a2646;
assign na2976 = ~a2976;
assign na2964 = ~a2964;
assign na2952 = ~a2952;
assign na2940 = ~a2940;
assign na2928 = ~a2928;
assign na2908 = ~a2908;
assign na2896 = ~a2896;
assign na2884 = ~a2884;
assign na2872 = ~a2872;
assign na2860 = ~a2860;
assign na2848 = ~a2848;
assign na2836 = ~a2836;
assign na2824 = ~a2824;
assign na2812 = ~a2812;
assign na2800 = ~a2800;
assign na2788 = ~a2788;
assign na2776 = ~a2776;
assign na2764 = ~a2764;
assign na2752 = ~a2752;
assign na2740 = ~a2740;
assign na2728 = ~a2728;
assign na2716 = ~a2716;
assign a2628 = ~a2626 & ~a2624;
assign na2608 = ~a2608;
assign na2504 = ~a2504;
assign z1 = l196;
assign na2448 = ~a2448;
assign na2432 = ~a2432;
assign na6990 = ~a6990;
assign na7008 = ~a7008;
assign na7026 = ~a7026;
assign na2412 = ~a2412;
assign na7020 = ~a7020;
assign na7002 = ~a7002;
assign na6984 = ~a6984;
assign na2368 = ~a2368;
assign na2350 = ~a2350;
assign na2332 = ~a2332;
assign na2320 = ~a2320;
assign na7032 = ~a7032;
assign na2290 = ~a2290;
assign na2270 = ~a2270;
assign na2258 = ~a2258;
assign na2246 = ~a2246;
assign a2218 = ~a2216 & ~a2214;
assign na7036 = ~a7036;
assign na7052 = ~a7052;
assign na7058 = ~a7058;
assign na7046 = ~a7046;
assign na7070 = ~a7070;
assign na7074 = ~a7074;
assign a7064 = ~a7062 & ~a7060;
assign na2180 = ~a2180;
assign na2162 = ~a2162;
assign na2148 = ~a2148;
assign na2096 = ~a2096;
assign na2084 = ~a2084;
assign na2072 = ~a2072;
assign na2054 = ~a2054;
assign na2008 = ~a2008;
assign na7086 = ~a7086;
assign na7106 = ~a7106;
assign na7118 = ~a7118;
assign na7140 = ~a7140;
assign na7134 = ~a7134;
assign na7112 = ~a7112;
assign na7100 = ~a7100;
assign na7080 = ~a7080;
assign na1940 = ~a1940;
assign na1758 = ~a1758;
assign na1564 = ~a1564;
assign na1544 = ~a1544;
assign na1524 = ~a1524;
assign na1500 = ~a1500;
assign na1480 = ~a1480;
assign a1168 = ~l68 & ~l66;
assign a1170 = ~a1168 & ~l60;
assign a1172 = ~l162 & l160;
assign a1174 = a1172 & l158;
assign a1176 = a1174 & l84;
assign a1178 = l168 & l166;
assign a1180 = l170 & ~l168;
assign a1182 = ~a1180 & ~a1178;
assign a1184 = ~a1182 & ~l172;
assign a1186 = ~a1184 & ~l126;
assign a1188 = ~a1186 & l164;
assign a1190 = ~a1188 & ~a1176;
assign a1192 = l164 & l84;
assign a1194 = a1192 & a1190;
assign a1196 = ~l82 & ~l80;
assign a1198 = a1196 & ~l60;
assign a1200 = ~a1198 & ~a1194;
assign a1202 = ~l148 & ~l146;
assign a1204 = l152 & ~l150;
assign a1206 = a1204 & a1202;
assign a1208 = l184 & l182;
assign a1210 = l186 & ~l84;
assign a1212 = a1210 & a1208;
assign a1214 = a1212 & ~a1206;
assign a1216 = ~l188 & ~l174;
assign a1218 = a1216 & ~a1214;
assign a1220 = ~a1218 & ~l180;
assign a1222 = l92 & l90;
assign a1224 = l96 & l94;
assign a1226 = a1224 & a1222;
assign a1228 = l100 & ~l98;
assign a1230 = l104 & l102;
assign a1232 = a1230 & a1228;
assign a1234 = a1232 & a1226;
assign a1236 = l108 & l106;
assign a1238 = l112 & l110;
assign a1240 = a1238 & a1236;
assign a1242 = l116 & l114;
assign a1244 = l120 & l118;
assign a1246 = a1244 & ~a1242;
assign a1248 = a1246 & a1240;
assign a1250 = a1248 & a1234;
assign a1252 = a1250 & l88;
assign a1254 = ~a1252 & l86;
assign a1256 = l122 & l84;
assign a1258 = a1256 & ~a1254;
assign a1260 = a1258 & a1206;
assign a1262 = ~a1260 & ~a1220;
assign a1264 = a1262 & a1200;
assign a1266 = ~a1264 & a1168;
assign a1268 = ~a1266 & ~a1170;
assign a1270 = ~a1268 & l64;
assign a1272 = ~l64 & ~l60;
assign a1276 = l72 & l70;
assign a1278 = l78 & ~l76;
assign a1280 = a1278 & l74;
assign a1282 = a1280 & a1276;
assign a1284 = a1282 & a1168;
assign a1286 = a1284 & l62;
assign a1288 = a1168 & ~l60;
assign a1290 = a1288 & ~a1196;
assign a1292 = ~a1290 & ~l62;
assign a1294 = ~a1292 & ~a1286;
assign a1296 = a1294 & l64;
assign a1298 = ~l64 & l62;
assign a1300 = ~a1298 & ~a1296;
assign a1304 = ~l666 & ~l660;
assign a1306 = ~l624 & ~l618;
assign a1308 = a1306 & a1304;
assign a1310 = ~l648 & ~l636;
assign a1312 = ~l654 & ~l642;
assign a1314 = a1312 & a1310;
assign a1316 = a1314 & a1308;
assign a1318 = a1316 & l758;
assign a1320 = l760 & l450;
assign a1322 = ~l764 & ~l762;
assign a1324 = a1322 & a1320;
assign a1326 = ~l768 & l766;
assign a1328 = l772 & ~l770;
assign a1330 = a1328 & a1326;
assign a1332 = a1330 & a1324;
assign a1334 = l848 & l126;
assign a1336 = l68 & ~l66;
assign a1338 = ~a1336 & ~a1334;
assign a1340 = l848 & l476;
assign a1342 = l848 & l132;
assign a1344 = ~a1342 & ~a1340;
assign a1346 = a1344 & a1338;
assign a1348 = a1346 & ~a1332;
assign a1350 = a1348 & ~a1318;
assign a1352 = l134 & l132;
assign a1354 = l138 & l136;
assign a1356 = a1354 & a1352;
assign a1358 = l180 & l152;
assign a1360 = a1358 & a1356;
assign a1362 = ~l470 & ~l158;
assign a1364 = ~a1362 & l848;
assign a1366 = ~a1196 & l866;
assign a1368 = ~a1366 & ~a1364;
assign a1370 = a1368 & ~a1360;
assign a1372 = a1316 & l114;
assign a1374 = ~l150 & l146;
assign a1376 = ~a1374 & ~a1202;
assign a1378 = l152 & ~l80;
assign a1380 = a1378 & a1376;
assign a1382 = ~l178 & ~l124;
assign a1384 = ~a1382 & l848;
assign a1386 = l848 & l128;
assign a1388 = l870 & l60;
assign a1390 = ~a1388 & ~a1386;
assign a1392 = a1390 & ~a1384;
assign a1394 = a1392 & ~a1380;
assign a1396 = a1394 & ~a1372;
assign a1398 = a1396 & a1370;
assign a1400 = a1398 & a1350;
assign a1402 = ~a1400 & l64;
assign a1404 = l68 & ~l64;
assign a1406 = ~a1404 & ~a1402;
assign a1408 = l192 & ~l190;
assign a1410 = a1408 & l64;
assign a1412 = ~l74 & ~l72;
assign a1414 = l178 & ~l70;
assign a1416 = a1414 & a1278;
assign a1418 = a1416 & a1412;
assign a1420 = a1418 & a1168;
assign a1422 = l852 & l476;
assign a1424 = a1422 & a1168;
assign a1426 = a1424 & a1252;
assign a1428 = ~a1426 & ~l178;
assign a1430 = ~a1428 & ~a1420;
assign a1432 = a1430 & ~l178;
assign a1434 = l776 & ~l774;
assign a1436 = l778 & l450;
assign a1438 = a1436 & a1434;
assign a1440 = l782 & l780;
assign a1442 = l788 & l786;
assign a1444 = a1442 & l784;
assign a1446 = a1444 & a1440;
assign a1448 = a1446 & a1438;
assign a1450 = a1448 & l790;
assign a1452 = ~a1450 & ~a1174;
assign a1454 = a1294 & ~l62;
assign a1456 = ~a1454 & a1452;
assign a1458 = a1456 & ~a1432;
assign a1460 = ~l178 & ~l62;
assign a1462 = l126 & ~l84;
assign a1464 = ~a1462 & ~l128;
assign a1466 = a1464 & a1460;
assign a1468 = a1466 & l70;
assign a1470 = ~a1466 & l72;
assign a1472 = ~a1470 & ~a1468;
assign a1474 = a1472 & a1458;
assign a1476 = ~a1474 & l64;
assign a1478 = l1166 & ~l64;
assign a1480 = ~a1478 & ~a1476;
assign a1482 = ~a1480 & ~a1410;
assign a1484 = a1410 & l70;
assign a1486 = ~a1484 & ~a1482;
assign a1488 = a1466 & l72;
assign a1490 = ~a1466 & l78;
assign a1492 = ~a1490 & ~a1488;
assign a1494 = a1492 & a1458;
assign a1496 = ~a1494 & l64;
assign a1498 = l1164 & ~l64;
assign a1500 = ~a1498 & ~a1496;
assign a1502 = ~a1500 & ~a1410;
assign a1504 = a1410 & l72;
assign a1506 = ~a1504 & ~a1502;
assign a1508 = a1466 & l74;
assign a1510 = ~l78 & l76;
assign a1512 = ~a1510 & ~a1278;
assign a1514 = ~a1512 & ~a1466;
assign a1516 = ~a1514 & ~a1508;
assign a1518 = a1516 & a1458;
assign a1520 = ~a1518 & l64;
assign a1522 = l1162 & ~l64;
assign a1524 = ~a1522 & ~a1520;
assign a1526 = ~a1524 & ~a1410;
assign a1528 = a1410 & l74;
assign a1530 = ~a1528 & ~a1526;
assign a1532 = a1466 & l76;
assign a1534 = ~a1466 & l70;
assign a1536 = ~a1534 & ~a1532;
assign a1538 = a1536 & a1458;
assign a1540 = ~a1538 & l64;
assign a1542 = l1160 & ~l64;
assign a1544 = ~a1542 & ~a1540;
assign a1546 = ~a1544 & ~a1410;
assign a1548 = a1410 & l76;
assign a1550 = ~a1548 & ~a1546;
assign a1552 = a1466 & l78;
assign a1554 = ~a1466 & l74;
assign a1556 = ~a1554 & ~a1552;
assign a1558 = a1556 & a1458;
assign a1560 = ~a1558 & l64;
assign a1562 = l1158 & ~l64;
assign a1564 = ~a1562 & ~a1560;
assign a1566 = ~a1564 & ~a1410;
assign a1568 = a1410 & l78;
assign a1570 = ~a1568 & ~a1566;
assign a1572 = ~a1168 & l182;
assign a1574 = a1174 & ~l126;
assign a1576 = ~l128 & ~l126;
assign a1578 = ~a1576 & ~l84;
assign a1580 = a1578 & a1282;
assign a1582 = ~a1580 & a1462;
assign a1584 = ~a1582 & ~a1574;
assign a1586 = ~a1584 & a1168;
assign a1588 = ~a1168 & l126;
assign a1590 = ~a1588 & ~a1586;
assign a1592 = a1590 & l126;
assign a1594 = ~a1592 & ~l182;
assign a1596 = a1218 & a1168;
assign a1598 = a1596 & ~a1194;
assign a1600 = a1598 & ~a1594;
assign a1602 = ~a1600 & ~a1572;
assign a1604 = a1602 & a1206;
assign a1606 = a1174 & a1168;
assign a1608 = a1258 & ~a1206;
assign a1610 = ~l142 & ~l140;
assign a1612 = ~a1610 & l144;
assign a1614 = a1612 & l142;
assign a1616 = a1418 & ~l176;
assign a1618 = ~a1616 & ~a1614;
assign a1620 = a1618 & ~a1608;
assign a1622 = ~a1620 & a1168;
assign a1624 = ~a1622 & ~l158;
assign a1626 = ~a1624 & ~a1606;
assign a1628 = ~a1626 & a1590;
assign a1630 = a1420 & l176;
assign a1632 = ~a1630 & ~l142;
assign a1634 = a1614 & a1168;
assign a1636 = ~a1634 & ~a1632;
assign a1638 = a1168 & l470;
assign a1640 = a1638 & a1172;
assign a1642 = ~a1640 & ~l476;
assign a1644 = ~a1642 & ~a1426;
assign a1646 = a1168 & l122;
assign a1648 = a1646 & ~l84;
assign a1650 = ~a1648 & ~l470;
assign a1652 = ~a1650 & ~a1640;
assign a1654 = ~a1652 & ~a1644;
assign a1656 = a1654 & ~a1430;
assign a1658 = a1656 & ~a1636;
assign a1660 = a1658 & a1628;
assign a1662 = ~a1660 & ~l84;
assign a1664 = ~a1662 & ~a1604;
assign a1666 = ~a1664 & l64;
assign a1668 = l80 & ~l64;
assign a1670 = ~a1668 & ~a1666;
assign a1672 = a1254 & l84;
assign a1674 = ~a1672 & a1646;
assign a1676 = ~l130 & l128;
assign a1678 = a1676 & a1580;
assign a1680 = a1356 & l84;
assign a1682 = a1612 & l140;
assign a1684 = ~a1682 & ~a1680;
assign a1686 = a1684 & ~a1678;
assign a1688 = ~a1686 & a1168;
assign a1690 = ~a1688 & ~l124;
assign a1692 = ~a1690 & ~a1674;
assign a1694 = a1692 & l84;
assign a1696 = l156 & ~l154;
assign a1698 = a1194 & ~l174;
assign a1700 = ~a1698 & l84;
assign a1702 = a1356 & a1168;
assign a1704 = ~a1286 & ~l132;
assign a1706 = ~a1704 & ~a1702;
assign a1708 = ~a1706 & ~a1294;
assign a1710 = a1708 & ~a1692;
assign a1712 = a1710 & a1268;
assign a1714 = a1712 & a1628;
assign a1716 = ~a1714 & a1700;
assign a1718 = ~a1716 & ~a1696;
assign a1720 = ~a1718 & ~a1206;
assign a1722 = ~a1720 & ~a1694;
assign a1724 = ~a1722 & l64;
assign a1726 = l82 & ~l64;
assign a1728 = ~a1726 & ~a1724;
assign a1730 = ~a1206 & l64;
assign a1732 = ~a1700 & ~a1696;
assign a1734 = ~a1732 & a1730;
assign a1736 = ~a1692 & l64;
assign a1738 = ~a1736 & l84;
assign a1740 = ~a1738 & ~a1734;
assign a1742 = ~l196 & l190;
assign a1744 = ~a1742 & l64;
assign a1746 = l872 & l326;
assign a1748 = a1746 & l458;
assign a1750 = ~a1746 & l86;
assign a1752 = ~a1750 & ~a1748;
assign a1754 = ~a1752 & l64;
assign a1756 = l1156 & ~l64;
assign a1758 = ~a1756 & ~a1754;
assign a1760 = ~a1758 & ~a1744;
assign a1762 = a1744 & l86;
assign a1764 = ~a1762 & ~a1760;
assign a1766 = l64 & i58;
assign a1768 = l88 & ~l64;
assign a1770 = ~a1768 & ~a1766;
assign a1772 = ~l476 & ~l470;
assign a1774 = ~a1772 & ~l84;
assign a1776 = ~l86 & l84;
assign a1778 = ~l1138 & ~l124;
assign a1780 = a1778 & ~a1776;
assign a1782 = a1780 & ~a1774;
assign a1784 = ~l1144 & ~l1142;
assign a1786 = a1784 & ~l1140;
assign a1788 = ~a1786 & ~a1250;
assign a1790 = a1788 & l92;
assign a1792 = ~a1790 & ~a1782;
assign a1794 = ~a1792 & l64;
assign a1796 = a1788 & l64;
assign a1798 = ~a1796 & l90;
assign a1800 = ~a1798 & ~a1794;
assign a1802 = a1788 & l96;
assign a1804 = ~a1802 & ~a1782;
assign a1806 = ~a1804 & l64;
assign a1808 = ~a1796 & l92;
assign a1810 = ~a1808 & ~a1806;
assign a1812 = a1788 & l100;
assign a1814 = ~a1812 & ~a1782;
assign a1816 = ~a1814 & l64;
assign a1818 = ~a1796 & l94;
assign a1820 = ~a1818 & ~a1816;
assign a1822 = a1788 & l112;
assign a1824 = ~a1822 & ~a1782;
assign a1826 = ~a1824 & l64;
assign a1828 = ~a1796 & l96;
assign a1830 = ~a1828 & ~a1826;
assign a1832 = a1788 & l106;
assign a1834 = ~a1832 & ~a1782;
assign a1836 = ~a1834 & l64;
assign a1838 = ~a1796 & l98;
assign a1840 = ~a1838 & ~a1836;
assign a1842 = a1788 & l90;
assign a1844 = ~a1842 & ~a1782;
assign a1846 = ~a1844 & l64;
assign a1848 = ~a1796 & l100;
assign a1850 = ~a1848 & ~a1846;
assign a1852 = a1788 & l118;
assign a1854 = ~a1852 & ~a1782;
assign a1856 = ~a1854 & l64;
assign a1858 = ~a1796 & l102;
assign a1860 = ~a1858 & ~a1856;
assign a1862 = a1788 & l120;
assign a1864 = ~a1862 & ~a1782;
assign a1866 = ~a1864 & l64;
assign a1868 = ~a1796 & l104;
assign a1870 = ~a1868 & ~a1866;
assign a1872 = a1788 & l108;
assign a1874 = ~a1872 & ~a1782;
assign a1876 = ~a1874 & l64;
assign a1878 = ~a1796 & l106;
assign a1880 = ~a1878 & ~a1876;
assign a1882 = a1788 & l102;
assign a1884 = ~a1882 & ~a1782;
assign a1886 = ~a1884 & l64;
assign a1888 = ~a1796 & l108;
assign a1890 = ~a1888 & ~a1886;
assign a1892 = a1788 & l94;
assign a1894 = ~a1892 & ~a1782;
assign a1896 = ~a1894 & l64;
assign a1898 = ~a1796 & l110;
assign a1900 = ~a1898 & ~a1896;
assign a1902 = ~l100 & l98;
assign a1904 = ~a1902 & ~a1228;
assign a1906 = ~l92 & ~l90;
assign a1908 = ~a1906 & ~a1222;
assign a1910 = a1908 & a1904;
assign a1912 = ~a1908 & ~a1904;
assign a1914 = ~a1912 & ~a1910;
assign a1916 = ~a1914 & a1788;
assign a1918 = ~a1916 & ~a1782;
assign a1920 = ~a1918 & l64;
assign a1922 = ~a1796 & l112;
assign a1924 = ~a1922 & ~a1920;
assign a1926 = l66 & l64;
assign a1928 = ~a1926 & ~l114;
assign a1930 = a1746 & l560;
assign a1932 = ~a1746 & l116;
assign a1934 = ~a1932 & ~a1930;
assign a1936 = ~a1934 & l64;
assign a1938 = l1154 & ~l64;
assign a1940 = ~a1938 & ~a1936;
assign a1942 = ~a1940 & ~a1744;
assign a1944 = a1744 & l116;
assign a1946 = ~a1944 & ~a1942;
assign a1948 = a1788 & l104;
assign a1950 = ~a1948 & ~a1782;
assign a1952 = ~a1950 & l64;
assign a1954 = ~a1796 & l118;
assign a1956 = ~a1954 & ~a1952;
assign a1958 = a1788 & l110;
assign a1960 = ~a1958 & ~a1782;
assign a1962 = ~a1960 & l64;
assign a1964 = ~a1796 & l120;
assign a1966 = ~a1964 & ~a1962;
assign a1968 = a1692 & l124;
assign a1970 = ~a1434 & ~l778;
assign a1972 = l782 & ~l84;
assign a1974 = l790 & l84;
assign a1976 = ~a1974 & ~a1972;
assign a1978 = a1976 & a1970;
assign a1980 = ~l780 & ~l774;
assign a1982 = ~a1980 & l84;
assign a1984 = ~a1982 & a1444;
assign a1986 = ~l782 & l84;
assign a1988 = l780 & l776;
assign a1990 = a1988 & l790;
assign a1992 = ~a1990 & ~l84;
assign a1994 = ~a1992 & ~a1986;
assign a1996 = a1994 & a1984;
assign a1998 = a1996 & a1978;
assign a2000 = ~a1998 & ~l122;
assign a2002 = ~a2000 & l64;
assign a2004 = a2002 & a1968;
assign a2006 = l1136 & ~l64;
assign a2008 = ~a2006 & ~a2004;
assign a2010 = ~a2008 & ~a1410;
assign a2012 = a1410 & l122;
assign a2014 = ~a2012 & ~a2010;
assign a2016 = ~l124 & ~l64;
assign a2020 = ~a1590 & l64;
assign a2022 = l126 & ~l64;
assign a2024 = ~a2022 & ~a2020;
assign a2026 = a1284 & l128;
assign a2028 = a2026 & ~l84;
assign a2030 = a2028 & l64;
assign a2032 = l790 & l64;
assign a2034 = a1168 & ~l180;
assign a2036 = a2034 & a2032;
assign a2038 = a2036 & a1448;
assign a2040 = ~a2038 & ~l128;
assign a2044 = a1746 & l462;
assign a2046 = ~a1746 & l130;
assign a2048 = ~a2046 & ~a2044;
assign a2050 = ~a2048 & l64;
assign a2052 = l1134 & ~l64;
assign a2054 = ~a2052 & ~a2050;
assign a2056 = ~a2054 & ~a1744;
assign a2058 = a1744 & l130;
assign a2060 = ~a2058 & ~a2056;
assign a2062 = a1706 & l64;
assign a2064 = l132 & ~l64;
assign a2066 = ~a2064 & ~a2062;
assign a2068 = l64 & i54;
assign a2070 = l1132 & ~l64;
assign a2072 = ~a2070 & ~a2068;
assign a2074 = ~a2072 & ~a1410;
assign a2076 = a1410 & l134;
assign a2078 = ~a2076 & ~a2074;
assign a2080 = l64 & i52;
assign a2082 = l1130 & ~l64;
assign a2084 = ~a2082 & ~a2080;
assign a2086 = ~a2084 & ~a1410;
assign a2088 = a1410 & l136;
assign a2090 = ~a2088 & ~a2086;
assign a2092 = l64 & i50;
assign a2094 = l1128 & ~l64;
assign a2096 = ~a2094 & ~a2092;
assign a2098 = ~a2096 & ~a1410;
assign a2100 = a1410 & l138;
assign a2102 = ~a2100 & ~a2098;
assign a2104 = a1168 & l64;
assign a2106 = a2104 & a1682;
assign a2108 = a2030 & l130;
assign a2110 = ~a2108 & ~l140;
assign a2114 = a1636 & l64;
assign a2116 = l142 & ~l64;
assign a2118 = ~a2116 & ~a2114;
assign a2120 = ~l1118 & l1116;
assign a2122 = l1118 & ~l1116;
assign a2124 = ~a2122 & ~a2120;
assign a2126 = l316 & l64;
assign a2128 = a2126 & l872;
assign a2130 = a2128 & ~a2124;
assign a2132 = a2130 & l424;
assign a2134 = l144 & ~l64;
assign a2136 = ~a2134 & ~a2132;
assign a2138 = a1746 & l472;
assign a2140 = ~a1746 & l146;
assign a2142 = ~a2140 & ~a2138;
assign a2144 = ~a2142 & l64;
assign a2146 = l1126 & ~l64;
assign a2148 = ~a2146 & ~a2144;
assign a2150 = ~a2148 & ~a1744;
assign a2152 = a1744 & l146;
assign a2154 = ~a2152 & ~a2150;
assign a2156 = l196 & l64;
assign a2158 = l64 & i48;
assign a2160 = l1124 & ~l64;
assign a2162 = ~a2160 & ~a2158;
assign a2164 = ~a2162 & ~a2156;
assign a2166 = a2156 & l148;
assign a2168 = ~a2166 & ~a2164;
assign a2170 = a1746 & l478;
assign a2172 = ~a1746 & l150;
assign a2174 = ~a2172 & ~a2170;
assign a2176 = ~a2174 & l64;
assign a2178 = l1122 & ~l64;
assign a2180 = ~a2178 & ~a2176;
assign a2182 = ~a2180 & ~a1744;
assign a2184 = a1744 & l150;
assign a2186 = ~a2184 & ~a2182;
assign a2188 = ~l62 & l60;
assign a2190 = ~l182 & ~l126;
assign a2192 = a2190 & ~l158;
assign a2194 = a2192 & a2188;
assign a2196 = a2194 & ~a1968;
assign a2198 = a2196 & a1664;
assign a2200 = l1108 & l64;
assign a2202 = a2200 & ~a2198;
assign a2204 = l152 & ~l64;
assign a2206 = ~a2204 & ~a2202;
assign a2208 = a1746 & l522;
assign a2210 = ~a1746 & ~l154;
assign a2212 = ~a2210 & ~a2208;
assign a2214 = ~a2212 & l64;
assign a2216 = ~l1106 & ~l64;
assign a2220 = ~a2218 & ~a1744;
assign a2222 = a1744 & ~l154;
assign a2226 = ~l126 & i44;
assign a2228 = a2226 & ~l158;
assign a2230 = a2228 & a1730;
assign a2232 = l156 & ~l64;
assign a2234 = ~a2232 & ~a2230;
assign a2236 = a1626 & l64;
assign a2238 = l158 & ~l64;
assign a2240 = ~a2238 & ~a2236;
assign a2242 = l162 & l64;
assign a2244 = l1104 & ~l64;
assign a2246 = ~a2244 & ~a2242;
assign a2248 = ~a2246 & ~a1410;
assign a2250 = a1410 & l160;
assign a2252 = ~a2250 & ~a2248;
assign a2254 = l64 & i42;
assign a2256 = l1102 & ~l64;
assign a2258 = ~a2256 & ~a2254;
assign a2260 = ~a2258 & ~a1410;
assign a2262 = a2242 & a1408;
assign a2264 = ~a2262 & ~a2260;
assign a2266 = ~a1190 & l64;
assign a2268 = l1100 & ~l64;
assign a2270 = ~a2268 & ~a2266;
assign a2272 = ~a2270 & ~a1410;
assign a2274 = l164 & l64;
assign a2276 = a2274 & a1408;
assign a2278 = ~a2276 & ~a2272;
assign a2280 = a1746 & l546;
assign a2282 = ~a1746 & l166;
assign a2284 = ~a2282 & ~a2280;
assign a2286 = ~a2284 & l64;
assign a2288 = l1098 & ~l64;
assign a2290 = ~a2288 & ~a2286;
assign a2292 = ~a2290 & ~a1744;
assign a2294 = a1744 & l166;
assign a2296 = ~a2294 & ~a2292;
assign a2298 = a1696 & l1096;
assign a2300 = ~a1698 & l168;
assign a2302 = ~a2300 & ~a2298;
assign a2304 = ~a2302 & a1730;
assign a2306 = ~a1736 & l168;
assign a2308 = ~a2306 & ~a2304;
assign a2310 = a1746 & l550;
assign a2312 = ~a1746 & l170;
assign a2314 = ~a2312 & ~a2310;
assign a2316 = ~a2314 & l64;
assign a2318 = l1094 & ~l64;
assign a2320 = ~a2318 & ~a2316;
assign a2322 = ~a2320 & ~a1744;
assign a2324 = a1744 & l170;
assign a2326 = ~a2324 & ~a2322;
assign a2328 = a2274 & ~a1182;
assign a2330 = l1092 & ~l64;
assign a2332 = ~a2330 & ~a2328;
assign a2334 = ~a2332 & ~a2156;
assign a2336 = a2156 & l172;
assign a2338 = ~a2336 & ~a2334;
assign a2340 = ~l84 & l64;
assign a2342 = l182 & ~l174;
assign a2344 = a2342 & a2340;
assign a2346 = a2344 & a1206;
assign a2348 = l1090 & ~l64;
assign a2350 = ~a2348 & ~a2346;
assign a2352 = ~a2350 & ~a1410;
assign a2354 = a1410 & l174;
assign a2356 = ~a2354 & ~a2352;
assign a2358 = a1746 & l466;
assign a2360 = ~a1746 & l176;
assign a2362 = ~a2360 & ~a2358;
assign a2364 = ~a2362 & l64;
assign a2366 = l1088 & ~l64;
assign a2368 = ~a2366 & ~a2364;
assign a2370 = ~a2368 & ~a1744;
assign a2372 = a1744 & l176;
assign a2374 = ~a2372 & ~a2370;
assign a2376 = a1430 & l64;
assign a2378 = l178 & ~l64;
assign a2380 = ~a2378 & ~a2376;
assign a2382 = ~l1074 & ~l526;
assign a2384 = l1074 & l526;
assign a2386 = ~a2384 & l60;
assign a2388 = a2386 & ~a2382;
assign a2390 = l1076 & l520;
assign a2392 = l1078 & ~l512;
assign a2394 = ~a2392 & ~a2390;
assign a2396 = ~l1076 & ~l520;
assign a2398 = ~l1078 & l512;
assign a2400 = ~a2398 & ~a2396;
assign a2402 = a2400 & a2394;
assign a2404 = a2402 & a2388;
assign a2406 = ~a2404 & ~l180;
assign a2408 = ~a2406 & l64;
assign a2410 = l1080 & ~l64;
assign a2412 = ~a2410 & ~a2408;
assign a2414 = ~a2412 & ~a1410;
assign a2416 = a1410 & l180;
assign a2418 = ~a2416 & ~a2414;
assign a2420 = ~a1602 & l64;
assign a2422 = l182 & ~l64;
assign a2424 = ~a2422 & ~a2420;
assign a2426 = ~a1208 & ~i38;
assign a2428 = ~a2426 & l64;
assign a2430 = l1072 & ~l64;
assign a2432 = ~a2430 & ~a2428;
assign a2434 = ~a2432 & ~a1410;
assign a2436 = a1410 & l184;
assign a2438 = ~a2436 & ~a2434;
assign a2440 = l186 & l182;
assign a2442 = ~a2440 & ~i36;
assign a2444 = ~a2442 & l64;
assign a2446 = l1070 & ~l64;
assign a2448 = ~a2446 & ~a2444;
assign a2450 = ~a2448 & ~a1410;
assign a2452 = a1410 & l186;
assign a2454 = ~a2452 & ~a2450;
assign a2456 = l182 & l64;
assign a2458 = a1696 & ~l188;
assign a2460 = a2458 & a2456;
assign a2462 = l194 & ~l64;
assign a2464 = ~a2462 & ~a2460;
assign a2466 = ~a2464 & ~a1410;
assign a2468 = a1410 & l188;
assign a2470 = ~a2468 & ~a2466;
assign a2472 = ~l198 & l64;
assign a2474 = l204 & ~l202;
assign a2476 = a2474 & l200;
assign a2478 = ~a2476 & l190;
assign a2480 = ~a2478 & a2472;
assign a2482 = ~l206 & ~l64;
assign a2486 = ~a2484 & ~a2156;
assign a2488 = a2156 & ~l190;
assign a2492 = ~a1696 & ~a1206;
assign a2494 = a2492 & a1270;
assign a2496 = l192 & ~l64;
assign a2498 = ~a2496 & ~a2494;
assign a2500 = l64 & i34;
assign a2502 = l1062 & ~l64;
assign a2504 = ~a2502 & ~a2500;
assign a2506 = ~a2504 & ~a2156;
assign a2508 = a2156 & l198;
assign a2510 = ~a2508 & ~a2506;
assign a2512 = ~l430 & ~l358;
assign a2514 = ~a2512 & l362;
assign a2516 = a2514 & ~l202;
assign a2518 = ~a2516 & ~l198;
assign a2520 = ~l290 & ~l288;
assign a2522 = a2520 & ~l286;
assign a2524 = ~l294 & ~l292;
assign a2526 = ~l298 & ~l296;
assign a2528 = a2526 & a2524;
assign a2530 = a2528 & a2522;
assign a2532 = ~l302 & ~l300;
assign a2534 = ~l306 & ~l304;
assign a2536 = a2534 & a2532;
assign a2538 = ~l310 & ~l308;
assign a2540 = ~l314 & ~l312;
assign a2542 = a2540 & a2538;
assign a2544 = a2542 & a2536;
assign a2546 = a2544 & a2530;
assign a2548 = ~l930 & ~l928;
assign a2550 = ~l406 & ~l326;
assign a2552 = ~l934 & ~l932;
assign a2554 = a2552 & a2550;
assign a2556 = a2554 & a2548;
assign a2558 = a2556 & a2546;
assign a2560 = l936 & l208;
assign a2562 = a2560 & l280;
assign a2564 = a2562 & ~a2558;
assign a2566 = a2564 & ~l242;
assign a2568 = ~l318 & ~l316;
assign a2570 = ~l322 & ~l320;
assign a2572 = a2570 & a2568;
assign a2574 = ~l328 & ~l326;
assign a2576 = a2574 & ~l324;
assign a2578 = ~l332 & ~l330;
assign a2580 = ~l336 & ~l334;
assign a2582 = a2580 & a2578;
assign a2584 = a2582 & a2576;
assign a2586 = a2584 & a2572;
assign a2588 = a2586 & a2546;
assign a2590 = l338 & l280;
assign a2592 = a2590 & ~l208;
assign a2594 = a2592 & ~a2588;
assign a2596 = ~a2474 & l200;
assign a2598 = a2596 & ~a2594;
assign a2600 = a2598 & ~a2566;
assign a2602 = ~a2600 & a2518;
assign a2604 = ~a2602 & l64;
assign a2606 = l1060 & ~l64;
assign a2608 = ~a2606 & ~a2604;
assign a2610 = ~a2608 & ~a2156;
assign a2612 = a2156 & l200;
assign a2614 = ~a2612 & ~a2610;
assign a2616 = l918 & l428;
assign a2618 = ~a2616 & ~l198;
assign a2620 = ~l346 & ~l202;
assign a2622 = ~a2620 & a2618;
assign a2624 = ~a2622 & l64;
assign a2626 = ~l1058 & ~l64;
assign a2630 = ~a2628 & ~a2156;
assign a2632 = a2156 & ~l202;
assign a2636 = ~l210 & ~l208;
assign a2638 = ~l214 & ~l212;
assign a2640 = a2638 & a2636;
assign a2642 = ~l220 & ~l218;
assign a2644 = a2642 & ~l216;
assign a2646 = ~l222 & l64;
assign a2648 = ~l226 & ~l224;
assign a2650 = a2648 & a2646;
assign a2652 = a2650 & a2644;
assign a2654 = a2652 & a2640;
assign a2656 = ~l230 & ~l228;
assign a2658 = ~l234 & ~l232;
assign a2660 = a2658 & a2656;
assign a2662 = ~l238 & ~l236;
assign a2664 = ~l244 & ~l242;
assign a2666 = a2664 & ~l240;
assign a2668 = a2666 & a2662;
assign a2670 = a2668 & a2660;
assign a2672 = ~l248 & ~l246;
assign a2674 = ~l252 & ~l250;
assign a2676 = a2674 & a2672;
assign a2678 = ~l256 & ~l254;
assign a2680 = ~l258 & ~l198;
assign a2682 = a2680 & a2678;
assign a2684 = a2682 & a2676;
assign a2686 = a2684 & a2670;
assign a2688 = a2686 & a2654;
assign a2690 = l260 & ~l64;
assign a2692 = ~a2690 & ~a2688;
assign a2694 = ~a2692 & ~a2156;
assign a2696 = a2156 & l204;
assign a2698 = ~a2696 & ~a2694;
assign a2700 = a2564 & l242;
assign a2702 = ~l266 & ~l264;
assign a2704 = l268 & ~l200;
assign a2706 = a2704 & ~a2702;
assign a2708 = ~a2706 & ~l256;
assign a2710 = a2708 & ~a2700;
assign a2712 = ~a2710 & l64;
assign a2714 = l1056 & ~l64;
assign a2716 = ~a2714 & ~a2712;
assign a2718 = ~a2716 & ~a1744;
assign a2720 = a1744 & l208;
assign a2722 = ~a2720 & ~a2718;
assign a2724 = l220 & l64;
assign a2726 = l1054 & ~l64;
assign a2728 = ~a2726 & ~a2724;
assign a2730 = ~a2728 & ~a1744;
assign a2732 = a1744 & l210;
assign a2734 = ~a2732 & ~a2730;
assign a2736 = l228 & l64;
assign a2738 = l1052 & ~l64;
assign a2740 = ~a2738 & ~a2736;
assign a2742 = ~a2740 & ~a1744;
assign a2744 = a1744 & l212;
assign a2746 = ~a2744 & ~a2742;
assign a2748 = l234 & l64;
assign a2750 = l1050 & ~l64;
assign a2752 = ~a2750 & ~a2748;
assign a2754 = ~a2752 & ~a1744;
assign a2756 = a1744 & l214;
assign a2758 = ~a2756 & ~a2754;
assign a2760 = l218 & l64;
assign a2762 = l1048 & ~l64;
assign a2764 = ~a2762 & ~a2760;
assign a2766 = ~a2764 & ~a1744;
assign a2768 = a1744 & l216;
assign a2770 = ~a2768 & ~a2766;
assign a2772 = l208 & l64;
assign a2774 = l1046 & ~l64;
assign a2776 = ~a2774 & ~a2772;
assign a2778 = ~a2776 & ~a1744;
assign a2780 = a1744 & l218;
assign a2782 = ~a2780 & ~a2778;
assign a2784 = l216 & l64;
assign a2786 = l1044 & ~l64;
assign a2788 = ~a2786 & ~a2784;
assign a2790 = ~a2788 & ~a1744;
assign a2792 = a1744 & l220;
assign a2794 = ~a2792 & ~a2790;
assign a2796 = l244 & l64;
assign a2798 = l1042 & ~l64;
assign a2800 = ~a2798 & ~a2796;
assign a2802 = ~a2800 & ~a1744;
assign a2804 = a1744 & l222;
assign a2806 = ~a2804 & ~a2802;
assign a2808 = l210 & l64;
assign a2810 = l1040 & ~l64;
assign a2812 = ~a2810 & ~a2808;
assign a2814 = ~a2812 & ~a1744;
assign a2816 = a1744 & l224;
assign a2818 = ~a2816 & ~a2814;
assign a2820 = l214 & l64;
assign a2822 = l1038 & ~l64;
assign a2824 = ~a2822 & ~a2820;
assign a2826 = ~a2824 & ~a1744;
assign a2828 = a1744 & l226;
assign a2830 = ~a2828 & ~a2826;
assign a2832 = l240 & l64;
assign a2834 = l1036 & ~l64;
assign a2836 = ~a2834 & ~a2832;
assign a2838 = ~a2836 & ~a1744;
assign a2840 = a1744 & l228;
assign a2842 = ~a2840 & ~a2838;
assign a2844 = l232 & l64;
assign a2846 = l1034 & ~l64;
assign a2848 = ~a2846 & ~a2844;
assign a2850 = ~a2848 & ~a1744;
assign a2852 = a1744 & l230;
assign a2854 = ~a2852 & ~a2850;
assign a2856 = l212 & l64;
assign a2858 = l1032 & ~l64;
assign a2860 = ~a2858 & ~a2856;
assign a2862 = ~a2860 & ~a1744;
assign a2864 = a1744 & l232;
assign a2866 = ~a2864 & ~a2862;
assign a2868 = l230 & l64;
assign a2870 = l1030 & ~l64;
assign a2872 = ~a2870 & ~a2868;
assign a2874 = ~a2872 & ~a1744;
assign a2876 = a1744 & l234;
assign a2878 = ~a2876 & ~a2874;
assign a2880 = l250 & l64;
assign a2882 = l1028 & ~l64;
assign a2884 = ~a2882 & ~a2880;
assign a2886 = ~a2884 & ~a1744;
assign a2888 = a1744 & l236;
assign a2890 = ~a2888 & ~a2886;
assign a2892 = l248 & l64;
assign a2894 = l1026 & ~l64;
assign a2896 = ~a2894 & ~a2892;
assign a2898 = ~a2896 & ~a1744;
assign a2900 = a1744 & l238;
assign a2902 = ~a2900 & ~a2898;
assign a2904 = l224 & l64;
assign a2906 = l1024 & ~l64;
assign a2908 = ~a2906 & ~a2904;
assign a2910 = ~a2908 & ~a1744;
assign a2912 = a1744 & l240;
assign a2914 = ~a2912 & ~a2910;
assign a2916 = a2700 & ~l256;
assign a2918 = ~a2916 & l254;
assign a2920 = a2700 & a2678;
assign a2922 = ~a2920 & ~a2918;
assign a2924 = ~a2922 & l64;
assign a2926 = l1022 & ~l64;
assign a2928 = ~a2926 & ~a2924;
assign a2930 = ~a2928 & ~a2156;
assign a2932 = a2156 & l242;
assign a2934 = ~a2932 & ~a2930;
assign a2936 = l238 & l64;
assign a2938 = l1020 & ~l64;
assign a2940 = ~a2938 & ~a2936;
assign a2942 = ~a2940 & ~a1744;
assign a2944 = a1744 & l244;
assign a2946 = ~a2944 & ~a2942;
assign a2948 = l226 & l64;
assign a2950 = l1018 & ~l64;
assign a2952 = ~a2950 & ~a2948;
assign a2954 = ~a2952 & ~a1744;
assign a2956 = a1744 & l246;
assign a2958 = ~a2956 & ~a2954;
assign a2960 = l236 & l64;
assign a2962 = l1016 & ~l64;
assign a2964 = ~a2962 & ~a2960;
assign a2966 = ~a2964 & ~a1744;
assign a2968 = a1744 & l248;
assign a2970 = ~a2968 & ~a2966;
assign a2972 = l246 & l64;
assign a2974 = l1014 & ~l64;
assign a2976 = ~a2974 & ~a2972;
assign a2978 = ~a2976 & ~a1744;
assign a2980 = a1744 & l250;
assign a2982 = ~a2980 & ~a2978;
assign a2984 = ~l1012 & ~l64;
assign a2988 = a2986 & ~a1744;
assign a2990 = a1744 & l252;
assign a2992 = ~a2990 & ~a2988;
assign a2994 = l222 & l198;
assign a2996 = a2994 & l242;
assign a2998 = a2996 & ~l270;
assign a3000 = ~a2996 & ~l258;
assign a3002 = ~a3000 & l64;
assign a3004 = a3002 & ~a2998;
assign a3006 = l1010 & ~l64;
assign a3008 = ~a3006 & ~a3004;
assign a3010 = ~a3008 & ~a2156;
assign a3012 = a2156 & l254;
assign a3014 = ~a3012 & ~a3010;
assign a3016 = a2706 & ~l256;
assign a3018 = a3016 & ~l242;
assign a3020 = l270 & ~l258;
assign a3022 = ~l270 & l258;
assign a3024 = ~a3022 & ~a3020;
assign a3026 = ~a3024 & a2994;
assign a3028 = ~a3016 & l242;
assign a3030 = ~a3028 & ~a3026;
assign a3032 = a3030 & ~a3018;
assign a3034 = ~a3032 & l64;
assign a3036 = l272 & ~l64;
assign a3038 = ~a3036 & ~a3034;
assign a3040 = ~a3038 & ~a2156;
assign a3042 = a2156 & l256;
assign a3044 = ~a3042 & ~a3040;
assign a3046 = l198 & l64;
assign a3048 = l262 & ~l64;
assign a3050 = ~a3048 & ~a3046;
assign a3052 = ~a3050 & ~a2156;
assign a3054 = a2156 & l258;
assign a3056 = ~a3054 & ~a3052;
assign a3058 = a2566 & l200;
assign a3060 = ~a3058 & ~l264;
assign a3062 = l264 & l202;
assign a3064 = ~a3062 & a2472;
assign a3066 = a3064 & ~a3060;
assign a3068 = l1008 & ~l64;
assign a3070 = ~a3068 & ~a3066;
assign a3072 = ~a3070 & ~a1744;
assign a3074 = a1744 & l264;
assign a3076 = ~a3074 & ~a3072;
assign a3078 = a2594 & l200;
assign a3080 = ~a3078 & ~l266;
assign a3082 = l342 & l340;
assign a3084 = a3082 & l266;
assign a3086 = ~a3084 & a2472;
assign a3088 = a3086 & ~a3080;
assign a3090 = l344 & ~l64;
assign a3092 = ~a3090 & ~a3088;
assign a3094 = ~a3092 & ~a1744;
assign a3096 = a1744 & l266;
assign a3098 = ~a3096 & ~a3094;
assign a3100 = l280 & l64;
assign a3102 = l282 & ~l64;
assign a3104 = ~a3102 & ~a3100;
assign a3106 = ~a3104 & ~a1744;
assign a3108 = a1744 & l268;
assign a3110 = ~a3108 & ~a3106;
assign a3112 = a3024 & l274;
assign a3114 = ~l274 & ~l198;
assign a3116 = a3114 & ~l270;
assign a3118 = ~a3116 & l64;
assign a3120 = a3118 & ~a3112;
assign a3122 = l276 & ~l64;
assign a3124 = ~a3122 & ~a3120;
assign a3126 = ~a3124 & ~a2156;
assign a3128 = a2156 & l270;
assign a3130 = ~a3128 & ~a3126;
assign a3132 = ~a3114 & a2646;
assign a3134 = l278 & ~l64;
assign a3136 = ~a3134 & ~a3132;
assign a3138 = ~a3136 & ~a2156;
assign a3140 = a2156 & l274;
assign a3142 = ~a3140 & ~a3138;
assign a3144 = a3046 & l222;
assign a3146 = l284 & ~l64;
assign a3148 = ~a3146 & ~a3144;
assign a3150 = ~a3148 & ~a1744;
assign a3152 = a1744 & l280;
assign a3154 = ~a3152 & ~a3150;
assign a3156 = l224 & ~l210;
assign a3158 = a3156 & a2994;
assign a3160 = l220 & ~l216;
assign a3162 = a3160 & a3158;
assign a3164 = a3162 & ~l208;
assign a3166 = a3164 & ~l218;
assign a3168 = l918 & l350;
assign a3170 = a3168 & a2514;
assign a3172 = ~a3170 & ~l198;
assign a3174 = a3172 & l286;
assign a3176 = ~a3174 & ~a3166;
assign a3178 = ~a3176 & l64;
assign a3180 = l1006 & ~l64;
assign a3182 = ~a3180 & ~a3178;
assign a3184 = ~a3182 & ~a1744;
assign a3186 = a1744 & l286;
assign a3188 = ~a3186 & ~a3184;
assign a3190 = a3162 & l208;
assign a3192 = a3190 & ~l218;
assign a3194 = a3172 & l288;
assign a3196 = ~a3194 & ~a3192;
assign a3198 = ~a3196 & l64;
assign a3200 = l1004 & ~l64;
assign a3202 = ~a3200 & ~a3198;
assign a3204 = ~a3202 & ~a1744;
assign a3206 = a1744 & l288;
assign a3208 = ~a3206 & ~a3204;
assign a3210 = ~l220 & l208;
assign a3212 = l218 & l216;
assign a3214 = a3212 & a3158;
assign a3216 = a3214 & a3210;
assign a3218 = a3172 & l290;
assign a3220 = ~a3218 & ~a3216;
assign a3222 = ~a3220 & l64;
assign a3224 = l1002 & ~l64;
assign a3226 = ~a3224 & ~a3222;
assign a3228 = ~a3226 & ~a1744;
assign a3230 = a1744 & l290;
assign a3232 = ~a3230 & ~a3228;
assign a3234 = a2994 & ~l224;
assign a3236 = a3234 & a2636;
assign a3238 = ~l218 & ~l216;
assign a3240 = a3238 & l220;
assign a3242 = a3240 & a3236;
assign a3244 = a3172 & l292;
assign a3246 = ~a3244 & ~a3242;
assign a3248 = ~a3246 & l64;
assign a3250 = l1000 & ~l64;
assign a3252 = ~a3250 & ~a3248;
assign a3254 = ~a3252 & ~a1744;
assign a3256 = a1744 & l292;
assign a3258 = ~a3256 & ~a3254;
assign a3260 = a3236 & a2644;
assign a3262 = a3172 & l294;
assign a3264 = ~a3262 & ~a3260;
assign a3266 = ~a3264 & l64;
assign a3268 = l998 & ~l64;
assign a3270 = ~a3268 & ~a3266;
assign a3272 = ~a3270 & ~a1744;
assign a3274 = a1744 & l294;
assign a3276 = ~a3274 & ~a3272;
assign a3278 = ~l220 & ~l208;
assign a3280 = a3278 & a3214;
assign a3282 = a3172 & l296;
assign a3284 = ~a3282 & ~a3280;
assign a3286 = ~a3284 & l64;
assign a3288 = l996 & ~l64;
assign a3290 = ~a3288 & ~a3286;
assign a3292 = ~a3290 & ~a1744;
assign a3294 = a1744 & l296;
assign a3296 = ~a3294 & ~a3292;
assign a3298 = ~l218 & l216;
assign a3300 = a3298 & l220;
assign a3302 = ~l210 & l208;
assign a3304 = a3302 & a3234;
assign a3306 = a3304 & a3300;
assign a3308 = a3172 & l298;
assign a3310 = ~a3308 & ~a3306;
assign a3312 = ~a3310 & l64;
assign a3314 = l994 & ~l64;
assign a3316 = ~a3314 & ~a3312;
assign a3318 = ~a3316 & ~a1744;
assign a3320 = a1744 & l298;
assign a3322 = ~a3320 & ~a3318;
assign a3324 = l218 & ~l216;
assign a3326 = a3324 & a3158;
assign a3328 = a3326 & a3210;
assign a3330 = a3172 & l300;
assign a3332 = ~a3330 & ~a3328;
assign a3334 = ~a3332 & l64;
assign a3336 = l992 & ~l64;
assign a3338 = ~a3336 & ~a3334;
assign a3340 = ~a3338 & ~a1744;
assign a3342 = a1744 & l300;
assign a3344 = ~a3342 & ~a3340;
assign a3346 = a3238 & a3158;
assign a3348 = a3346 & a3278;
assign a3350 = a3172 & l302;
assign a3352 = ~a3350 & ~a3348;
assign a3354 = ~a3352 & l64;
assign a3356 = l990 & ~l64;
assign a3358 = ~a3356 & ~a3354;
assign a3360 = ~a3358 & ~a1744;
assign a3362 = a1744 & l302;
assign a3364 = ~a3362 & ~a3360;
assign a3366 = a3324 & l220;
assign a3368 = a3366 & a3304;
assign a3370 = a3172 & l304;
assign a3372 = ~a3370 & ~a3368;
assign a3374 = ~a3372 & l64;
assign a3376 = l988 & ~l64;
assign a3378 = ~a3376 & ~a3374;
assign a3380 = ~a3378 & ~a1744;
assign a3382 = a1744 & l304;
assign a3384 = ~a3382 & ~a3380;
assign a3386 = ~l220 & l218;
assign a3388 = a3386 & l216;
assign a3390 = a3388 & a3304;
assign a3392 = a3172 & l306;
assign a3394 = ~a3392 & ~a3390;
assign a3396 = ~a3394 & l64;
assign a3398 = l986 & ~l64;
assign a3400 = ~a3398 & ~a3396;
assign a3402 = ~a3400 & ~a1744;
assign a3404 = a1744 & l306;
assign a3406 = ~a3404 & ~a3402;
assign a3408 = a3366 & a3236;
assign a3410 = a3172 & l308;
assign a3412 = ~a3410 & ~a3408;
assign a3414 = ~a3412 & l64;
assign a3416 = l984 & ~l64;
assign a3418 = ~a3416 & ~a3414;
assign a3420 = ~a3418 & ~a1744;
assign a3422 = a1744 & l308;
assign a3424 = ~a3422 & ~a3420;
assign a3426 = a3304 & a3240;
assign a3428 = a3172 & l310;
assign a3430 = ~a3428 & ~a3426;
assign a3432 = ~a3430 & l64;
assign a3434 = l982 & ~l64;
assign a3436 = ~a3434 & ~a3432;
assign a3438 = ~a3436 & ~a1744;
assign a3440 = a1744 & l310;
assign a3442 = ~a3440 & ~a3438;
assign a3444 = a3388 & a3236;
assign a3446 = a3172 & l312;
assign a3448 = ~a3446 & ~a3444;
assign a3450 = ~a3448 & l64;
assign a3452 = l980 & ~l64;
assign a3454 = ~a3452 & ~a3450;
assign a3456 = ~a3454 & ~a1744;
assign a3458 = a1744 & l312;
assign a3460 = ~a3458 & ~a3456;
assign a3462 = a3386 & ~l216;
assign a3464 = a3462 & a3304;
assign a3466 = a3172 & l314;
assign a3468 = ~a3466 & ~a3464;
assign a3470 = ~a3468 & l64;
assign a3472 = l978 & ~l64;
assign a3474 = ~a3472 & ~a3470;
assign a3476 = ~a3474 & ~a1744;
assign a3478 = a1744 & l314;
assign a3480 = ~a3478 & ~a3476;
assign a3482 = a3234 & l210;
assign a3484 = a3482 & a3238;
assign a3486 = a3484 & a3278;
assign a3488 = a3172 & l316;
assign a3490 = ~a3488 & ~a3486;
assign a3492 = ~a3490 & l64;
assign a3494 = l976 & ~l64;
assign a3496 = ~a3494 & ~a3492;
assign a3498 = ~a3496 & ~a1744;
assign a3500 = a1744 & l316;
assign a3502 = ~a3500 & ~a3498;
assign a3504 = a2642 & l216;
assign a3506 = a3504 & a3304;
assign a3508 = a3172 & l318;
assign a3510 = ~a3508 & ~a3506;
assign a3512 = ~a3510 & l64;
assign a3514 = l974 & ~l64;
assign a3516 = ~a3514 & ~a3512;
assign a3518 = ~a3516 & ~a1744;
assign a3520 = a1744 & l318;
assign a3522 = ~a3520 & ~a3518;
assign a3524 = a3482 & a3324;
assign a3526 = a3524 & a3210;
assign a3528 = a3172 & l320;
assign a3530 = ~a3528 & ~a3526;
assign a3532 = ~a3530 & l64;
assign a3534 = l972 & ~l64;
assign a3536 = ~a3534 & ~a3532;
assign a3538 = ~a3536 & ~a1744;
assign a3540 = a1744 & l320;
assign a3542 = ~a3540 & ~a3538;
assign a3544 = a3504 & a3236;
assign a3546 = a3172 & l322;
assign a3548 = ~a3546 & ~a3544;
assign a3550 = ~a3548 & l64;
assign a3552 = l970 & ~l64;
assign a3554 = ~a3552 & ~a3550;
assign a3556 = ~a3554 & ~a1744;
assign a3558 = a1744 & l322;
assign a3560 = ~a3558 & ~a3556;
assign a3562 = a3346 & a3210;
assign a3564 = a3172 & l324;
assign a3566 = ~a3564 & ~a3562;
assign a3568 = ~a3566 & l64;
assign a3570 = l968 & ~l64;
assign a3572 = ~a3570 & ~a3568;
assign a3574 = ~a3572 & ~a1744;
assign a3576 = a1744 & l324;
assign a3578 = ~a3576 & ~a3574;
assign a3580 = a3484 & a3210;
assign a3582 = a3172 & l326;
assign a3584 = ~a3582 & ~a3580;
assign a3586 = ~a3584 & l64;
assign a3588 = l966 & ~l64;
assign a3590 = ~a3588 & ~a3586;
assign a3592 = ~a3590 & ~a1744;
assign a3594 = a1744 & l326;
assign a3596 = ~a3594 & ~a3592;
assign a3598 = a3298 & a3158;
assign a3600 = a3598 & a3278;
assign a3602 = a3172 & l328;
assign a3604 = ~a3602 & ~a3600;
assign a3606 = ~a3604 & l64;
assign a3608 = l964 & ~l64;
assign a3610 = ~a3608 & ~a3606;
assign a3612 = ~a3610 & ~a1744;
assign a3614 = a1744 & l328;
assign a3616 = ~a3614 & ~a3612;
assign a3618 = a3598 & a3210;
assign a3620 = a3172 & l330;
assign a3622 = ~a3620 & ~a3618;
assign a3624 = ~a3622 & l64;
assign a3626 = l962 & ~l64;
assign a3628 = ~a3626 & ~a3624;
assign a3630 = ~a3628 & ~a1744;
assign a3632 = a1744 & l330;
assign a3634 = ~a3632 & ~a3630;
assign a3636 = a3326 & a3278;
assign a3638 = a3172 & l332;
assign a3640 = ~a3638 & ~a3636;
assign a3642 = ~a3640 & l64;
assign a3644 = l960 & ~l64;
assign a3646 = ~a3644 & ~a3642;
assign a3648 = ~a3646 & ~a1744;
assign a3650 = a1744 & l332;
assign a3652 = ~a3650 & ~a3648;
assign a3654 = a3304 & a2644;
assign a3656 = a3172 & l334;
assign a3658 = ~a3656 & ~a3654;
assign a3660 = ~a3658 & l64;
assign a3662 = l958 & ~l64;
assign a3664 = ~a3662 & ~a3660;
assign a3666 = ~a3664 & ~a1744;
assign a3668 = a1744 & l334;
assign a3670 = ~a3668 & ~a3666;
assign a3672 = a3462 & a3236;
assign a3674 = a3172 & l336;
assign a3676 = ~a3674 & ~a3672;
assign a3678 = ~a3676 & l64;
assign a3680 = l956 & ~l64;
assign a3682 = ~a3680 & ~a3678;
assign a3684 = ~a3682 & ~a1744;
assign a3686 = a1744 & l336;
assign a3688 = ~a3686 & ~a3684;
assign a3690 = ~l246 & i26;
assign a3692 = ~l250 & i28;
assign a3694 = ~a3692 & ~a3690;
assign a3696 = a3694 & ~a3026;
assign a3698 = ~l214 & i30;
assign a3700 = ~l226 & i32;
assign a3702 = ~a3700 & ~a3698;
assign a3704 = a2856 & l248;
assign a3706 = a3704 & a3702;
assign a3708 = a3706 & a2670;
assign a3710 = a3708 & a3696;
assign a3712 = l954 & ~l64;
assign a3714 = ~a3712 & ~a3710;
assign a3716 = ~a3714 & ~a1744;
assign a3718 = a1744 & l338;
assign a3720 = ~a3718 & ~a3716;
assign a3722 = ~l358 & ~l264;
assign a3724 = a3722 & ~l428;
assign a3726 = l202 & l64;
assign a3728 = ~l424 & ~l340;
assign a3730 = ~a3728 & a3726;
assign a3732 = a3730 & a3724;
assign a3734 = l952 & ~l64;
assign a3736 = ~a3734 & ~a3732;
assign a3738 = ~a3736 & ~a2156;
assign a3740 = a2156 & l340;
assign a3742 = ~a3740 & ~a3738;
assign a3744 = l348 & ~l346;
assign a3746 = ~l348 & l346;
assign a3748 = ~a3746 & ~a3744;
assign a3750 = ~l352 & l350;
assign a3752 = a3750 & a3748;
assign a3754 = ~a3752 & ~l342;
assign a3756 = ~a3754 & a3726;
assign a3758 = l354 & ~l64;
assign a3760 = ~a3758 & ~a3756;
assign a3762 = ~a3760 & ~a2156;
assign a3764 = a2156 & l342;
assign a3766 = ~a3764 & ~a3762;
assign a3768 = ~a2550 & l408;
assign a3770 = ~a3722 & l410;
assign a3772 = a3770 & ~a3768;
assign a3774 = l202 & l200;
assign a3776 = ~a3774 & a3722;
assign a3778 = ~a3776 & l412;
assign a3780 = ~a3778 & ~l414;
assign a3782 = a3780 & ~a3772;
assign a3784 = ~a3782 & l64;
assign a3786 = l416 & ~l64;
assign a3788 = ~a3786 & ~a3784;
assign a3790 = ~a3788 & ~a2156;
assign a3792 = a2156 & l346;
assign a3794 = ~a3792 & ~a3790;
assign a3796 = ~a3748 & l376;
assign a3798 = l348 & ~l198;
assign a3800 = a3798 & ~l376;
assign a3802 = ~a3800 & ~a3796;
assign a3804 = ~a3802 & l64;
assign a3806 = l404 & ~l64;
assign a3808 = ~a3806 & ~a3804;
assign a3810 = ~a3808 & ~a2156;
assign a3812 = a2156 & l348;
assign a3814 = ~a3812 & ~a3810;
assign a3816 = l372 & ~l370;
assign a3818 = l376 & l374;
assign a3820 = a3818 & a3816;
assign a3822 = ~l380 & ~l378;
assign a3824 = l384 & l382;
assign a3826 = a3824 & a3822;
assign a3828 = a3826 & a3820;
assign a3830 = ~l350 & l64;
assign a3832 = a3830 & ~l198;
assign a3834 = a3832 & a3828;
assign a3836 = l386 & ~l64;
assign a3838 = ~a3836 & ~a3834;
assign a3840 = ~a3838 & ~a2156;
assign a3842 = a2156 & l350;
assign a3844 = ~a3842 & ~a3840;
assign a3846 = a3722 & l350;
assign a3848 = a3846 & ~a3748;
assign a3850 = ~a3848 & ~l356;
assign a3852 = a3848 & l356;
assign a3854 = ~a3852 & ~a3850;
assign a3856 = ~a3854 & l348;
assign a3858 = a3854 & ~l348;
assign a3860 = ~a3858 & ~a3856;
assign a3862 = ~a3860 & l350;
assign a3864 = ~l350 & l346;
assign a3866 = ~a3864 & ~a3862;
assign a3868 = ~a3866 & l64;
assign a3870 = l360 & ~l64;
assign a3872 = ~a3870 & ~a3868;
assign a3874 = ~a3872 & ~a2156;
assign a3876 = a2156 & l352;
assign a3878 = ~a3876 & ~a3874;
assign a3880 = a3830 & l356;
assign a3882 = l368 & ~l64;
assign a3884 = ~a3882 & ~a3880;
assign a3886 = ~a3884 & ~a1744;
assign a3888 = a1744 & l356;
assign a3890 = ~a3888 & ~a3886;
assign a3892 = ~a3062 & ~l358;
assign a3894 = l362 & ~l202;
assign a3896 = a3894 & l358;
assign a3898 = ~a3896 & a2472;
assign a3900 = a3898 & ~a3892;
assign a3902 = l364 & ~l64;
assign a3904 = ~a3902 & ~a3900;
assign a3906 = ~a3904 & ~a1744;
assign a3908 = a1744 & l358;
assign a3910 = ~a3908 & ~a3906;
assign a3912 = l64 & i4;
assign a3914 = a3912 & i2;
assign a3916 = l366 & ~l64;
assign a3918 = ~a3916 & ~a3914;
assign a3920 = ~a3918 & ~a2156;
assign a3922 = a2156 & l362;
assign a3924 = ~a3922 & ~a3920;
assign a3926 = l402 & ~l64;
assign a3928 = a3726 & l380;
assign a3930 = ~a3928 & ~a3926;
assign a3932 = a3930 & ~a2156;
assign a3934 = a2156 & ~l370;
assign a3938 = ~l372 & l370;
assign a3940 = ~a3938 & l202;
assign a3942 = a3940 & ~a3816;
assign a3944 = ~a3942 & l64;
assign a3946 = ~l400 & ~l64;
assign a3950 = ~a3948 & ~a2156;
assign a3952 = a2156 & ~l372;
assign a3956 = l398 & ~l64;
assign a3958 = a3726 & l382;
assign a3960 = ~a3958 & ~a3956;
assign a3962 = a3960 & ~a2156;
assign a3964 = a2156 & ~l374;
assign a3968 = l346 & ~l202;
assign a3970 = ~a3968 & ~l376;
assign a3972 = ~a3970 & a2472;
assign a3974 = a3972 & ~a3828;
assign a3976 = l396 & ~l64;
assign a3978 = ~a3976 & ~a3974;
assign a3980 = ~a3978 & ~a2156;
assign a3982 = a2156 & l376;
assign a3984 = ~a3982 & ~a3980;
assign a3986 = l394 & ~l64;
assign a3988 = a3726 & l384;
assign a3990 = ~a3988 & ~a3986;
assign a3992 = a3990 & ~a2156;
assign a3994 = a2156 & ~l378;
assign a3998 = l392 & ~l64;
assign a4000 = a3726 & l378;
assign a4002 = ~a4000 & ~a3998;
assign a4004 = a4002 & ~a2156;
assign a4006 = a2156 & ~l380;
assign a4010 = l390 & ~l64;
assign a4012 = a3726 & l372;
assign a4014 = ~a4012 & ~a4010;
assign a4016 = a4014 & ~a2156;
assign a4018 = a2156 & ~l382;
assign a4022 = l388 & ~l64;
assign a4024 = a3726 & l374;
assign a4026 = ~a4024 & ~a4022;
assign a4028 = a4026 & ~a2156;
assign a4030 = a2156 & ~l384;
assign a4034 = a3524 & a3278;
assign a4036 = a3172 & l406;
assign a4038 = ~a4036 & ~a4034;
assign a4040 = ~a4038 & l64;
assign a4042 = l950 & ~l64;
assign a4044 = ~a4042 & ~a4040;
assign a4046 = ~a4044 & ~a1744;
assign a4048 = a1744 & l406;
assign a4050 = ~a4048 & ~a4046;
assign a4052 = ~a3058 & ~l408;
assign a4054 = ~a3768 & l64;
assign a4056 = a4054 & a2618;
assign a4058 = a4056 & ~a4052;
assign a4060 = l938 & ~l64;
assign a4062 = ~a4060 & ~a4058;
assign a4064 = ~a4062 & ~a1744;
assign a4066 = a1744 & l408;
assign a4068 = ~a4066 & ~a4064;
assign a4070 = ~l422 & ~l64;
assign a4072 = a4054 & ~l424;
assign a4076 = a4074 & ~a1744;
assign a4078 = a1744 & l410;
assign a4080 = ~a4078 & ~a4076;
assign a4082 = ~i10 & ~i8;
assign a4084 = ~a4082 & l64;
assign a4086 = l420 & ~l64;
assign a4088 = ~a4086 & ~a4084;
assign a4090 = ~a4088 & ~a2156;
assign a4092 = a2156 & l412;
assign a4094 = ~a4092 & ~a4090;
assign a4096 = l64 & i6;
assign a4098 = l418 & ~l64;
assign a4100 = ~a4098 & ~a4096;
assign a4102 = ~a4100 & ~a2156;
assign a4104 = a2156 & l414;
assign a4106 = ~a4104 & ~a4102;
assign a4108 = l426 & l326;
assign a4110 = l406 & ~l60;
assign a4112 = ~a4110 & ~a4108;
assign a4114 = ~a4112 & a3768;
assign a4116 = l424 & l340;
assign a4118 = l430 & l428;
assign a4120 = ~a4118 & ~l340;
assign a4122 = a4120 & l432;
assign a4124 = ~a4122 & ~a4116;
assign a4126 = ~a4124 & ~a3768;
assign a4128 = ~a4126 & ~a4114;
assign a4130 = ~a4128 & l64;
assign a4132 = l434 & ~l64;
assign a4134 = ~a4132 & ~a4130;
assign a4136 = ~a4134 & ~a1744;
assign a4138 = a1744 & l424;
assign a4140 = ~a4138 & ~a4136;
assign a4142 = a1746 & l424;
assign a4144 = ~a1746 & l426;
assign a4146 = ~a4144 & ~a4142;
assign a4148 = ~a4146 & l64;
assign a4150 = l926 & ~l64;
assign a4152 = ~a4150 & ~a4148;
assign a4154 = ~a4152 & ~a1744;
assign a4156 = a1744 & l426;
assign a4158 = ~a4156 & ~a4154;
assign a4160 = a3938 & ~l382;
assign a4162 = ~l384 & ~l374;
assign a4164 = a4162 & a3822;
assign a4166 = a4164 & a4160;
assign a4168 = a3082 & l876;
assign a4170 = ~a4168 & a3722;
assign a4172 = a4170 & ~a4166;
assign a4174 = ~a4172 & l916;
assign a4176 = ~a4174 & ~l428;
assign a4178 = ~a2616 & a2472;
assign a4180 = a4178 & ~a4176;
assign a4182 = l920 & ~l64;
assign a4184 = ~a4182 & ~a4180;
assign a4186 = ~a4184 & ~a2156;
assign a4188 = a2156 & l428;
assign a4190 = ~a4188 & ~a4186;
assign a4192 = ~a3084 & ~l430;
assign a4194 = a3894 & l430;
assign a4196 = ~a4194 & a2472;
assign a4198 = a4196 & ~a4192;
assign a4200 = l914 & ~l64;
assign a4202 = ~a4200 & ~a4198;
assign a4204 = ~a4202 & ~a1744;
assign a4206 = a1744 & l430;
assign a4208 = ~a4206 & ~a4204;
assign a4210 = l436 & l326;
assign a4212 = l406 & l62;
assign a4214 = ~a4212 & ~a4210;
assign a4216 = ~a4214 & a3768;
assign a4218 = l432 & l340;
assign a4220 = a4120 & l438;
assign a4222 = ~a4220 & ~a4218;
assign a4224 = ~a4222 & ~a3768;
assign a4226 = ~a4224 & ~a4216;
assign a4228 = ~a4226 & l64;
assign a4230 = l440 & ~l64;
assign a4232 = ~a4230 & ~a4228;
assign a4234 = ~a4232 & ~a1744;
assign a4236 = a1744 & l432;
assign a4238 = ~a4236 & ~a4234;
assign a4240 = a1746 & l432;
assign a4242 = ~a1746 & l436;
assign a4244 = ~a4242 & ~a4240;
assign a4246 = ~a4244 & l64;
assign a4248 = l912 & ~l64;
assign a4250 = ~a4248 & ~a4246;
assign a4252 = ~a4250 & ~a1744;
assign a4254 = a1744 & l436;
assign a4256 = ~a4254 & ~a4252;
assign a4258 = l442 & l326;
assign a4260 = l406 & l132;
assign a4262 = ~a4260 & ~a4258;
assign a4264 = ~a4262 & a3768;
assign a4266 = l438 & l340;
assign a4268 = a4120 & l444;
assign a4270 = ~a4268 & ~a4266;
assign a4272 = ~a4270 & ~a3768;
assign a4274 = ~a4272 & ~a4264;
assign a4276 = ~a4274 & l64;
assign a4278 = l446 & ~l64;
assign a4280 = ~a4278 & ~a4276;
assign a4282 = ~a4280 & ~a1744;
assign a4284 = a1744 & l438;
assign a4286 = ~a4284 & ~a4282;
assign a4288 = a1746 & l438;
assign a4290 = ~a1746 & l442;
assign a4292 = ~a4290 & ~a4288;
assign a4294 = ~a4292 & l64;
assign a4296 = l910 & ~l64;
assign a4298 = ~a4296 & ~a4294;
assign a4300 = ~a4298 & ~a1744;
assign a4302 = a1744 & l442;
assign a4304 = ~a4302 & ~a4300;
assign a4306 = l448 & l326;
assign a4308 = l450 & l406;
assign a4310 = ~a4308 & ~a4306;
assign a4312 = ~a4310 & a3768;
assign a4314 = l444 & l340;
assign a4316 = a4120 & l452;
assign a4318 = ~a4316 & ~a4314;
assign a4320 = ~a4318 & ~a3768;
assign a4322 = ~a4320 & ~a4312;
assign a4324 = ~a4322 & l64;
assign a4326 = l454 & ~l64;
assign a4328 = ~a4326 & ~a4324;
assign a4330 = ~a4328 & ~a1744;
assign a4332 = a1744 & l444;
assign a4334 = ~a4332 & ~a4330;
assign a4336 = a1746 & l444;
assign a4338 = ~a1746 & l448;
assign a4340 = ~a4338 & ~a4336;
assign a4342 = ~a4340 & l64;
assign a4344 = l908 & ~l64;
assign a4346 = ~a4344 & ~a4342;
assign a4348 = ~a4346 & ~a1744;
assign a4350 = a1744 & l448;
assign a4352 = ~a4350 & ~a4348;
assign a4354 = a1450 & a1168;
assign a4356 = a1702 & ~l84;
assign a4358 = ~a4356 & ~l450;
assign a4360 = ~a4358 & ~a4354;
assign a4362 = a4360 & l64;
assign a4364 = l450 & ~l64;
assign a4366 = ~a4364 & ~a4362;
assign a4368 = l456 & l326;
assign a4370 = l406 & l128;
assign a4372 = ~a4370 & ~a4368;
assign a4374 = ~a4372 & a3768;
assign a4376 = l452 & l340;
assign a4378 = a4120 & l458;
assign a4380 = ~a4378 & ~a4376;
assign a4382 = ~a4380 & ~a3768;
assign a4384 = ~a4382 & ~a4374;
assign a4386 = ~a4384 & l64;
assign a4388 = l460 & ~l64;
assign a4390 = ~a4388 & ~a4386;
assign a4392 = ~a4390 & ~a1744;
assign a4394 = a1744 & l452;
assign a4396 = ~a4394 & ~a4392;
assign a4398 = a1746 & l452;
assign a4400 = ~a1746 & l456;
assign a4402 = ~a4400 & ~a4398;
assign a4404 = ~a4402 & l64;
assign a4406 = l906 & ~l64;
assign a4408 = ~a4406 & ~a4404;
assign a4410 = ~a4408 & ~a1744;
assign a4412 = a1744 & l456;
assign a4414 = ~a4412 & ~a4410;
assign a4416 = l326 & l86;
assign a4418 = l406 & l140;
assign a4420 = ~a4418 & ~a4416;
assign a4422 = ~a4420 & a3768;
assign a4424 = l458 & l340;
assign a4426 = a4120 & l462;
assign a4428 = ~a4426 & ~a4424;
assign a4430 = ~a4428 & ~a3768;
assign a4432 = ~a4430 & ~a4422;
assign a4434 = ~a4432 & l64;
assign a4436 = l464 & ~l64;
assign a4438 = ~a4436 & ~a4434;
assign a4440 = ~a4438 & ~a1744;
assign a4442 = a1744 & l458;
assign a4444 = ~a4442 & ~a4440;
assign a4446 = l326 & l130;
assign a4448 = l406 & l124;
assign a4450 = ~a4448 & ~a4446;
assign a4452 = ~a4450 & a3768;
assign a4454 = l462 & l340;
assign a4456 = a4120 & l466;
assign a4458 = ~a4456 & ~a4454;
assign a4460 = ~a4458 & ~a3768;
assign a4462 = ~a4460 & ~a4452;
assign a4464 = ~a4462 & l64;
assign a4466 = l468 & ~l64;
assign a4468 = ~a4466 & ~a4464;
assign a4470 = ~a4468 & ~a1744;
assign a4472 = a1744 & l462;
assign a4474 = ~a4472 & ~a4470;
assign a4476 = l326 & l176;
assign a4478 = l470 & l406;
assign a4480 = ~a4478 & ~a4476;
assign a4482 = ~a4480 & a3768;
assign a4484 = l466 & l340;
assign a4486 = a4120 & l472;
assign a4488 = ~a4486 & ~a4484;
assign a4490 = ~a4488 & ~a3768;
assign a4492 = ~a4490 & ~a4482;
assign a4494 = ~a4492 & l64;
assign a4496 = l474 & ~l64;
assign a4498 = ~a4496 & ~a4494;
assign a4500 = ~a4498 & ~a1744;
assign a4502 = a1744 & l466;
assign a4504 = ~a4502 & ~a4500;
assign a4506 = a1652 & l64;
assign a4508 = l470 & ~l64;
assign a4510 = ~a4508 & ~a4506;
assign a4512 = l326 & l146;
assign a4514 = l476 & l406;
assign a4516 = ~a4514 & ~a4512;
assign a4518 = ~a4516 & a3768;
assign a4520 = l472 & l340;
assign a4522 = a4120 & l478;
assign a4524 = ~a4522 & ~a4520;
assign a4526 = ~a4524 & ~a3768;
assign a4528 = ~a4526 & ~a4518;
assign a4530 = ~a4528 & l64;
assign a4532 = l480 & ~l64;
assign a4534 = ~a4532 & ~a4530;
assign a4536 = ~a4534 & ~a1744;
assign a4538 = a1744 & l472;
assign a4540 = ~a4538 & ~a4536;
assign a4542 = a1644 & l64;
assign a4544 = l476 & ~l64;
assign a4546 = ~a4544 & ~a4542;
assign a4548 = l326 & l150;
assign a4550 = l406 & l178;
assign a4552 = ~a4550 & ~a4548;
assign a4554 = ~a4552 & a3768;
assign a4556 = l478 & l340;
assign a4558 = a4120 & l482;
assign a4560 = ~a4558 & ~a4556;
assign a4562 = ~a4560 & ~a3768;
assign a4564 = ~a4562 & ~a4554;
assign a4566 = ~a4564 & l64;
assign a4568 = l484 & ~l64;
assign a4570 = ~a4568 & ~a4566;
assign a4572 = ~a4570 & ~a1744;
assign a4574 = a1744 & l478;
assign a4576 = ~a4574 & ~a4572;
assign a4578 = l486 & l326;
assign a4580 = l406 & l142;
assign a4582 = ~a4580 & ~a4578;
assign a4584 = ~a4582 & a3768;
assign a4586 = l482 & l340;
assign a4588 = a4120 & l488;
assign a4590 = ~a4588 & ~a4586;
assign a4592 = ~a4590 & ~a3768;
assign a4594 = ~a4592 & ~a4584;
assign a4596 = ~a4594 & l64;
assign a4598 = l490 & ~l64;
assign a4600 = ~a4598 & ~a4596;
assign a4602 = ~a4600 & ~a1744;
assign a4604 = a1744 & l482;
assign a4606 = ~a4604 & ~a4602;
assign a4608 = a1746 & l482;
assign a4610 = ~a1746 & l486;
assign a4612 = ~a4610 & ~a4608;
assign a4614 = ~a4612 & l64;
assign a4616 = l904 & ~l64;
assign a4618 = ~a4616 & ~a4614;
assign a4620 = ~a4618 & ~a1744;
assign a4622 = a1744 & l486;
assign a4624 = ~a4622 & ~a4620;
assign a4626 = l492 & l326;
assign a4628 = l406 & l158;
assign a4630 = ~a4628 & ~a4626;
assign a4632 = ~a4630 & a3768;
assign a4634 = l488 & l340;
assign a4636 = a4120 & l494;
assign a4638 = ~a4636 & ~a4634;
assign a4640 = ~a4638 & ~a3768;
assign a4642 = ~a4640 & ~a4632;
assign a4644 = ~a4642 & l64;
assign a4646 = l496 & ~l64;
assign a4648 = ~a4646 & ~a4644;
assign a4650 = ~a4648 & ~a1744;
assign a4652 = a1744 & l488;
assign a4654 = ~a4652 & ~a4650;
assign a4656 = a1746 & l488;
assign a4658 = ~a1746 & l492;
assign a4660 = ~a4658 & ~a4656;
assign a4662 = ~a4660 & l64;
assign a4664 = l902 & ~l64;
assign a4666 = ~a4664 & ~a4662;
assign a4668 = ~a4666 & ~a1744;
assign a4670 = a1744 & l492;
assign a4672 = ~a4670 & ~a4668;
assign a4674 = l498 & l326;
assign a4676 = l406 & l126;
assign a4678 = ~a4676 & ~a4674;
assign a4680 = ~a4678 & a3768;
assign a4682 = l494 & l340;
assign a4684 = a4120 & l500;
assign a4686 = ~a4684 & ~a4682;
assign a4688 = ~a4686 & ~a3768;
assign a4690 = ~a4688 & ~a4680;
assign a4692 = ~a4690 & l64;
assign a4694 = l502 & ~l64;
assign a4696 = ~a4694 & ~a4692;
assign a4698 = ~a4696 & ~a1744;
assign a4700 = a1744 & l494;
assign a4702 = ~a4700 & ~a4698;
assign a4704 = a1746 & l494;
assign a4706 = ~a1746 & l498;
assign a4708 = ~a4706 & ~a4704;
assign a4710 = ~a4708 & l64;
assign a4712 = l900 & ~l64;
assign a4714 = ~a4712 & ~a4710;
assign a4716 = ~a4714 & ~a1744;
assign a4718 = a1744 & l498;
assign a4720 = ~a4718 & ~a4716;
assign a4722 = l504 & l326;
assign a4724 = l406 & l182;
assign a4726 = ~a4724 & ~a4722;
assign a4728 = ~a4726 & a3768;
assign a4730 = l500 & l340;
assign a4732 = a4120 & l506;
assign a4734 = ~a4732 & ~a4730;
assign a4736 = ~a4734 & ~a3768;
assign a4738 = ~a4736 & ~a4728;
assign a4740 = ~a4738 & l64;
assign a4742 = l508 & ~l64;
assign a4744 = ~a4742 & ~a4740;
assign a4746 = ~a4744 & ~a1744;
assign a4748 = a1744 & l500;
assign a4750 = ~a4748 & ~a4746;
assign a4752 = a1746 & l500;
assign a4754 = ~a1746 & l504;
assign a4756 = ~a4754 & ~a4752;
assign a4758 = ~a4756 & l64;
assign a4760 = l898 & ~l64;
assign a4762 = ~a4760 & ~a4758;
assign a4764 = ~a4762 & ~a1744;
assign a4766 = a1744 & l504;
assign a4768 = ~a4766 & ~a4764;
assign a4770 = l510 & l326;
assign a4772 = l512 & l406;
assign a4774 = ~a4772 & ~a4770;
assign a4776 = ~a4774 & a3768;
assign a4778 = l506 & l340;
assign a4780 = a4120 & l514;
assign a4782 = ~a4780 & ~a4778;
assign a4784 = ~a4782 & ~a3768;
assign a4786 = ~a4784 & ~a4776;
assign a4788 = ~a4786 & l64;
assign a4790 = l516 & ~l64;
assign a4792 = ~a4790 & ~a4788;
assign a4794 = ~a4792 & ~a1744;
assign a4796 = a1744 & l506;
assign a4798 = ~a4796 & ~a4794;
assign a4800 = a1746 & l506;
assign a4802 = ~a1746 & l510;
assign a4804 = ~a4802 & ~a4800;
assign a4806 = ~a4804 & l64;
assign a4808 = l896 & ~l64;
assign a4810 = ~a4808 & ~a4806;
assign a4812 = ~a4810 & ~a1744;
assign a4814 = a1744 & l510;
assign a4816 = ~a4814 & ~a4812;
assign a4818 = l872 & l320;
assign a4820 = a4818 & l424;
assign a4822 = ~a4818 & l512;
assign a4824 = ~a4822 & ~a4820;
assign a4826 = ~a4824 & l64;
assign a4828 = l894 & ~l64;
assign a4830 = ~a4828 & ~a4826;
assign a4832 = ~a4830 & ~a1744;
assign a4834 = a1744 & l512;
assign a4836 = ~a4834 & ~a4832;
assign a4838 = l518 & l326;
assign a4840 = ~l520 & l406;
assign a4842 = ~a4840 & ~a4838;
assign a4844 = ~a4842 & a3768;
assign a4846 = l514 & l340;
assign a4848 = a4120 & l522;
assign a4850 = ~a4848 & ~a4846;
assign a4852 = ~a4850 & ~a3768;
assign a4854 = ~a4852 & ~a4844;
assign a4856 = ~a4854 & l64;
assign a4858 = l524 & ~l64;
assign a4860 = ~a4858 & ~a4856;
assign a4862 = ~a4860 & ~a1744;
assign a4864 = a1744 & l514;
assign a4866 = ~a4864 & ~a4862;
assign a4868 = a1746 & l514;
assign a4870 = ~a1746 & l518;
assign a4872 = ~a4870 & ~a4868;
assign a4874 = ~a4872 & l64;
assign a4876 = l892 & ~l64;
assign a4878 = ~a4876 & ~a4874;
assign a4880 = ~a4878 & ~a1744;
assign a4882 = a1744 & l518;
assign a4884 = ~a4882 & ~a4880;
assign a4886 = a4818 & l432;
assign a4888 = ~a4818 & ~l520;
assign a4890 = ~a4888 & ~a4886;
assign a4892 = ~a4890 & l64;
assign a4894 = ~l890 & ~l64;
assign a4898 = ~a4896 & ~a1744;
assign a4900 = a1744 & ~l520;
assign a4904 = l326 & ~l154;
assign a4906 = ~l526 & l406;
assign a4908 = ~a4906 & ~a4904;
assign a4910 = ~a4908 & a3768;
assign a4912 = l522 & l340;
assign a4914 = a4120 & l528;
assign a4916 = ~a4914 & ~a4912;
assign a4918 = ~a4916 & ~a3768;
assign a4920 = ~a4918 & ~a4910;
assign a4922 = ~a4920 & l64;
assign a4924 = l530 & ~l64;
assign a4926 = ~a4924 & ~a4922;
assign a4928 = ~a4926 & ~a1744;
assign a4930 = a1744 & l522;
assign a4932 = ~a4930 & ~a4928;
assign a4934 = a4818 & l438;
assign a4936 = ~a4818 & ~l526;
assign a4938 = ~a4936 & ~a4934;
assign a4940 = ~a4938 & l64;
assign a4942 = ~l888 & ~l64;
assign a4946 = ~a4944 & ~a1744;
assign a4948 = a1744 & ~l526;
assign a4952 = a3768 & l326;
assign a4954 = a4952 & l532;
assign a4956 = l528 & l340;
assign a4958 = a4120 & l534;
assign a4960 = ~a4958 & ~a4956;
assign a4962 = ~a4960 & ~a3768;
assign a4964 = ~a4962 & ~a4954;
assign a4966 = ~a4964 & l64;
assign a4968 = l536 & ~l64;
assign a4970 = ~a4968 & ~a4966;
assign a4972 = ~a4970 & ~a1744;
assign a4974 = a1744 & l528;
assign a4976 = ~a4974 & ~a4972;
assign a4978 = a1746 & l528;
assign a4980 = ~a1746 & l532;
assign a4982 = ~a4980 & ~a4978;
assign a4984 = ~a4982 & l64;
assign a4986 = l886 & ~l64;
assign a4988 = ~a4986 & ~a4984;
assign a4990 = ~a4988 & ~a1744;
assign a4992 = a1744 & l532;
assign a4994 = ~a4992 & ~a4990;
assign a4996 = a4952 & l538;
assign a4998 = l534 & l340;
assign a5000 = a4120 & l540;
assign a5002 = ~a5000 & ~a4998;
assign a5004 = ~a5002 & ~a3768;
assign a5006 = ~a5004 & ~a4996;
assign a5008 = ~a5006 & l64;
assign a5010 = l542 & ~l64;
assign a5012 = ~a5010 & ~a5008;
assign a5014 = ~a5012 & ~a1744;
assign a5016 = a1744 & l534;
assign a5018 = ~a5016 & ~a5014;
assign a5020 = a1746 & l534;
assign a5022 = ~a1746 & l538;
assign a5024 = ~a5022 & ~a5020;
assign a5026 = ~a5024 & l64;
assign a5028 = l884 & ~l64;
assign a5030 = ~a5028 & ~a5026;
assign a5032 = ~a5030 & ~a1744;
assign a5034 = a1744 & l538;
assign a5036 = ~a5034 & ~a5032;
assign a5038 = a4952 & l544;
assign a5040 = l540 & l340;
assign a5042 = a4120 & l546;
assign a5044 = ~a5042 & ~a5040;
assign a5046 = ~a5044 & ~a3768;
assign a5048 = ~a5046 & ~a5038;
assign a5050 = ~a5048 & l64;
assign a5052 = l548 & ~l64;
assign a5054 = ~a5052 & ~a5050;
assign a5056 = ~a5054 & ~a1744;
assign a5058 = a1744 & l540;
assign a5060 = ~a5058 & ~a5056;
assign a5062 = a1746 & l540;
assign a5064 = ~a1746 & l544;
assign a5066 = ~a5064 & ~a5062;
assign a5068 = ~a5066 & l64;
assign a5070 = l882 & ~l64;
assign a5072 = ~a5070 & ~a5068;
assign a5074 = ~a5072 & ~a1744;
assign a5076 = a1744 & l544;
assign a5078 = ~a5076 & ~a5074;
assign a5080 = a4952 & l166;
assign a5082 = l546 & l340;
assign a5084 = a4120 & l550;
assign a5086 = ~a5084 & ~a5082;
assign a5088 = ~a5086 & ~a3768;
assign a5090 = ~a5088 & ~a5080;
assign a5092 = ~a5090 & l64;
assign a5094 = l552 & ~l64;
assign a5096 = ~a5094 & ~a5092;
assign a5098 = ~a5096 & ~a1744;
assign a5100 = a1744 & l546;
assign a5102 = ~a5100 & ~a5098;
assign a5104 = a4952 & l170;
assign a5106 = l550 & l340;
assign a5108 = a4120 & l554;
assign a5110 = ~a5108 & ~a5106;
assign a5112 = ~a5110 & ~a3768;
assign a5114 = ~a5112 & ~a5104;
assign a5116 = ~a5114 & l64;
assign a5118 = l556 & ~l64;
assign a5120 = ~a5118 & ~a5116;
assign a5122 = ~a5120 & ~a1744;
assign a5124 = a1744 & l550;
assign a5126 = ~a5124 & ~a5122;
assign a5128 = a4952 & l558;
assign a5130 = l554 & l340;
assign a5132 = a4120 & l560;
assign a5134 = ~a5132 & ~a5130;
assign a5136 = ~a5134 & ~a3768;
assign a5138 = ~a5136 & ~a5128;
assign a5140 = ~a5138 & l64;
assign a5142 = l562 & ~l64;
assign a5144 = ~a5142 & ~a5140;
assign a5146 = ~a5144 & ~a1744;
assign a5148 = a1744 & l554;
assign a5150 = ~a5148 & ~a5146;
assign a5152 = a1746 & l554;
assign a5154 = ~a1746 & l558;
assign a5156 = ~a5154 & ~a5152;
assign a5158 = ~a5156 & l64;
assign a5160 = l874 & ~l64;
assign a5162 = ~a5160 & ~a5158;
assign a5164 = ~a5162 & ~a1744;
assign a5166 = a1744 & l558;
assign a5168 = ~a5166 & ~a5164;
assign a5170 = a4952 & l116;
assign a5172 = l560 & l340;
assign a5174 = a4120 & l564;
assign a5176 = ~a5174 & ~a5172;
assign a5178 = ~a5176 & ~a3768;
assign a5180 = ~a5178 & ~a5170;
assign a5182 = ~a5180 & l64;
assign a5184 = l566 & ~l64;
assign a5186 = ~a5184 & ~a5182;
assign a5188 = ~a5186 & ~a1744;
assign a5190 = a1744 & l560;
assign a5192 = ~a5190 & ~a5188;
assign a5194 = l564 & l340;
assign a5196 = a4120 & l568;
assign a5198 = ~a5196 & ~a5194;
assign a5200 = ~a5198 & a4054;
assign a5202 = l570 & ~l64;
assign a5204 = ~a5202 & ~a5200;
assign a5206 = ~a5204 & ~a1744;
assign a5208 = a1744 & l564;
assign a5210 = ~a5208 & ~a5206;
assign a5212 = l568 & l340;
assign a5214 = a4120 & l572;
assign a5216 = ~a5214 & ~a5212;
assign a5218 = ~a5216 & a4054;
assign a5220 = l574 & ~l64;
assign a5222 = ~a5220 & ~a5218;
assign a5224 = ~a5222 & ~a1744;
assign a5226 = a1744 & l568;
assign a5228 = ~a5226 & ~a5224;
assign a5230 = l572 & l340;
assign a5232 = a4120 & l576;
assign a5234 = ~a5232 & ~a5230;
assign a5236 = ~a5234 & a4054;
assign a5238 = l578 & ~l64;
assign a5240 = ~a5238 & ~a5236;
assign a5242 = ~a5240 & ~a1744;
assign a5244 = a1744 & l572;
assign a5246 = ~a5244 & ~a5242;
assign a5248 = l576 & l340;
assign a5250 = a4120 & l580;
assign a5252 = ~a5250 & ~a5248;
assign a5254 = ~a5252 & a4054;
assign a5256 = l582 & ~l64;
assign a5258 = ~a5256 & ~a5254;
assign a5260 = ~a5258 & ~a1744;
assign a5262 = a1744 & l576;
assign a5264 = ~a5262 & ~a5260;
assign a5266 = l580 & l340;
assign a5268 = a4120 & l584;
assign a5270 = ~a5268 & ~a5266;
assign a5272 = ~a5270 & a4054;
assign a5274 = l586 & ~l64;
assign a5276 = ~a5274 & ~a5272;
assign a5278 = ~a5276 & ~a1744;
assign a5280 = a1744 & l580;
assign a5282 = ~a5280 & ~a5278;
assign a5284 = l584 & l340;
assign a5286 = a4120 & l588;
assign a5288 = ~a5286 & ~a5284;
assign a5290 = ~a5288 & a4054;
assign a5292 = l590 & ~l64;
assign a5294 = ~a5292 & ~a5290;
assign a5296 = ~a5294 & ~a1744;
assign a5298 = a1744 & l584;
assign a5300 = ~a5298 & ~a5296;
assign a5302 = l588 & l340;
assign a5304 = a4120 & l592;
assign a5306 = ~a5304 & ~a5302;
assign a5308 = ~a5306 & a4054;
assign a5310 = l594 & ~l64;
assign a5312 = ~a5310 & ~a5308;
assign a5314 = ~a5312 & ~a1744;
assign a5316 = a1744 & l588;
assign a5318 = ~a5316 & ~a5314;
assign a5320 = l592 & l340;
assign a5322 = a4120 & l596;
assign a5324 = ~a5322 & ~a5320;
assign a5326 = ~a5324 & a4054;
assign a5328 = l598 & ~l64;
assign a5330 = ~a5328 & ~a5326;
assign a5332 = ~a5330 & ~a1744;
assign a5334 = a1744 & l592;
assign a5336 = ~a5334 & ~a5332;
assign a5338 = a3768 & l406;
assign a5340 = a5338 & l600;
assign a5342 = l596 & l340;
assign a5344 = a4120 & l602;
assign a5346 = ~a5344 & ~a5342;
assign a5348 = ~a5346 & ~a3768;
assign a5350 = ~a5348 & ~a5340;
assign a5352 = ~a5350 & l64;
assign a5354 = l604 & ~l64;
assign a5356 = ~a5354 & ~a5352;
assign a5358 = ~a5356 & ~a1744;
assign a5360 = a1744 & l596;
assign a5362 = ~a5360 & ~a5358;
assign a5364 = a1388 & l64;
assign a5366 = ~a5364 & ~l600;
assign a5368 = a5338 & l606;
assign a5370 = l602 & l340;
assign a5372 = a4120 & l608;
assign a5374 = ~a5372 & ~a5370;
assign a5376 = ~a5374 & ~a3768;
assign a5378 = ~a5376 & ~a5368;
assign a5380 = ~a5378 & l64;
assign a5382 = l610 & ~l64;
assign a5384 = ~a5382 & ~a5380;
assign a5386 = ~a5384 & ~a1744;
assign a5388 = a1744 & l602;
assign a5390 = ~a5388 & ~a5386;
assign a5392 = a1380 & l64;
assign a5394 = ~a5392 & ~l606;
assign a5396 = a5338 & l612;
assign a5398 = l608 & l340;
assign a5400 = a4120 & l614;
assign a5402 = ~a5400 & ~a5398;
assign a5404 = ~a5402 & ~a3768;
assign a5406 = ~a5404 & ~a5396;
assign a5408 = ~a5406 & l64;
assign a5410 = l616 & ~l64;
assign a5412 = ~a5410 & ~a5408;
assign a5414 = ~a5412 & ~a1744;
assign a5416 = a1744 & l608;
assign a5418 = ~a5416 & ~a5414;
assign a5420 = a1366 & l64;
assign a5422 = ~a5420 & ~l612;
assign a5424 = a5338 & l618;
assign a5426 = l614 & l340;
assign a5428 = a4120 & l620;
assign a5430 = ~a5428 & ~a5426;
assign a5432 = ~a5430 & ~a3768;
assign a5434 = ~a5432 & ~a5424;
assign a5436 = ~a5434 & l64;
assign a5438 = l622 & ~l64;
assign a5440 = ~a5438 & ~a5436;
assign a5442 = ~a5440 & ~a1744;
assign a5444 = a1744 & l614;
assign a5446 = ~a5444 & ~a5442;
assign a5448 = a1360 & l64;
assign a5450 = ~a5448 & ~l618;
assign a5452 = a5338 & l624;
assign a5454 = l620 & l340;
assign a5456 = a4120 & l626;
assign a5458 = ~a5456 & ~a5454;
assign a5460 = ~a5458 & ~a3768;
assign a5462 = ~a5460 & ~a5452;
assign a5464 = ~a5462 & l64;
assign a5466 = l628 & ~l64;
assign a5468 = ~a5466 & ~a5464;
assign a5470 = ~a5468 & ~a1744;
assign a5472 = a1744 & l620;
assign a5474 = ~a5472 & ~a5470;
assign a5476 = l158 & l152;
assign a5478 = a5476 & a2340;
assign a5480 = ~a5478 & ~l624;
assign a5482 = a5338 & l630;
assign a5484 = l626 & l340;
assign a5486 = a4120 & l632;
assign a5488 = ~a5486 & ~a5484;
assign a5490 = ~a5488 & ~a3768;
assign a5492 = ~a5490 & ~a5482;
assign a5494 = ~a5492 & l64;
assign a5496 = l634 & ~l64;
assign a5498 = ~a5496 & ~a5494;
assign a5500 = ~a5498 & ~a1744;
assign a5502 = a1744 & l626;
assign a5504 = ~a5502 & ~a5500;
assign a5506 = a1342 & l64;
assign a5508 = ~a5506 & ~l630;
assign a5510 = a5338 & l636;
assign a5512 = l632 & l340;
assign a5514 = a4120 & l638;
assign a5516 = ~a5514 & ~a5512;
assign a5518 = ~a5516 & ~a3768;
assign a5520 = ~a5518 & ~a5510;
assign a5522 = ~a5520 & l64;
assign a5524 = l640 & ~l64;
assign a5526 = ~a5524 & ~a5522;
assign a5528 = ~a5526 & ~a1744;
assign a5530 = a1744 & l632;
assign a5532 = ~a5530 & ~a5528;
assign a5534 = a1340 & l64;
assign a5536 = ~a5534 & ~l636;
assign a5538 = a5338 & l642;
assign a5540 = l638 & l340;
assign a5542 = a4120 & l644;
assign a5544 = ~a5542 & ~a5540;
assign a5546 = ~a5544 & ~a3768;
assign a5548 = ~a5546 & ~a5538;
assign a5550 = ~a5548 & l64;
assign a5552 = l646 & ~l64;
assign a5554 = ~a5552 & ~a5550;
assign a5556 = ~a5554 & ~a1744;
assign a5558 = a1744 & l638;
assign a5560 = ~a5558 & ~a5556;
assign a5562 = a1386 & l64;
assign a5564 = ~a5562 & ~l642;
assign a5566 = a5338 & l648;
assign a5568 = l644 & l340;
assign a5570 = a4120 & l650;
assign a5572 = ~a5570 & ~a5568;
assign a5574 = ~a5572 & ~a3768;
assign a5576 = ~a5574 & ~a5566;
assign a5578 = ~a5576 & l64;
assign a5580 = l652 & ~l64;
assign a5582 = ~a5580 & ~a5578;
assign a5584 = ~a5582 & ~a1744;
assign a5586 = a1744 & l644;
assign a5588 = ~a5586 & ~a5584;
assign a5590 = a1384 & l64;
assign a5592 = ~a5590 & ~l648;
assign a5594 = a5338 & l654;
assign a5596 = l650 & l340;
assign a5598 = a4120 & l656;
assign a5600 = ~a5598 & ~a5596;
assign a5602 = ~a5600 & ~a3768;
assign a5604 = ~a5602 & ~a5594;
assign a5606 = ~a5604 & l64;
assign a5608 = l658 & ~l64;
assign a5610 = ~a5608 & ~a5606;
assign a5612 = ~a5610 & ~a1744;
assign a5614 = a1744 & l650;
assign a5616 = ~a5614 & ~a5612;
assign a5618 = a1364 & l64;
assign a5620 = ~a5618 & ~l654;
assign a5622 = a5338 & l660;
assign a5624 = l656 & l340;
assign a5626 = a4120 & l662;
assign a5628 = ~a5626 & ~a5624;
assign a5630 = ~a5628 & ~a3768;
assign a5632 = ~a5630 & ~a5622;
assign a5634 = ~a5632 & l64;
assign a5636 = l664 & ~l64;
assign a5638 = ~a5636 & ~a5634;
assign a5640 = ~a5638 & ~a1744;
assign a5642 = a1744 & l656;
assign a5644 = ~a5642 & ~a5640;
assign a5646 = a1334 & l64;
assign a5648 = ~a5646 & ~l660;
assign a5650 = a5338 & l666;
assign a5652 = l662 & l340;
assign a5654 = a4120 & l668;
assign a5656 = ~a5654 & ~a5652;
assign a5658 = ~a5656 & ~a3768;
assign a5660 = ~a5658 & ~a5650;
assign a5662 = ~a5660 & l64;
assign a5664 = l670 & ~l64;
assign a5666 = ~a5664 & ~a5662;
assign a5668 = ~a5666 & ~a1744;
assign a5670 = a1744 & l662;
assign a5672 = ~a5670 & ~a5668;
assign a5674 = a1332 & l64;
assign a5676 = ~a5674 & ~l666;
assign a5678 = a5338 & l672;
assign a5680 = l668 & l340;
assign a5682 = a4120 & l674;
assign a5684 = ~a5682 & ~a5680;
assign a5686 = ~a5684 & ~a3768;
assign a5688 = ~a5686 & ~a5678;
assign a5690 = ~a5688 & l64;
assign a5692 = l676 & ~l64;
assign a5694 = ~a5692 & ~a5690;
assign a5696 = ~a5694 & ~a1744;
assign a5698 = a1744 & l668;
assign a5700 = ~a5698 & ~a5696;
assign a5702 = a1318 & l64;
assign a5704 = ~a5702 & ~l672;
assign a5706 = a5338 & l678;
assign a5708 = l674 & l340;
assign a5710 = a4120 & l680;
assign a5712 = ~a5710 & ~a5708;
assign a5714 = ~a5712 & ~a3768;
assign a5716 = ~a5714 & ~a5706;
assign a5718 = ~a5716 & l64;
assign a5720 = l682 & ~l64;
assign a5722 = ~a5720 & ~a5718;
assign a5724 = ~a5722 & ~a1744;
assign a5726 = a1744 & l674;
assign a5728 = ~a5726 & ~a5724;
assign a5730 = a1372 & l64;
assign a5732 = ~a5730 & ~l678;
assign a5734 = l680 & l340;
assign a5736 = a4120 & l684;
assign a5738 = ~a5736 & ~a5734;
assign a5740 = ~a5738 & a4054;
assign a5742 = l686 & ~l64;
assign a5744 = ~a5742 & ~a5740;
assign a5746 = ~a5744 & ~a1744;
assign a5748 = a1744 & l680;
assign a5750 = ~a5748 & ~a5746;
assign a5752 = l684 & l340;
assign a5754 = a4120 & l688;
assign a5756 = ~a5754 & ~a5752;
assign a5758 = ~a5756 & a4054;
assign a5760 = l690 & ~l64;
assign a5762 = ~a5760 & ~a5758;
assign a5764 = ~a5762 & ~a1744;
assign a5766 = a1744 & l684;
assign a5768 = ~a5766 & ~a5764;
assign a5770 = l688 & l340;
assign a5772 = a4120 & l692;
assign a5774 = ~a5772 & ~a5770;
assign a5776 = ~a5774 & a4054;
assign a5778 = l694 & ~l64;
assign a5780 = ~a5778 & ~a5776;
assign a5782 = ~a5780 & ~a1744;
assign a5784 = a1744 & l688;
assign a5786 = ~a5784 & ~a5782;
assign a5788 = l692 & l340;
assign a5790 = a4120 & l696;
assign a5792 = ~a5790 & ~a5788;
assign a5794 = ~a5792 & a4054;
assign a5796 = l698 & ~l64;
assign a5798 = ~a5796 & ~a5794;
assign a5800 = ~a5798 & ~a1744;
assign a5802 = a1744 & l692;
assign a5804 = ~a5802 & ~a5800;
assign a5806 = l696 & l340;
assign a5808 = a4120 & l700;
assign a5810 = ~a5808 & ~a5806;
assign a5812 = ~a5810 & a4054;
assign a5814 = l702 & ~l64;
assign a5816 = ~a5814 & ~a5812;
assign a5818 = ~a5816 & ~a1744;
assign a5820 = a1744 & l696;
assign a5822 = ~a5820 & ~a5818;
assign a5824 = l700 & l340;
assign a5826 = a4120 & l704;
assign a5828 = ~a5826 & ~a5824;
assign a5830 = ~a5828 & a4054;
assign a5832 = l706 & ~l64;
assign a5834 = ~a5832 & ~a5830;
assign a5836 = ~a5834 & ~a1744;
assign a5838 = a1744 & l700;
assign a5840 = ~a5838 & ~a5836;
assign a5842 = l704 & l340;
assign a5844 = a4120 & l708;
assign a5846 = ~a5844 & ~a5842;
assign a5848 = ~a5846 & a4054;
assign a5850 = l710 & ~l64;
assign a5852 = ~a5850 & ~a5848;
assign a5854 = ~a5852 & ~a1744;
assign a5856 = a1744 & l704;
assign a5858 = ~a5856 & ~a5854;
assign a5860 = l708 & l340;
assign a5862 = a4120 & l712;
assign a5864 = ~a5862 & ~a5860;
assign a5866 = ~a5864 & a4054;
assign a5868 = l714 & ~l64;
assign a5870 = ~a5868 & ~a5866;
assign a5872 = ~a5870 & ~a1744;
assign a5874 = a1744 & l708;
assign a5876 = ~a5874 & ~a5872;
assign a5878 = l712 & l340;
assign a5880 = a4120 & l716;
assign a5882 = ~a5880 & ~a5878;
assign a5884 = ~a5882 & a4054;
assign a5886 = l718 & ~l64;
assign a5888 = ~a5886 & ~a5884;
assign a5890 = ~a5888 & ~a1744;
assign a5892 = a1744 & l712;
assign a5894 = ~a5892 & ~a5890;
assign a5896 = l716 & l340;
assign a5898 = a4120 & l720;
assign a5900 = ~a5898 & ~a5896;
assign a5902 = ~a5900 & a4054;
assign a5904 = l722 & ~l64;
assign a5906 = ~a5904 & ~a5902;
assign a5908 = ~a5906 & ~a1744;
assign a5910 = a1744 & l716;
assign a5912 = ~a5910 & ~a5908;
assign a5914 = l720 & l340;
assign a5916 = a4120 & l724;
assign a5918 = ~a5916 & ~a5914;
assign a5920 = ~a5918 & a4054;
assign a5922 = l726 & ~l64;
assign a5924 = ~a5922 & ~a5920;
assign a5926 = ~a5924 & ~a1744;
assign a5928 = a1744 & l720;
assign a5930 = ~a5928 & ~a5926;
assign a5932 = l724 & l340;
assign a5934 = a4120 & l728;
assign a5936 = ~a5934 & ~a5932;
assign a5938 = ~a5936 & a4054;
assign a5940 = l730 & ~l64;
assign a5942 = ~a5940 & ~a5938;
assign a5944 = ~a5942 & ~a1744;
assign a5946 = a1744 & l724;
assign a5948 = ~a5946 & ~a5944;
assign a5950 = l728 & l340;
assign a5952 = a4120 & l732;
assign a5954 = ~a5952 & ~a5950;
assign a5956 = ~a5954 & a4054;
assign a5958 = l734 & ~l64;
assign a5960 = ~a5958 & ~a5956;
assign a5962 = ~a5960 & ~a1744;
assign a5964 = a1744 & l728;
assign a5966 = ~a5964 & ~a5962;
assign a5968 = l732 & l340;
assign a5970 = a4120 & l736;
assign a5972 = ~a5970 & ~a5968;
assign a5974 = ~a5972 & a4054;
assign a5976 = l738 & ~l64;
assign a5978 = ~a5976 & ~a5974;
assign a5980 = ~a5978 & ~a1744;
assign a5982 = a1744 & l732;
assign a5984 = ~a5982 & ~a5980;
assign a5986 = l736 & l340;
assign a5988 = a4120 & l740;
assign a5990 = ~a5988 & ~a5986;
assign a5992 = ~a5990 & a4054;
assign a5994 = l742 & ~l64;
assign a5996 = ~a5994 & ~a5992;
assign a5998 = ~a5996 & ~a1744;
assign a6000 = a1744 & l736;
assign a6002 = ~a6000 & ~a5998;
assign a6004 = l740 & l340;
assign a6006 = a4120 & l744;
assign a6008 = ~a6006 & ~a6004;
assign a6010 = ~a6008 & a4054;
assign a6012 = l746 & ~l64;
assign a6014 = ~a6012 & ~a6010;
assign a6016 = ~a6014 & ~a1744;
assign a6018 = a1744 & l740;
assign a6020 = ~a6018 & ~a6016;
assign a6022 = l744 & l340;
assign a6024 = a4120 & l748;
assign a6026 = ~a6024 & ~a6022;
assign a6028 = ~a6026 & a4054;
assign a6030 = l750 & ~l64;
assign a6032 = ~a6030 & ~a6028;
assign a6034 = ~a6032 & ~a1744;
assign a6036 = a1744 & l744;
assign a6038 = ~a6036 & ~a6034;
assign a6040 = l748 & l340;
assign a6042 = a3722 & l752;
assign a6044 = a6042 & a4120;
assign a6046 = ~a6044 & ~a6040;
assign a6048 = ~a6046 & a4054;
assign a6050 = l754 & ~l64;
assign a6052 = ~a6050 & ~a6048;
assign a6054 = ~a6052 & ~a1744;
assign a6056 = a1744 & l748;
assign a6058 = ~a6056 & ~a6054;
assign a6060 = ~a3850 & l350;
assign a6062 = ~a6060 & ~l352;
assign a6064 = ~a6062 & l64;
assign a6066 = l756 & ~l64;
assign a6068 = ~a6066 & ~a6064;
assign a6070 = ~a6068 & ~a2156;
assign a6072 = a2156 & l752;
assign a6074 = ~a6072 & ~a6070;
assign a6076 = l62 & ~l60;
assign a6078 = ~a6076 & ~a2188;
assign a6080 = a6078 & l132;
assign a6082 = ~a6078 & ~l132;
assign a6084 = ~a6082 & ~a6080;
assign a6086 = l140 & ~l124;
assign a6088 = ~l140 & l124;
assign a6090 = ~a6088 & ~a6086;
assign a6092 = ~l450 & ~l128;
assign a6094 = l450 & l128;
assign a6096 = ~a6094 & ~a6092;
assign a6098 = a6096 & a6090;
assign a6100 = ~a6096 & ~a6090;
assign a6102 = ~a6100 & ~a6098;
assign a6104 = a6102 & a6084;
assign a6106 = ~a6102 & ~a6084;
assign a6108 = ~a6106 & ~a6104;
assign a6110 = l182 & l126;
assign a6112 = ~a6110 & ~a2190;
assign a6114 = ~a6112 & l476;
assign a6116 = a6112 & ~l476;
assign a6118 = ~a6116 & ~a6114;
assign a6120 = l470 & l158;
assign a6122 = ~a6120 & ~a1362;
assign a6124 = ~l178 & l142;
assign a6126 = l178 & ~l142;
assign a6128 = ~a6126 & ~a6124;
assign a6130 = ~a6128 & ~a6122;
assign a6132 = a6128 & a6122;
assign a6134 = ~a6132 & ~a6130;
assign a6136 = a6134 & ~a6118;
assign a6138 = ~a6134 & a6118;
assign a6140 = ~a6138 & ~a6136;
assign a6142 = ~a6140 & ~a6108;
assign a6144 = a6140 & a6108;
assign a6146 = ~l176 & l142;
assign a6148 = l140 & ~l130;
assign a6150 = ~a6148 & ~a6146;
assign a6152 = a1610 & ~l178;
assign a6154 = a6092 & a1772;
assign a6156 = a6154 & a6152;
assign a6158 = ~a6156 & l84;
assign a6160 = ~a6158 & a6150;
assign a6162 = a6160 & ~a6144;
assign a6164 = a6162 & ~a6142;
assign a6166 = ~a6164 & l64;
assign a6168 = l758 & ~l64;
assign a6170 = ~a6168 & ~a6166;
assign a6172 = a4360 & ~l450;
assign a6174 = l792 & l450;
assign a6176 = ~a6174 & l760;
assign a6178 = a6174 & l770;
assign a6180 = ~a6178 & ~a6176;
assign a6182 = a6180 & ~a6172;
assign a6184 = ~a6182 & l64;
assign a6186 = l846 & ~l64;
assign a6188 = ~a6186 & ~a6184;
assign a6190 = ~a6188 & ~a1410;
assign a6192 = a1410 & l760;
assign a6194 = ~a6192 & ~a6190;
assign a6196 = ~a6174 & l762;
assign a6198 = a6174 & l764;
assign a6200 = ~a6198 & ~a6196;
assign a6202 = a6200 & ~a6172;
assign a6204 = ~a6202 & l64;
assign a6206 = l844 & ~l64;
assign a6208 = ~a6206 & ~a6204;
assign a6210 = ~a6208 & ~a1410;
assign a6212 = a1410 & l762;
assign a6214 = ~a6212 & ~a6210;
assign a6216 = a6174 & l760;
assign a6218 = a6216 & l764;
assign a6220 = ~a6216 & ~l764;
assign a6222 = ~a6220 & ~a6218;
assign a6224 = ~a6222 & ~a6172;
assign a6226 = ~a6224 & l64;
assign a6228 = l842 & ~l64;
assign a6230 = ~a6228 & ~a6226;
assign a6232 = ~a6230 & ~a1410;
assign a6234 = a1410 & l764;
assign a6236 = ~a6234 & ~a6232;
assign a6238 = ~a6174 & l766;
assign a6240 = a6174 & l768;
assign a6242 = ~a6240 & ~a6238;
assign a6244 = a6242 & ~a6172;
assign a6246 = ~a6244 & l64;
assign a6248 = l840 & ~l64;
assign a6250 = ~a6248 & ~a6246;
assign a6252 = ~a6250 & ~a1410;
assign a6254 = a1410 & l766;
assign a6256 = ~a6254 & ~a6252;
assign a6258 = ~a6174 & l768;
assign a6260 = a6174 & l762;
assign a6262 = ~a6260 & ~a6258;
assign a6264 = a6262 & ~a6172;
assign a6266 = ~a6264 & l64;
assign a6268 = l838 & ~l64;
assign a6270 = ~a6268 & ~a6266;
assign a6272 = ~a6270 & ~a1410;
assign a6274 = a1410 & l768;
assign a6276 = ~a6274 & ~a6272;
assign a6278 = ~a6174 & l770;
assign a6280 = a6174 & l772;
assign a6282 = ~a6280 & ~a6278;
assign a6284 = a6282 & ~a6172;
assign a6286 = ~a6284 & l64;
assign a6288 = l836 & ~l64;
assign a6290 = ~a6288 & ~a6286;
assign a6292 = ~a6290 & ~a1410;
assign a6294 = a1410 & l770;
assign a6296 = ~a6294 & ~a6292;
assign a6298 = ~a6174 & l772;
assign a6300 = a6174 & l766;
assign a6302 = ~a6300 & ~a6298;
assign a6304 = a6302 & ~a6172;
assign a6306 = ~a6304 & l64;
assign a6308 = l794 & ~l64;
assign a6310 = ~a6308 & ~a6306;
assign a6312 = ~a6310 & ~a1410;
assign a6314 = a1410 & l772;
assign a6316 = ~a6314 & ~a6312;
assign a6318 = a1692 & ~l124;
assign a6320 = ~l806 & ~l804;
assign a6322 = a6320 & ~l802;
assign a6324 = ~a6322 & l450;
assign a6326 = ~a6324 & ~a6172;
assign a6328 = a6326 & ~a6318;
assign a6330 = ~l450 & ~l124;
assign a6332 = a6330 & l774;
assign a6334 = ~a6330 & l776;
assign a6336 = ~a6334 & ~a6332;
assign a6338 = a6336 & a6328;
assign a6340 = ~a6338 & l64;
assign a6342 = l834 & ~l64;
assign a6344 = ~a6342 & ~a6340;
assign a6346 = ~a6344 & ~a1410;
assign a6348 = a1410 & l774;
assign a6350 = ~a6348 & ~a6346;
assign a6352 = a6330 & l776;
assign a6354 = ~a6330 & l778;
assign a6356 = ~a6354 & ~a6352;
assign a6358 = a6356 & a6328;
assign a6360 = ~a6358 & l64;
assign a6362 = l832 & ~l64;
assign a6364 = ~a6362 & ~a6360;
assign a6366 = ~a6364 & ~a1410;
assign a6368 = a1410 & l776;
assign a6370 = ~a6368 & ~a6366;
assign a6372 = a6330 & l778;
assign a6374 = ~a6330 & l780;
assign a6376 = ~a6374 & ~a6372;
assign a6378 = a6376 & a6328;
assign a6380 = ~a6378 & l64;
assign a6382 = l830 & ~l64;
assign a6384 = ~a6382 & ~a6380;
assign a6386 = ~a6384 & ~a1410;
assign a6388 = a1410 & l778;
assign a6390 = ~a6388 & ~a6386;
assign a6392 = a6330 & l780;
assign a6394 = ~a6330 & l786;
assign a6396 = ~a6394 & ~a6392;
assign a6398 = a6396 & a6328;
assign a6400 = ~a6398 & l64;
assign a6402 = l828 & ~l64;
assign a6404 = ~a6402 & ~a6400;
assign a6406 = ~a6404 & ~a1410;
assign a6408 = a1410 & l780;
assign a6410 = ~a6408 & ~a6406;
assign a6412 = a6330 & l782;
assign a6414 = ~a6330 & l788;
assign a6416 = ~a6414 & ~a6412;
assign a6418 = a6416 & a6328;
assign a6420 = ~a6418 & l64;
assign a6422 = l826 & ~l64;
assign a6424 = ~a6422 & ~a6420;
assign a6426 = ~a6424 & ~a1410;
assign a6428 = a1410 & l782;
assign a6430 = ~a6428 & ~a6426;
assign a6432 = a6330 & l784;
assign a6434 = ~a6330 & l790;
assign a6436 = ~a6434 & ~a6432;
assign a6438 = a6436 & a6328;
assign a6440 = ~a6438 & l64;
assign a6442 = l824 & ~l64;
assign a6444 = ~a6442 & ~a6440;
assign a6446 = ~a6444 & ~a1410;
assign a6448 = a1410 & l784;
assign a6450 = ~a6448 & ~a6446;
assign a6452 = a6330 & l786;
assign a6454 = ~a6330 & l782;
assign a6456 = ~a6454 & ~a6452;
assign a6458 = a6456 & a6328;
assign a6460 = ~a6458 & l64;
assign a6462 = l822 & ~l64;
assign a6464 = ~a6462 & ~a6460;
assign a6466 = ~a6464 & ~a1410;
assign a6468 = a1410 & l786;
assign a6470 = ~a6468 & ~a6466;
assign a6472 = a6330 & l788;
assign a6474 = ~a6330 & l784;
assign a6476 = ~a6474 & ~a6472;
assign a6478 = a6476 & a6328;
assign a6480 = ~a6478 & l64;
assign a6482 = l820 & ~l64;
assign a6484 = ~a6482 & ~a6480;
assign a6486 = ~a6484 & ~a1410;
assign a6488 = a1410 & l788;
assign a6490 = ~a6488 & ~a6486;
assign a6492 = a6330 & l790;
assign a6494 = l782 & ~l774;
assign a6496 = ~l782 & l774;
assign a6498 = ~a6496 & ~a6494;
assign a6500 = ~a6498 & ~a6330;
assign a6502 = ~a6500 & ~a6492;
assign a6504 = a6502 & a6328;
assign a6506 = ~a6504 & l64;
assign a6508 = l808 & ~l64;
assign a6510 = ~a6508 & ~a6506;
assign a6512 = ~a6510 & ~a1410;
assign a6514 = a2032 & a1408;
assign a6516 = ~a6514 & ~a6512;
assign a6518 = l798 & l64;
assign a6520 = a6518 & ~l796;
assign a6522 = l792 & ~l64;
assign a6524 = ~a6522 & ~a6520;
assign a6526 = l796 & ~l64;
assign a6528 = ~a6526 & ~a6518;
assign a6530 = l64 & i12;
assign a6532 = l800 & ~l64;
assign a6534 = ~a6532 & ~a6530;
assign a6536 = ~a6534 & ~a2156;
assign a6538 = a2156 & l798;
assign a6540 = ~a6538 & ~a6536;
assign a6542 = l810 & l64;
assign a6544 = l64 & i18;
assign a6546 = l818 & ~l64;
assign a6548 = ~a6546 & ~a6544;
assign a6550 = ~a6548 & ~a6542;
assign a6552 = a6542 & l802;
assign a6554 = ~a6552 & ~a6550;
assign a6556 = l64 & i16;
assign a6558 = l816 & ~l64;
assign a6560 = ~a6558 & ~a6556;
assign a6562 = ~a6560 & ~a6542;
assign a6564 = a6542 & l804;
assign a6566 = ~a6564 & ~a6562;
assign a6568 = l64 & i14;
assign a6570 = l812 & ~l64;
assign a6572 = ~a6570 & ~a6568;
assign a6574 = ~a6572 & ~a6542;
assign a6576 = a6542 & l806;
assign a6578 = ~a6576 & ~a6574;
assign a6580 = ~a1692 & l124;
assign a6582 = ~a1606 & l64;
assign a6584 = a6582 & ~a1640;
assign a6586 = a6584 & ~a2028;
assign a6588 = a6586 & ~a1702;
assign a6590 = a6588 & ~a1592;
assign a6592 = a6590 & ~a1426;
assign a6594 = a6592 & ~a6580;
assign a6596 = a6594 & l850;
assign a6598 = l854 & ~l64;
assign a6600 = ~a6598 & ~a6596;
assign a6602 = ~a6600 & ~a1410;
assign a6604 = a1410 & l848;
assign a6606 = ~a6604 & ~a6602;
assign a6608 = l858 & l792;
assign a6610 = a6608 & l856;
assign a6612 = ~a6610 & ~l850;
assign a6614 = ~a6612 & ~l66;
assign a6616 = a6614 & a6594;
assign a6618 = l860 & ~l64;
assign a6620 = ~a6618 & ~a6616;
assign a6622 = ~a6620 & ~a1410;
assign a6624 = a1410 & l850;
assign a6626 = ~a6624 & ~a6622;
assign a6628 = l64 & i20;
assign a6630 = l852 & ~l64;
assign a6632 = ~a6630 & ~a6628;
assign a6634 = ~a6608 & ~l856;
assign a6636 = ~a6634 & a6594;
assign a6638 = l864 & ~l64;
assign a6640 = ~a6638 & ~a6636;
assign a6642 = ~a6640 & ~a1410;
assign a6644 = a1410 & l856;
assign a6646 = ~a6644 & ~a6642;
assign a6648 = a1362 & ~l132;
assign a6650 = ~l476 & ~l124;
assign a6652 = a6650 & a1576;
assign a6654 = a6652 & a6648;
assign a6656 = ~a6654 & a6594;
assign a6658 = l862 & ~l64;
assign a6660 = ~a6658 & ~a6656;
assign a6662 = ~a6660 & ~a1410;
assign a6664 = a1410 & l858;
assign a6666 = ~a6664 & ~a6662;
assign a6668 = l64 & i22;
assign a6670 = l868 & ~l64;
assign a6672 = ~a6670 & ~a6668;
assign a6674 = ~a6672 & ~a2156;
assign a6676 = a2156 & l866;
assign a6678 = ~a6676 & ~a6674;
assign a6680 = l64 & i24;
assign a6682 = l870 & ~l64;
assign a6684 = ~a6682 & ~a6680;
assign a6686 = ~l876 & l872;
assign a6688 = a6686 & ~l198;
assign a6690 = ~a6688 & ~a3084;
assign a6692 = ~a6690 & l64;
assign a6694 = l878 & ~l64;
assign a6696 = ~a6694 & ~a6692;
assign a6698 = ~a6696 & ~a2156;
assign a6700 = a2156 & l872;
assign a6702 = ~a6700 & ~a6698;
assign a6704 = ~l880 & ~l64;
assign a6706 = a2156 & ~l876;
assign a6710 = ~l916 & ~l350;
assign a6712 = ~a6710 & a2472;
assign a6714 = a6712 & ~a4174;
assign a6716 = l924 & ~l64;
assign a6718 = ~a6716 & ~a6714;
assign a6720 = ~a6718 & ~a2156;
assign a6722 = a2156 & l916;
assign a6724 = ~a6722 & ~a6720;
assign a6726 = ~l482 & ~l472;
assign a6728 = ~l650 & ~l638;
assign a6730 = a6728 & a6726;
assign a6732 = ~l478 & ~l466;
assign a6734 = ~l500 & ~l488;
assign a6736 = a6734 & a6732;
assign a6738 = a6736 & a6730;
assign a6740 = ~l462 & ~l452;
assign a6742 = ~l674 & ~l662;
assign a6744 = a6742 & a6740;
assign a6746 = ~l692 & ~l684;
assign a6748 = ~l708 & ~l700;
assign a6750 = a6748 & a6746;
assign a6752 = a6750 & a6744;
assign a6754 = a6752 & a6738;
assign a6756 = ~l632 & ~l620;
assign a6758 = ~l528 & ~l514;
assign a6760 = a6758 & a6756;
assign a6762 = ~l608 & ~l596;
assign a6764 = ~l550 & ~l540;
assign a6766 = a6764 & a6762;
assign a6768 = a6766 & a6760;
assign a6770 = ~l438 & ~l432;
assign a6772 = ~l740 & ~l732;
assign a6774 = a6772 & a6770;
assign a6776 = ~l458 & ~l444;
assign a6778 = ~l752 & ~l748;
assign a6780 = a6778 & a6776;
assign a6782 = a6780 & a6774;
assign a6784 = a6782 & a6768;
assign a6786 = a6784 & a6754;
assign a6788 = ~l744 & ~l736;
assign a6790 = ~l696 & ~l688;
assign a6792 = a6790 & a6788;
assign a6794 = ~l728 & ~l720;
assign a6796 = ~l680 & ~l668;
assign a6798 = a6796 & a6794;
assign a6800 = a6798 & a6792;
assign a6802 = ~l534 & ~l522;
assign a6804 = ~l568 & ~l560;
assign a6806 = a6804 & a6802;
assign a6808 = ~l506 & ~l494;
assign a6810 = ~l584 & ~l576;
assign a6812 = a6810 & a6808;
assign a6814 = a6812 & a6806;
assign a6816 = a6814 & a6800;
assign a6818 = ~l602 & ~l592;
assign a6820 = ~l626 & ~l614;
assign a6822 = a6820 & a6818;
assign a6824 = ~l588 & ~l580;
assign a6826 = ~l572 & ~l564;
assign a6828 = a6826 & a6824;
assign a6830 = a6828 & a6822;
assign a6832 = ~l424 & ~l352;
assign a6834 = ~l346 & l64;
assign a6836 = a6834 & ~l410;
assign a6838 = a6836 & a6832;
assign a6840 = ~l656 & ~l644;
assign a6842 = ~l724 & ~l716;
assign a6844 = a6842 & a6840;
assign a6846 = ~l712 & ~l704;
assign a6848 = ~l554 & ~l546;
assign a6850 = a6848 & a6846;
assign a6852 = a6850 & a6844;
assign a6854 = a6852 & a6838;
assign a6856 = a6854 & a6830;
assign a6858 = a6856 & a6816;
assign a6860 = a6858 & a6786;
assign a6862 = l922 & ~l64;
assign a6864 = ~a6862 & ~a6860;
assign a6866 = ~a6864 & ~a2156;
assign a6868 = a2156 & l918;
assign a6870 = ~a6868 & ~a6866;
assign a6872 = a3300 & a3236;
assign a6874 = a3172 & l928;
assign a6876 = ~a6874 & ~a6872;
assign a6878 = ~a6876 & l64;
assign a6880 = l948 & ~l64;
assign a6882 = ~a6880 & ~a6878;
assign a6884 = ~a6882 & ~a1744;
assign a6886 = a1744 & l928;
assign a6888 = ~a6886 & ~a6884;
assign a6890 = a3212 & l220;
assign a6892 = a6890 & a3236;
assign a6894 = a3172 & l930;
assign a6896 = ~a6894 & ~a6892;
assign a6898 = ~a6896 & l64;
assign a6900 = l946 & ~l64;
assign a6902 = ~a6900 & ~a6898;
assign a6904 = ~a6902 & ~a1744;
assign a6906 = a1744 & l930;
assign a6908 = ~a6906 & ~a6904;
assign a6910 = a3164 & l218;
assign a6912 = a3172 & l932;
assign a6914 = ~a6912 & ~a6910;
assign a6916 = ~a6914 & l64;
assign a6918 = l944 & ~l64;
assign a6920 = ~a6918 & ~a6916;
assign a6922 = ~a6920 & ~a1744;
assign a6924 = a1744 & l932;
assign a6926 = ~a6924 & ~a6922;
assign a6928 = a3190 & l218;
assign a6930 = a3172 & l934;
assign a6932 = ~a6930 & ~a6928;
assign a6934 = ~a6932 & l64;
assign a6936 = l942 & ~l64;
assign a6938 = ~a6936 & ~a6934;
assign a6940 = ~a6938 & ~a1744;
assign a6942 = a1744 & l934;
assign a6944 = ~a6942 & ~a6940;
assign a6946 = l214 & ~i30;
assign a6948 = l226 & ~i32;
assign a6950 = ~a6948 & ~a6946;
assign a6952 = l246 & ~i26;
assign a6954 = l250 & ~i28;
assign a6956 = ~a6954 & ~a6952;
assign a6958 = a6956 & a6950;
assign a6960 = a6958 & a3710;
assign a6962 = l940 & ~l64;
assign a6964 = ~a6962 & ~a6960;
assign a6966 = ~a6964 & ~a1744;
assign a6968 = a1744 & l936;
assign a6970 = ~a6968 & ~a6966;
assign a6972 = ~a1214 & l64;
assign a6974 = l1074 & l174;
assign a6976 = ~l1074 & ~l174;
assign a6978 = ~a6976 & ~a6974;
assign a6980 = a6978 & a6972;
assign a6982 = l1086 & ~l64;
assign a6984 = ~a6982 & ~a6980;
assign a6986 = ~a6984 & ~a1410;
assign a6988 = a1410 & l1074;
assign a6990 = ~a6988 & ~a6986;
assign a6992 = a6974 & l1076;
assign a6994 = ~a6974 & ~l1076;
assign a6996 = ~a6994 & ~a6992;
assign a6998 = a6996 & a6972;
assign a7000 = l1084 & ~l64;
assign a7002 = ~a7000 & ~a6998;
assign a7004 = ~a7002 & ~a1410;
assign a7006 = a1410 & l1076;
assign a7008 = ~a7006 & ~a7004;
assign a7010 = a6992 & l1078;
assign a7012 = ~a6992 & ~l1078;
assign a7014 = ~a7012 & ~a7010;
assign a7016 = a7014 & a6972;
assign a7018 = l1082 & ~l64;
assign a7020 = ~a7018 & ~a7016;
assign a7022 = ~a7020 & ~a1410;
assign a7024 = a1410 & l1078;
assign a7026 = ~a7024 & ~a7022;
assign a7028 = l64 & i40;
assign a7030 = l1096 & ~l64;
assign a7032 = ~a7030 & ~a7028;
assign a7034 = ~l1110 & l1108;
assign a7036 = ~a7034 & ~i46;
assign a7038 = a1430 & ~a1242;
assign a7040 = ~a7038 & ~l1112;
assign a7042 = ~a7040 & l64;
assign a7044 = l1114 & ~l64;
assign a7046 = ~a7044 & ~a7042;
assign a7048 = ~a7046 & ~a1410;
assign a7050 = a1410 & l1110;
assign a7052 = ~a7050 & ~a7048;
assign a7054 = a2130 & l444;
assign a7056 = l1112 & ~l64;
assign a7058 = ~a7056 & ~a7054;
assign a7060 = l1116 & l64;
assign a7062 = ~l1120 & ~l64;
assign a7066 = a7064 & ~a2156;
assign a7068 = a2156 & l1116;
assign a7070 = ~a7068 & ~a7066;
assign a7072 = l1118 & ~l64;
assign a7074 = ~a7072 & ~a7060;
assign a7076 = l1142 & l64;
assign a7078 = l1152 & ~l64;
assign a7080 = ~a7078 & ~a7076;
assign a7082 = ~a7080 & ~a2156;
assign a7084 = a2156 & l1138;
assign a7086 = ~a7084 & ~a7082;
assign a7088 = ~a1242 & l64;
assign a7090 = a6318 & ~l84;
assign a7092 = ~a1420 & l1140;
assign a7094 = ~a7092 & ~a7090;
assign a7096 = ~a7094 & a7088;
assign a7098 = l1150 & ~l64;
assign a7100 = ~a7098 & ~a7096;
assign a7102 = ~a7100 & ~a1410;
assign a7104 = a1410 & l1140;
assign a7106 = ~a7104 & ~a7102;
assign a7108 = l64 & i56;
assign a7110 = l1148 & ~l64;
assign a7112 = ~a7110 & ~a7108;
assign a7114 = ~a7112 & ~a2156;
assign a7116 = a2156 & l1142;
assign a7118 = ~a7116 & ~a7114;
assign a7120 = ~a1692 & a1656;
assign a7122 = ~a7120 & l1144;
assign a7124 = a1694 & l86;
assign a7126 = ~a7124 & ~a7090;
assign a7128 = a7126 & ~a7122;
assign a7130 = ~a7128 & a7088;
assign a7132 = l1146 & ~l64;
assign a7134 = ~a7132 & ~a7130;
assign a7136 = ~a7134 & ~a1410;
assign a7138 = a1410 & l1144;
assign a7140 = ~a7138 & ~a7136;
assign p0 = a6076;

assert property (~p0);

endmodule
