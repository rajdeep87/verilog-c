module m6s12 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120;

output p0;

wire na1780,a3436,a3566,a3590,na4050,na4058,na4066,na4074,na4082,na4090,na4098,na4106,na4114,na4122,a4124,
a4126,a4128,a4130,a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4402,a4446,a4448,a4450,a4452,
a4454,a4516,a4570,a4572,a4586,na4686,a4698,ni104,na4708,na4718,na4726,na4732,na4738,na4744,na4750,
na4756,na4762,na4768,na4774,ni108,ni116,a238,a240,a242,a244,a246,a248,a250,a252,a254,
a256,a258,a260,a262,a264,a266,a268,a270,a272,a274,a276,a278,a280,a282,a284,
a286,a288,a290,a292,a294,a296,a298,a300,a302,a304,a306,a308,a310,a312,a314,
a316,a318,a320,a322,a324,a326,a328,a330,a332,a334,a336,a338,a340,a342,a344,
a346,a348,a350,a352,a354,a356,a358,a360,a362,a364,a366,a368,a370,a372,a374,
a376,a378,a380,a382,a384,a386,a388,a390,a392,a394,a396,a398,a400,a402,a404,
a406,a408,a410,a412,a414,a416,a418,a420,a422,a424,a426,a428,a430,a432,a434,
a436,a438,a440,a442,a444,a446,a448,a450,a452,a454,a456,a458,a460,a462,a464,
a466,a468,a470,a472,a474,a476,a478,a480,a482,a484,a486,a488,a490,a492,a494,
a496,a498,a500,a502,a504,a506,a508,a510,a512,a514,a516,a518,a520,a522,a524,
a526,a528,a530,a532,a534,a536,a538,a540,a542,a544,a546,a548,a550,a552,a554,
a556,a558,a560,a562,a564,a566,a568,a570,a572,a574,a576,a578,a580,a582,a584,
a586,a588,a590,a592,a594,a596,a598,a600,a602,a604,a606,a608,a610,a612,a614,
a616,a618,a620,a622,a624,a626,a628,a630,a632,a634,a636,a638,a640,a642,a644,
a646,a648,a650,a652,a654,a656,a658,a660,a662,a664,a666,a668,a670,a672,a674,
a676,a678,a680,a682,a684,a686,a688,a690,a692,a694,a696,a698,a700,a702,a704,
a706,a708,a710,a712,a714,a716,a718,a720,a722,a724,a726,a728,a730,a732,a734,
a736,a738,a740,a742,a744,a746,a748,a750,a752,a754,a756,a758,a760,a762,a764,
a766,a768,a770,a772,a774,a776,a778,a780,a782,a784,a786,a788,a790,a792,a794,
a796,a798,a800,a802,a804,a806,a808,a810,a812,a814,a816,a818,a820,a822,a824,
a826,a828,a830,a832,a834,a836,a838,a840,a842,a844,a846,a848,a850,a852,a854,
a856,a858,a860,a862,a864,a866,a868,a870,a872,a874,a876,a878,a880,a882,a884,
a886,a888,a890,a892,a894,a896,a898,a900,a902,a904,a906,a908,a910,a912,a914,
a916,a918,a920,a922,a924,a926,a928,a930,a932,a934,a936,a938,a940,a942,a944,
a946,a948,a950,a952,a954,a956,a958,a960,a962,a964,a966,a968,a970,a972,a974,
a976,a978,a980,a982,a984,a986,a988,a990,a992,a994,a996,a998,a1000,a1002,a1004,
a1006,a1008,a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,a1034,
a1036,a1038,a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,a1062,a1064,
a1066,a1068,a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,a1092,a1094,
a1096,a1098,a1100,a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,a1124,
a1126,a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,a1154,
a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,a1178,a1180,a1182,a1184,
a1186,a1188,a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,a1208,a1210,a1212,a1214,
a1216,a1218,a1220,a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1242,a1244,
a1246,a1248,a1250,a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,a1268,a1270,a1272,a1274,
a1276,a1278,a1280,a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,
a1306,a1308,a1310,a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,a1334,
a1336,a1338,a1340,a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,
a1366,a1368,a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,a1388,a1390,a1392,a1394,
a1396,a1398,a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1424,
a1426,a1428,a1430,a1432,a1434,a1436,a1438,a1440,a1442,a1444,a1446,a1448,a1450,a1452,a1454,
a1456,a1458,a1460,a1462,a1464,a1466,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1482,a1484,
a1486,a1488,a1490,a1492,a1494,a1496,a1498,a1500,a1502,a1504,a1506,a1508,a1510,a1512,a1514,
a1516,a1518,a1520,a1522,a1524,a1526,a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,
a1546,a1548,a1550,a1552,a1554,a1556,a1558,a1560,a1562,a1564,a1566,a1568,a1570,a1572,a1574,
a1576,a1578,a1580,a1582,a1584,a1586,a1588,a1590,a1592,a1594,a1596,a1598,a1600,a1602,a1604,
a1606,a1608,a1610,a1612,a1614,a1616,a1618,a1620,a1622,a1624,a1626,a1628,a1630,a1632,a1634,
a1636,a1638,a1640,a1642,a1644,a1646,a1648,a1650,a1652,a1654,a1656,a1658,a1660,a1662,a1664,
a1666,a1668,a1670,a1672,a1674,a1676,a1678,a1680,a1682,a1684,a1686,a1688,a1690,a1692,a1694,
a1696,a1698,a1700,a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,
a1726,a1728,a1730,a1732,a1734,a1736,a1738,a1740,a1742,a1744,a1746,a1748,a1750,a1752,a1754,
a1756,a1758,a1760,a1762,a1764,a1766,a1768,a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,
a1786,a1788,a1790,a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,
a1816,a1818,a1820,a1822,a1824,a1826,a1828,a1830,a1832,a1834,a1836,a1838,a1840,a1842,a1844,
a1846,a1848,a1850,a1852,a1854,a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,
a1876,a1878,a1880,a1882,a1884,a1886,a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,
a1906,a1908,a1910,a1912,a1914,a1916,a1918,a1920,a1922,a1924,a1926,a1928,a1930,a1932,a1934,
a1936,a1938,a1940,a1942,a1944,a1946,a1948,a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,
a1966,a1968,a1970,a1972,a1974,a1976,a1978,a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,
a1996,a1998,a2000,a2002,a2004,a2006,a2008,a2010,a2012,a2014,a2016,a2018,a2020,a2022,a2024,
a2026,a2028,a2030,a2032,a2034,a2036,a2038,a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,
a2056,a2058,a2060,a2062,a2064,a2066,a2068,a2070,a2072,a2074,a2076,a2078,a2080,a2082,a2084,
a2086,a2088,a2090,a2092,a2094,a2096,a2098,a2100,a2102,a2104,a2106,a2108,a2110,a2112,a2114,
a2116,a2118,a2120,a2122,a2124,a2126,a2128,a2130,a2132,a2134,a2136,a2138,a2140,a2142,a2144,
a2146,a2148,a2150,a2152,a2154,a2156,a2158,a2160,a2162,a2164,a2166,a2168,a2170,a2172,a2174,
a2176,a2178,a2180,a2182,a2184,a2186,a2188,a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,
a2206,a2208,a2210,a2212,a2214,a2216,a2218,a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,
a2236,a2238,a2240,a2242,a2244,a2246,a2248,a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,
a2266,a2268,a2270,a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,
a2296,a2298,a2300,a2302,a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,
a2326,a2328,a2330,a2332,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,
a2356,a2358,a2360,a2362,a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,
a2386,a2388,a2390,a2392,a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,
a2416,a2418,a2420,a2422,a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,
a2446,a2448,a2450,a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,
a2476,a2478,a2480,a2482,a2484,a2486,a2488,a2490,a2492,a2494,a2496,a2498,a2500,a2502,a2504,
a2506,a2508,a2510,a2512,a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,
a2536,a2538,a2540,a2542,a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,
a2566,a2568,a2570,a2572,a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,
a2596,a2598,a2600,a2602,a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,
a2626,a2628,a2630,a2632,a2634,a2636,a2638,a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,
a2656,a2658,a2660,a2662,a2664,a2666,a2668,a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,
a2686,a2688,a2690,a2692,a2694,a2696,a2698,a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,
a2716,a2718,a2720,a2722,a2724,a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,
a2746,a2748,a2750,a2752,a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,
a2776,a2778,a2780,a2782,a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,
a2806,a2808,a2810,a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,
a2836,a2838,a2840,a2842,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,
a2866,a2868,a2870,a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,
a2896,a2898,a2900,a2902,a2904,a2906,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,
a2926,a2928,a2930,a2932,a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,
a2956,a2958,a2960,a2962,a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,
a2986,a2988,a2990,a2992,a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,
a3016,a3018,a3020,a3022,a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,
a3046,a3048,a3050,a3052,a3054,a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,
a3076,a3078,a3080,a3082,a3084,a3086,a3088,a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,
a3106,a3108,a3110,a3112,a3114,a3116,a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,
a3136,a3138,a3140,a3142,a3144,a3146,a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,
a3166,a3168,a3170,a3172,a3174,a3176,a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,
a3196,a3198,a3200,a3202,a3204,a3206,a3208,a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,
a3226,a3228,a3230,a3232,a3234,a3236,a3238,a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,
a3256,a3258,a3260,a3262,a3264,a3266,a3268,a3270,a3272,a3274,a3276,a3278,a3280,a3282,a3284,
a3286,a3288,a3290,a3292,a3294,a3296,a3298,a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,
a3316,a3318,a3320,a3322,a3324,a3326,a3328,a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,
a3346,a3348,a3350,a3352,a3354,a3356,a3358,a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,
a3376,a3378,a3380,a3382,a3384,a3386,a3388,a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,
a3406,a3408,a3410,a3412,a3414,a3416,a3418,a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3434,
a3438,a3440,a3442,a3444,a3446,a3448,a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,
a3468,a3470,a3472,a3474,a3476,a3478,a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,
a3498,a3500,a3502,a3504,a3506,a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,
a3528,a3530,a3532,a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,
a3558,a3560,a3562,a3564,a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,a3588,
a3592,a3594,a3596,a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,a3618,a3620,
a3622,a3624,a3626,a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3648,a3650,
a3652,a3654,a3656,a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,a3678,a3680,
a3682,a3684,a3686,a3688,a3690,a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,
a3712,a3714,a3716,a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,a3738,a3740,
a3742,a3744,a3746,a3748,a3750,a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,a3768,a3770,
a3772,a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,a3798,a3800,
a3802,a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,a3828,a3830,
a3832,a3834,a3836,a3838,a3840,a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,a3858,a3860,
a3862,a3864,a3866,a3868,a3870,a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,a3888,a3890,
a3892,a3894,a3896,a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,a3918,a3920,
a3922,a3924,a3926,a3928,a3930,a3932,a3934,a3936,a3938,a3940,a3942,a3944,a3946,a3948,a3950,
a3952,a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,a3978,a3980,
a3982,a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,a4008,a4010,
a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,a4038,a4040,
a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,a4068,a4070,
a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,a4096,a4098,a4100,
a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4146,a4148,a4150,a4152,
a4154,a4156,a4158,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,
a4184,a4186,a4188,a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,
a4214,a4216,a4218,a4220,a4222,a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,
a4244,a4246,a4248,a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,
a4274,a4276,a4278,a4280,a4282,a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,
a4304,a4306,a4308,a4310,a4312,a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,
a4334,a4336,a4338,a4340,a4342,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,
a4364,a4366,a4368,a4370,a4372,a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,
a4394,a4396,a4398,a4400,a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,
a4426,a4428,a4430,a4432,a4434,a4436,a4438,a4440,a4442,a4444,a4456,a4458,a4460,a4462,a4464,
a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4482,a4484,a4486,a4488,a4490,a4492,a4494,
a4496,a4498,a4500,a4502,a4504,a4506,a4508,a4510,a4512,a4514,a4518,a4520,a4522,a4524,a4526,
a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,a4554,a4556,
a4558,a4560,a4562,a4564,a4566,a4568,a4574,a4576,a4578,a4580,a4582,a4584,a4588,a4590,a4592,
a4594,a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,a4612,a4614,a4616,a4618,a4620,a4622,
a4624,a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,a4642,a4644,a4646,a4648,a4650,a4652,
a4654,a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,a4672,a4674,a4676,a4678,a4680,a4682,
a4684,a4686,a4688,a4690,a4692,a4694,a4696,a4700,a4702,a4704,a4706,a4708,a4710,a4712,a4714,
a4716,a4718,a4720,a4722,a4724,a4726,a4728,a4730,a4732,a4734,a4736,a4738,a4740,a4742,a4744,
a4746,a4748,a4750,a4752,a4754,a4756,a4758,a4760,a4762,a4764,a4766,a4768,a4770,a4772,a4774,
a4776,a4778,a4780,p0;

reg l122,l124,l126,l128,l130,l132,l134,l136,l138,l140,l142,l144,l146,l148,l150,
l152,l154,l156,l158,l160,l162,l164,l166,l168,l170,l172,l174,l176,l178,l180,
l182,l184,l186,l188,l190,l192,l194,l196,l198,l200,l202,l204,l206,l208,l210,
l212,l214,l216,l218,l220,l222,l224,l226,l228,l230,l232,l234,l236;

initial
begin
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
end

always @(posedge na1780)
   l122 <= na1780;

always @(posedge a3436)
   l124 <= a3436;

always @(posedge l236)
   l126 <= l236;

always @(posedge i114)
   l128 <= i114;

always @(posedge i112)
   l130 <= i112;

always @(posedge i110)
   l132 <= i110;

always @(posedge a3566)
   l134 <= a3566;

always @(posedge a3590)
   l136 <= a3590;

always @(posedge na4050)
   l138 <= na4050;

always @(posedge na4058)
   l140 <= na4058;

always @(posedge na4066)
   l142 <= na4066;

always @(posedge na4074)
   l144 <= na4074;

always @(posedge na4082)
   l146 <= na4082;

always @(posedge na4090)
   l148 <= na4090;

always @(posedge na4098)
   l150 <= na4098;

always @(posedge na4106)
   l152 <= na4106;

always @(posedge na4114)
   l154 <= na4114;

always @(posedge na4122)
   l156 <= na4122;

always @(posedge a4124)
   l158 <= a4124;

always @(posedge a4126)
   l160 <= a4126;

always @(posedge a4128)
   l162 <= a4128;

always @(posedge a4130)
   l164 <= a4130;

always @(posedge a4132)
   l166 <= a4132;

always @(posedge a4134)
   l168 <= a4134;

always @(posedge a4136)
   l170 <= a4136;

always @(posedge a4138)
   l172 <= a4138;

always @(posedge a4140)
   l174 <= a4140;

always @(posedge a4142)
   l176 <= a4142;

always @(posedge a4144)
   l178 <= a4144;

always @(posedge a4402)
   l180 <= a4402;

always @(posedge a4446)
   l182 <= a4446;

always @(posedge a4448)
   l184 <= a4448;

always @(posedge a4450)
   l186 <= a4450;

always @(posedge a4452)
   l188 <= a4452;

always @(posedge i82)
   l190 <= i82;

always @(posedge a4454)
   l192 <= a4454;

always @(posedge a4516)
   l194 <= a4516;

always @(posedge a4570)
   l196 <= a4570;

always @(posedge a4572)
   l198 <= a4572;

always @(posedge a4586)
   l200 <= a4586;

always @(posedge na4686)
   l202 <= na4686;

always @(posedge a4698)
   l204 <= a4698;

always @(posedge ni104)
   l206 <= ni104;

always @(posedge na4708)
   l208 <= na4708;

always @(posedge i102)
   l210 <= i102;

always @(posedge i100)
   l212 <= i100;

always @(posedge na4718)
   l214 <= na4718;

always @(posedge na4726)
   l216 <= na4726;

always @(posedge na4732)
   l218 <= na4732;

always @(posedge na4738)
   l220 <= na4738;

always @(posedge na4744)
   l222 <= na4744;

always @(posedge na4750)
   l224 <= na4750;

always @(posedge na4756)
   l226 <= na4756;

always @(posedge na4762)
   l228 <= na4762;

always @(posedge na4768)
   l230 <= na4768;

always @(posedge na4774)
   l232 <= na4774;

always @(posedge ni108)
   l234 <= ni108;

always @(posedge ni116)
   l236 <= ni116;


assign na1780 = ~a1780;
assign a3436 = ~a3434 & ~i2;
assign a3566 = ~a3564 & ~i2;
assign a3590 = ~a3588 & ~i2;
assign na4050 = ~a4050;
assign na4058 = ~a4058;
assign na4066 = ~a4066;
assign na4074 = ~a4074;
assign na4082 = ~a4082;
assign na4090 = ~a4090;
assign na4098 = ~a4098;
assign na4106 = ~a4106;
assign na4114 = ~a4114;
assign na4122 = ~a4122;
assign a4124 = ~i98 & ~i2;
assign a4126 = ~i96 & ~i2;
assign a4128 = ~i94 & ~i2;
assign a4130 = ~i92 & ~i2;
assign a4132 = ~i90 & ~i2;
assign a4134 = l198 & ~i2;
assign a4136 = l190 & ~i2;
assign a4138 = l192 & ~i2;
assign a4140 = l184 & ~i2;
assign a4142 = l178 & ~i2;
assign a4144 = ~i86 & ~i2;
assign a4402 = ~a4400 & ~i2;
assign a4446 = ~a4444 & ~i2;
assign a4448 = ~i84 & ~i2;
assign a4450 = l158 & ~i2;
assign a4452 = l160 & ~i2;
assign a4454 = ~i80 & ~i2;
assign a4516 = ~a4514 & ~i2;
assign a4570 = ~a4568 & ~i2;
assign a4572 = ~i88 & ~i2;
assign a4586 = ~a4584 & ~a4578;
assign na4686 = ~a4686;
assign a4698 = a4696 & a4676;
assign ni104 = ~i104;
assign na4708 = ~a4708;
assign na4718 = ~a4718;
assign na4726 = ~a4726;
assign na4732 = ~a4732;
assign na4738 = ~a4738;
assign na4744 = ~a4744;
assign na4750 = ~a4750;
assign na4756 = ~a4756;
assign na4762 = ~a4762;
assign na4768 = ~a4768;
assign na4774 = ~a4774;
assign ni108 = ~i108;
assign ni116 = ~i116;
assign a238 = ~i8 & ~i6;
assign a240 = ~i12 & i10;
assign a242 = a240 & a238;
assign a244 = a242 & i4;
assign a246 = a244 & l126;
assign a248 = ~l144 & ~l142;
assign a250 = a248 & ~l140;
assign a252 = ~l150 & ~l148;
assign a254 = a252 & ~l146;
assign a256 = ~l156 & ~l154;
assign a258 = a256 & ~l152;
assign a260 = a258 & a254;
assign a262 = a260 & a250;
assign a264 = a262 & ~l138;
assign a266 = ~a264 & ~i22;
assign a268 = l126 & ~i32;
assign a270 = a268 & ~a266;
assign a272 = a270 & i34;
assign a274 = a272 & l166;
assign a276 = a266 & l156;
assign a278 = ~i26 & ~i24;
assign a280 = a278 & ~i28;
assign a282 = ~a268 & ~a266;
assign a284 = a282 & i30;
assign a286 = a284 & a280;
assign a288 = ~a286 & ~a276;
assign a290 = ~a288 & i52;
assign a292 = ~a290 & ~a274;
assign a294 = i26 & i24;
assign a296 = a294 & i28;
assign a298 = a282 & ~i30;
assign a300 = a298 & a296;
assign a302 = l182 & i36;
assign a304 = a302 & l180;
assign a306 = a304 & a270;
assign a308 = ~a306 & ~a300;
assign a310 = ~a308 & l172;
assign a312 = i26 & ~i24;
assign a314 = a312 & i28;
assign a316 = a314 & a298;
assign a318 = l182 & ~i36;
assign a320 = a318 & l180;
assign a322 = a320 & a270;
assign a324 = ~a322 & ~a316;
assign a326 = ~a324 & l174;
assign a328 = ~a326 & ~a310;
assign a330 = a328 & a292;
assign a332 = ~i26 & i24;
assign a334 = a332 & i28;
assign a336 = a334 & a298;
assign a338 = ~l182 & i36;
assign a340 = a338 & l180;
assign a342 = a340 & a270;
assign a344 = ~a342 & ~a336;
assign a346 = ~a344 & l176;
assign a348 = a278 & i28;
assign a350 = a348 & a298;
assign a352 = ~l182 & ~i36;
assign a354 = a352 & l180;
assign a356 = a354 & a270;
assign a358 = ~a356 & ~a350;
assign a360 = ~a358 & l186;
assign a362 = ~a360 & ~a346;
assign a364 = a294 & ~i28;
assign a366 = a364 & a298;
assign a368 = ~l180 & ~i34;
assign a370 = a368 & a302;
assign a372 = a370 & a270;
assign a374 = ~a372 & ~a366;
assign a376 = ~a374 & l188;
assign a378 = a312 & ~i28;
assign a380 = a378 & a298;
assign a382 = a368 & a318;
assign a384 = a382 & a270;
assign a386 = ~a384 & ~a380;
assign a388 = ~a386 & i40;
assign a390 = a266 & l138;
assign a392 = a390 & l168;
assign a394 = ~a392 & ~a388;
assign a396 = a394 & ~a376;
assign a398 = a396 & a362;
assign a400 = a398 & a330;
assign a402 = a266 & l140;
assign a404 = a402 & l170;
assign a406 = a296 & a284;
assign a408 = a266 & l144;
assign a410 = ~a408 & ~a406;
assign a412 = ~a410 & l172;
assign a414 = ~a412 & ~a404;
assign a416 = a266 & l142;
assign a418 = a314 & a284;
assign a420 = ~a418 & ~a416;
assign a422 = ~a420 & l174;
assign a424 = a266 & l146;
assign a426 = a334 & a284;
assign a428 = ~a426 & ~a424;
assign a430 = ~a428 & l176;
assign a432 = a348 & a284;
assign a434 = a266 & l148;
assign a436 = ~a434 & ~a432;
assign a438 = ~a436 & l186;
assign a440 = ~a438 & ~a430;
assign a442 = a440 & ~a422;
assign a444 = a442 & a414;
assign a446 = a364 & a284;
assign a448 = a266 & l150;
assign a450 = ~a448 & ~a446;
assign a452 = ~a450 & l188;
assign a454 = a378 & a284;
assign a456 = a266 & l152;
assign a458 = ~a456 & ~a454;
assign a460 = ~a458 & i40;
assign a462 = ~a460 & ~a452;
assign a464 = a298 & a280;
assign a466 = a368 & a352;
assign a468 = a466 & a270;
assign a470 = ~a468 & ~a464;
assign a472 = ~a470 & i52;
assign a474 = a332 & ~i28;
assign a476 = a474 & a284;
assign a478 = a266 & l154;
assign a480 = ~a478 & ~a476;
assign a482 = a474 & a298;
assign a484 = a368 & a338;
assign a486 = a484 & a270;
assign a488 = ~a486 & ~a482;
assign a490 = a488 & a480;
assign a492 = ~a490 & i42;
assign a494 = ~a492 & ~a472;
assign a496 = a494 & a462;
assign a498 = a496 & a444;
assign a500 = a498 & a400;
assign a502 = a272 & l164;
assign a504 = ~a288 & i42;
assign a506 = ~a504 & ~a502;
assign a508 = ~a308 & l166;
assign a510 = ~a324 & l172;
assign a512 = ~a510 & ~a508;
assign a514 = a512 & a506;
assign a516 = ~a344 & l174;
assign a518 = ~a358 & l176;
assign a520 = ~a518 & ~a516;
assign a522 = ~a374 & l186;
assign a524 = ~a386 & l188;
assign a526 = a390 & l166;
assign a528 = ~a526 & ~a524;
assign a530 = a528 & ~a522;
assign a532 = a530 & a520;
assign a534 = a532 & a514;
assign a536 = a402 & l168;
assign a538 = ~a410 & l170;
assign a540 = ~a538 & ~a536;
assign a542 = ~a420 & l172;
assign a544 = ~a428 & l174;
assign a546 = ~a436 & l176;
assign a548 = ~a546 & ~a544;
assign a550 = a548 & ~a542;
assign a552 = a550 & a540;
assign a554 = ~a450 & l186;
assign a556 = ~a458 & l188;
assign a558 = ~a556 & ~a554;
assign a560 = ~a470 & i42;
assign a562 = ~a490 & i40;
assign a564 = ~a562 & ~a560;
assign a566 = a564 & a558;
assign a568 = a566 & a552;
assign a570 = a568 & a534;
assign a572 = ~a570 & ~a500;
assign a574 = ~a572 & i64;
assign a576 = a570 & a500;
assign a578 = ~a576 & ~i64;
assign a580 = ~a578 & ~a574;
assign a582 = a272 & l192;
assign a584 = ~a288 & l172;
assign a586 = ~a584 & ~a582;
assign a588 = ~a308 & l184;
assign a590 = ~a324 & l178;
assign a592 = ~a590 & ~a588;
assign a594 = a592 & a586;
assign a596 = ~a344 & l158;
assign a598 = ~a358 & l160;
assign a600 = ~a598 & ~a596;
assign a602 = ~a374 & l162;
assign a604 = ~a386 & l164;
assign a606 = a390 & l184;
assign a608 = ~a606 & ~a604;
assign a610 = a608 & ~a602;
assign a612 = a610 & a600;
assign a614 = a612 & a594;
assign a616 = a402 & l178;
assign a618 = ~a410 & l158;
assign a620 = ~a618 & ~a616;
assign a622 = ~a420 & l160;
assign a624 = ~a428 & l162;
assign a626 = ~a436 & l164;
assign a628 = ~a626 & ~a624;
assign a630 = a628 & ~a622;
assign a632 = a630 & a620;
assign a634 = ~a450 & l166;
assign a636 = ~a458 & l168;
assign a638 = ~a636 & ~a634;
assign a640 = ~a480 & l170;
assign a642 = ~a488 & l166;
assign a644 = ~a470 & l172;
assign a646 = ~a644 & ~a642;
assign a648 = a646 & ~a640;
assign a650 = a648 & a638;
assign a652 = a650 & a632;
assign a654 = a652 & a614;
assign a656 = a272 & l184;
assign a658 = ~a288 & l174;
assign a660 = ~a658 & ~a656;
assign a662 = ~a308 & l178;
assign a664 = ~a324 & l158;
assign a666 = ~a664 & ~a662;
assign a668 = a666 & a660;
assign a670 = ~a344 & l160;
assign a672 = ~a358 & l162;
assign a674 = ~a672 & ~a670;
assign a676 = ~a374 & l164;
assign a678 = ~a386 & l166;
assign a680 = a390 & l178;
assign a682 = ~a680 & ~a678;
assign a684 = a682 & ~a676;
assign a686 = a684 & a674;
assign a688 = a686 & a668;
assign a690 = a402 & l158;
assign a692 = ~a410 & l160;
assign a694 = ~a692 & ~a690;
assign a696 = ~a420 & l162;
assign a698 = ~a428 & l164;
assign a700 = ~a436 & l166;
assign a702 = ~a700 & ~a698;
assign a704 = a702 & ~a696;
assign a706 = a704 & a694;
assign a708 = ~a450 & l168;
assign a710 = ~a458 & l170;
assign a712 = ~a710 & ~a708;
assign a714 = ~a470 & l174;
assign a716 = ~a490 & l172;
assign a718 = ~a716 & ~a714;
assign a720 = a718 & a712;
assign a722 = a720 & a706;
assign a724 = a722 & a688;
assign a726 = ~a724 & ~a654;
assign a728 = ~a726 & i64;
assign a730 = a724 & a654;
assign a732 = ~a730 & ~i64;
assign a734 = ~a732 & ~a728;
assign a736 = a734 & a580;
assign a738 = a272 & l162;
assign a740 = ~a288 & i40;
assign a742 = ~a740 & ~a738;
assign a744 = ~a308 & l164;
assign a746 = ~a324 & l166;
assign a748 = ~a746 & ~a744;
assign a750 = a748 & a742;
assign a752 = ~a344 & l172;
assign a754 = ~a358 & l174;
assign a756 = ~a754 & ~a752;
assign a758 = ~a374 & l176;
assign a760 = ~a386 & l186;
assign a762 = a390 & l164;
assign a764 = ~a762 & ~a760;
assign a766 = a764 & ~a758;
assign a768 = a766 & a756;
assign a770 = a768 & a750;
assign a772 = a402 & l166;
assign a774 = ~a410 & l168;
assign a776 = ~a774 & ~a772;
assign a778 = ~a420 & l170;
assign a780 = ~a428 & l172;
assign a782 = ~a436 & l174;
assign a784 = ~a782 & ~a780;
assign a786 = a784 & ~a778;
assign a788 = a786 & a776;
assign a790 = ~a450 & l176;
assign a792 = ~a458 & l186;
assign a794 = ~a792 & ~a790;
assign a796 = ~a470 & i40;
assign a798 = ~a490 & l188;
assign a800 = ~a798 & ~a796;
assign a802 = a800 & a794;
assign a804 = a802 & a788;
assign a806 = a804 & a770;
assign a808 = a272 & l160;
assign a810 = ~a288 & l188;
assign a812 = ~a810 & ~a808;
assign a814 = ~a308 & l162;
assign a816 = ~a324 & l164;
assign a818 = ~a816 & ~a814;
assign a820 = a818 & a812;
assign a822 = ~a344 & l166;
assign a824 = ~a358 & l172;
assign a826 = ~a824 & ~a822;
assign a828 = ~a374 & l174;
assign a830 = ~a386 & l176;
assign a832 = a390 & l162;
assign a834 = ~a832 & ~a830;
assign a836 = a834 & ~a828;
assign a838 = a836 & a826;
assign a840 = a838 & a820;
assign a842 = a402 & l164;
assign a844 = ~a410 & l166;
assign a846 = ~a844 & ~a842;
assign a848 = ~a420 & l168;
assign a850 = ~a428 & l170;
assign a852 = ~a436 & l172;
assign a854 = ~a852 & ~a850;
assign a856 = a854 & ~a848;
assign a858 = a856 & a846;
assign a860 = ~a450 & l174;
assign a862 = ~a458 & l176;
assign a864 = ~a862 & ~a860;
assign a866 = ~a470 & l188;
assign a868 = ~a490 & l186;
assign a870 = ~a868 & ~a866;
assign a872 = a870 & a864;
assign a874 = a872 & a858;
assign a876 = a874 & a840;
assign a878 = a876 & a806;
assign a880 = a272 & l178;
assign a882 = ~a288 & l176;
assign a884 = ~a882 & ~a880;
assign a886 = ~a308 & l158;
assign a888 = ~a324 & l160;
assign a890 = ~a888 & ~a886;
assign a892 = a890 & a884;
assign a894 = ~a344 & l162;
assign a896 = ~a358 & l164;
assign a898 = ~a896 & ~a894;
assign a900 = ~a374 & l166;
assign a902 = ~a386 & l172;
assign a904 = a390 & l158;
assign a906 = ~a904 & ~a902;
assign a908 = a906 & ~a900;
assign a910 = a908 & a898;
assign a912 = a910 & a892;
assign a914 = a402 & l160;
assign a916 = ~a410 & l162;
assign a918 = ~a916 & ~a914;
assign a920 = ~a420 & l164;
assign a922 = ~a428 & l166;
assign a924 = ~a436 & l168;
assign a926 = ~a924 & ~a922;
assign a928 = a926 & ~a920;
assign a930 = a928 & a918;
assign a932 = ~a450 & l170;
assign a934 = ~a458 & l172;
assign a936 = ~a934 & ~a932;
assign a938 = ~a470 & l176;
assign a940 = ~a490 & l174;
assign a942 = ~a940 & ~a938;
assign a944 = a942 & a936;
assign a946 = a944 & a930;
assign a948 = a946 & a912;
assign a950 = a272 & l158;
assign a952 = ~a288 & l186;
assign a954 = ~a952 & ~a950;
assign a956 = ~a308 & l160;
assign a958 = ~a324 & l162;
assign a960 = ~a958 & ~a956;
assign a962 = a960 & a954;
assign a964 = ~a344 & l164;
assign a966 = ~a358 & l166;
assign a968 = ~a966 & ~a964;
assign a970 = ~a374 & l172;
assign a972 = ~a386 & l174;
assign a974 = a390 & l160;
assign a976 = ~a974 & ~a972;
assign a978 = a976 & ~a970;
assign a980 = a978 & a968;
assign a982 = a980 & a962;
assign a984 = a402 & l162;
assign a986 = ~a410 & l164;
assign a988 = ~a986 & ~a984;
assign a990 = ~a420 & l166;
assign a992 = ~a428 & l168;
assign a994 = ~a436 & l170;
assign a996 = ~a994 & ~a992;
assign a998 = a996 & ~a990;
assign a1000 = a998 & a988;
assign a1002 = ~a450 & l172;
assign a1004 = ~a458 & l174;
assign a1006 = ~a1004 & ~a1002;
assign a1008 = ~a470 & l186;
assign a1010 = ~a490 & l176;
assign a1012 = ~a1010 & ~a1008;
assign a1014 = a1012 & a1006;
assign a1016 = a1014 & a1000;
assign a1018 = a1016 & a982;
assign a1020 = a1018 & a948;
assign a1022 = a1020 & a878;
assign a1024 = ~a1022 & ~i64;
assign a1026 = ~a876 & ~a806;
assign a1028 = ~a1018 & ~a948;
assign a1030 = a1028 & a1026;
assign a1032 = ~a1030 & i64;
assign a1034 = ~a1032 & ~a1024;
assign a1036 = a1034 & a736;
assign a1038 = ~a1036 & ~i62;
assign a1040 = ~a1038 & i118;
assign a1042 = a1040 & a246;
assign a1044 = ~i72 & ~i70;
assign a1046 = a1044 & ~l196;
assign a1048 = i76 & i74;
assign a1050 = ~a1048 & a1046;
assign a1052 = ~a1050 & l194;
assign a1054 = ~i12 & ~i10;
assign a1056 = a1054 & a238;
assign a1058 = a1056 & i4;
assign a1060 = a1058 & l126;
assign a1062 = a1028 & a726;
assign a1064 = a1062 & a1026;
assign a1066 = a1064 & a576;
assign a1068 = a1066 & a1060;
assign a1070 = a1068 & a1052;
assign a1072 = a1046 & ~i74;
assign a1074 = a1072 & ~i76;
assign a1076 = a1074 & ~i78;
assign a1078 = ~a1076 & l194;
assign a1080 = a878 & a576;
assign a1082 = a724 & ~a654;
assign a1084 = a1082 & a1020;
assign a1086 = a1084 & a1080;
assign a1088 = a1086 & a1060;
assign a1090 = a1088 & a1078;
assign a1092 = ~a1072 & l194;
assign a1094 = i12 & ~i10;
assign a1096 = a1094 & a238;
assign a1098 = a1096 & ~i4;
assign a1100 = a1098 & l126;
assign a1102 = a1020 & a730;
assign a1104 = a1026 & a572;
assign a1106 = a1104 & a1102;
assign a1108 = a1106 & a1100;
assign a1110 = a1108 & a1092;
assign a1112 = ~a1110 & ~a1090;
assign a1114 = a1112 & ~a1070;
assign a1116 = i78 & i76;
assign a1118 = a1116 & i74;
assign a1120 = ~a1118 & a1046;
assign a1122 = ~a1120 & l194;
assign a1124 = a1102 & a878;
assign a1126 = a570 & ~a500;
assign a1128 = a1126 & a1124;
assign a1130 = a1128 & a1100;
assign a1132 = a1130 & a1122;
assign a1134 = ~i78 & ~i76;
assign a1136 = ~a1134 & i74;
assign a1138 = ~a1136 & a1046;
assign a1140 = ~a1138 & l194;
assign a1142 = ~a876 & a806;
assign a1144 = a1142 & a1062;
assign a1146 = a1144 & a576;
assign a1148 = a1146 & a1060;
assign a1150 = a1148 & a1140;
assign a1152 = ~a1150 & ~a1132;
assign a1154 = a1152 & a1114;
assign a1156 = a1154 & ~a1042;
assign a1158 = a876 & ~a806;
assign a1160 = a1158 & a1102;
assign a1162 = a1160 & a572;
assign a1164 = a1162 & a1100;
assign a1166 = a1164 & a1140;
assign a1168 = ~a1116 & a1072;
assign a1170 = ~a1168 & l194;
assign a1172 = ~a948 & a726;
assign a1174 = a1172 & a1018;
assign a1176 = a1174 & a1080;
assign a1178 = a1176 & a1060;
assign a1180 = a1178 & a1170;
assign a1182 = ~a1180 & ~a1166;
assign a1184 = ~a570 & a500;
assign a1186 = a1184 & a1064;
assign a1188 = a1186 & a1060;
assign a1190 = a1188 & a1122;
assign a1192 = ~a724 & a654;
assign a1194 = a1192 & a1028;
assign a1196 = a1194 & a1104;
assign a1198 = a1196 & a1100;
assign a1200 = a1198 & a1078;
assign a1202 = a1080 & a1062;
assign a1204 = a1202 & a1060;
assign a1206 = a1204 & a1092;
assign a1208 = ~a1206 & ~a1200;
assign a1210 = a1208 & ~a1190;
assign a1212 = a1210 & a1182;
assign a1214 = a1124 & a572;
assign a1216 = a1214 & a1100;
assign a1218 = a1216 & a1052;
assign a1220 = a948 & a730;
assign a1222 = a1220 & ~a1018;
assign a1224 = a1222 & a1104;
assign a1226 = a1224 & a1100;
assign a1228 = a1226 & a1170;
assign a1230 = ~a1228 & ~a1218;
assign a1232 = ~a1074 & l194;
assign a1234 = a1028 & a730;
assign a1236 = a1234 & a1104;
assign a1238 = a1236 & a1100;
assign a1240 = a1238 & a1232;
assign a1242 = ~a1046 & l194;
assign a1244 = a1104 & a1062;
assign a1246 = a1244 & a1060;
assign a1248 = a1246 & a1242;
assign a1250 = ~a1248 & ~a1240;
assign a1252 = a1020 & a726;
assign a1254 = a1252 & a1080;
assign a1256 = a1254 & a1060;
assign a1258 = a1256 & a1232;
assign a1260 = a1102 & a1080;
assign a1262 = a1260 & a1100;
assign a1264 = a1262 & a1242;
assign a1266 = ~a1264 & ~a1258;
assign a1268 = a1266 & a1250;
assign a1270 = a1268 & a1230;
assign a1272 = a1270 & a1212;
assign a1274 = a1272 & a1156;
assign a1276 = i8 & ~i6;
assign a1278 = a1276 & a1054;
assign a1280 = a1278 & ~i4;
assign a1282 = a1280 & l126;
assign a1284 = a1282 & l128;
assign a1286 = l136 & l134;
assign a1288 = a242 & ~i4;
assign a1290 = a1288 & l126;
assign a1292 = a1290 & i68;
assign a1294 = a1292 & a1286;
assign a1296 = i12 & i10;
assign a1298 = a1296 & a238;
assign a1300 = a1298 & ~i4;
assign a1302 = a1300 & l126;
assign a1304 = ~a266 & ~i30;
assign a1306 = a500 & i46;
assign a1308 = ~a500 & ~i46;
assign a1310 = ~a1308 & ~a1306;
assign a1312 = a570 & i48;
assign a1314 = ~a570 & ~i48;
assign a1316 = ~a1314 & ~a1312;
assign a1318 = a1316 & a1310;
assign a1320 = a806 & i50;
assign a1322 = ~a806 & ~i50;
assign a1324 = ~a1322 & ~a1320;
assign a1326 = a876 & i20;
assign a1328 = ~a876 & ~i20;
assign a1330 = ~a1328 & ~a1326;
assign a1332 = a1330 & a1324;
assign a1334 = a1332 & a1318;
assign a1336 = a948 & i58;
assign a1338 = ~a948 & ~i58;
assign a1340 = ~a1338 & ~a1336;
assign a1342 = a1018 & i38;
assign a1344 = ~a1018 & ~i38;
assign a1346 = ~a1344 & ~a1342;
assign a1348 = a1346 & a1340;
assign a1350 = a654 & i56;
assign a1352 = ~a654 & ~i56;
assign a1354 = ~a1352 & ~a1350;
assign a1356 = a724 & i60;
assign a1358 = ~a724 & ~i60;
assign a1360 = ~a1358 & ~a1356;
assign a1362 = a1360 & a1354;
assign a1364 = a1362 & a1348;
assign a1366 = a1364 & a1334;
assign a1368 = a1366 & a1304;
assign a1370 = a654 & i58;
assign a1372 = ~a288 & l168;
assign a1374 = a390 & l190;
assign a1376 = ~a1374 & ~a1372;
assign a1378 = a402 & l192;
assign a1380 = ~a410 & l184;
assign a1382 = ~a1380 & ~a1378;
assign a1384 = ~a420 & l178;
assign a1386 = ~a428 & l158;
assign a1388 = ~a436 & l160;
assign a1390 = ~a1388 & ~a1386;
assign a1392 = a1390 & ~a1384;
assign a1394 = a1392 & a1382;
assign a1396 = ~a450 & l162;
assign a1398 = ~a458 & l164;
assign a1400 = ~a1398 & ~a1396;
assign a1402 = ~a480 & l166;
assign a1404 = ~a1402 & a1400;
assign a1406 = a1404 & a1394;
assign a1408 = a1406 & a1376;
assign a1410 = a1408 & i56;
assign a1412 = ~a1410 & ~a1370;
assign a1414 = ~a948 & ~i20;
assign a1416 = ~a724 & ~i38;
assign a1418 = ~a1416 & ~a1414;
assign a1420 = a1418 & a1412;
assign a1422 = a1018 & i50;
assign a1424 = a876 & i48;
assign a1426 = ~a1424 & ~a1422;
assign a1428 = ~a1018 & ~i50;
assign a1430 = ~a876 & ~i48;
assign a1432 = ~a1430 & ~a1428;
assign a1434 = a1432 & a1426;
assign a1436 = a1434 & a1420;
assign a1438 = a570 & i44;
assign a1440 = a806 & i46;
assign a1442 = ~a1440 & ~a1438;
assign a1444 = ~a500 & ~i54;
assign a1446 = a500 & i54;
assign a1448 = ~a1446 & ~a1304;
assign a1450 = a1448 & ~a1444;
assign a1452 = a1450 & a1442;
assign a1454 = ~a288 & l170;
assign a1456 = a390 & l192;
assign a1458 = ~a1456 & ~a1454;
assign a1460 = a402 & l184;
assign a1462 = ~a410 & l178;
assign a1464 = ~a1462 & ~a1460;
assign a1466 = ~a420 & l158;
assign a1468 = ~a428 & l160;
assign a1470 = ~a436 & l162;
assign a1472 = ~a1470 & ~a1468;
assign a1474 = a1472 & ~a1466;
assign a1476 = a1474 & a1464;
assign a1478 = ~a450 & l164;
assign a1480 = ~a458 & l166;
assign a1482 = ~a1480 & ~a1478;
assign a1484 = ~a480 & l168;
assign a1486 = ~a1484 & a1482;
assign a1488 = a1486 & a1476;
assign a1490 = a1488 & a1458;
assign a1492 = a1490 & i60;
assign a1494 = ~a1490 & ~i60;
assign a1496 = ~a1494 & ~a1492;
assign a1498 = ~a570 & ~i44;
assign a1500 = ~a806 & ~i46;
assign a1502 = ~a1500 & ~a1498;
assign a1504 = a1502 & a1496;
assign a1506 = a948 & i20;
assign a1508 = a724 & i38;
assign a1510 = ~a1508 & ~a1506;
assign a1512 = ~a654 & ~i58;
assign a1514 = ~a1408 & ~i56;
assign a1516 = ~a1514 & ~a1512;
assign a1518 = a1516 & a1510;
assign a1520 = a1518 & a1504;
assign a1522 = a1520 & a1452;
assign a1524 = a1522 & a1436;
assign a1526 = ~a1524 & ~a1368;
assign a1528 = ~a1526 & a1302;
assign a1530 = a1528 & a1286;
assign a1532 = ~a1530 & ~a1294;
assign a1534 = a1532 & ~a1284;
assign a1536 = a1534 & a1274;
assign a1538 = ~a1536 & ~i2;
assign a1540 = ~l128 & i14;
assign a1542 = a1540 & ~l130;
assign a1544 = a1542 & ~i16;
assign a1546 = ~l128 & ~i18;
assign a1548 = l130 & i14;
assign a1550 = a1548 & a1546;
assign a1552 = a1550 & a1282;
assign a1554 = a1546 & l132;
assign a1556 = a1554 & a1282;
assign a1558 = a1056 & ~i4;
assign a1560 = a1558 & l126;
assign a1562 = a1560 & ~i32;
assign a1564 = a1562 & a654;
assign a1566 = ~a1564 & ~a1556;
assign a1568 = a1566 & ~a1552;
assign a1570 = a1568 & ~a1544;
assign a1572 = ~a1570 & ~i2;
assign a1574 = ~a1572 & ~a1538;
assign a1576 = a1096 & i4;
assign a1578 = a1576 & l126;
assign a1580 = a1578 & i66;
assign a1582 = a1130 & ~a1122;
assign a1584 = ~a1244 & ~a1196;
assign a1586 = ~a1236 & ~a1224;
assign a1588 = a1586 & a1584;
assign a1590 = ~a1162 & ~a1106;
assign a1592 = ~a1184 & a1124;
assign a1594 = ~a1592 & a1590;
assign a1596 = a1594 & a1588;
assign a1598 = a1596 & a1100;
assign a1600 = ~a1598 & ~a1582;
assign a1602 = a1300 & ~l126;
assign a1604 = a1216 & ~a1052;
assign a1606 = ~a1604 & ~a1602;
assign a1608 = a1606 & a1600;
assign a1610 = a244 & ~l126;
assign a1612 = a1108 & ~a1092;
assign a1614 = ~a1612 & ~a1610;
assign a1616 = a1164 & ~a1140;
assign a1618 = a1226 & ~a1170;
assign a1620 = a1198 & ~a1078;
assign a1622 = ~a1620 & ~a1618;
assign a1624 = a1622 & ~a1616;
assign a1626 = a1624 & a1614;
assign a1628 = a1626 & a1608;
assign a1630 = a1098 & ~l126;
assign a1632 = ~i8 & i6;
assign a1634 = a1632 & a1054;
assign a1636 = a1634 & i4;
assign a1638 = a1636 & ~l126;
assign a1640 = ~a1638 & ~a1630;
assign a1642 = a1238 & ~a1232;
assign a1644 = a1634 & ~i4;
assign a1646 = a1644 & ~l126;
assign a1648 = ~a1646 & ~a1642;
assign a1650 = a1648 & a1640;
assign a1652 = a1288 & ~l126;
assign a1654 = ~a1260 & ~a1086;
assign a1656 = ~a1254 & ~a1176;
assign a1658 = a1656 & a1654;
assign a1660 = ~a1202 & ~a1146;
assign a1662 = ~a1126 & a1064;
assign a1664 = ~a1662 & a1660;
assign a1666 = a1664 & a1658;
assign a1668 = a1666 & a1060;
assign a1670 = ~a1668 & ~a1652;
assign a1672 = a1292 & ~a1286;
assign a1674 = a1296 & a1276;
assign a1676 = a1674 & ~l126;
assign a1678 = ~a1676 & ~a1672;
assign a1680 = a1678 & a1670;
assign a1682 = a1680 & a1650;
assign a1684 = a1682 & a1628;
assign a1686 = a1188 & ~a1122;
assign a1688 = a1054 & ~i4;
assign a1690 = ~a1688 & ~a240;
assign a1692 = ~a1690 & a1276;
assign a1694 = a1692 & ~l126;
assign a1696 = ~a1694 & ~a1686;
assign a1698 = a1058 & ~l126;
assign a1700 = a1148 & ~a1140;
assign a1702 = ~a1700 & ~a1698;
assign a1704 = a1276 & a1094;
assign a1706 = a1704 & i4;
assign a1708 = a1706 & ~l126;
assign a1710 = a1068 & ~a1052;
assign a1712 = a1204 & ~a1092;
assign a1714 = ~a1712 & ~a1710;
assign a1716 = a1714 & ~a1708;
assign a1718 = a1716 & a1702;
assign a1720 = a1718 & a1696;
assign a1722 = a1256 & ~a1232;
assign a1724 = a1038 & a246;
assign a1726 = ~a1724 & ~a1722;
assign a1728 = ~a1278 & i4;
assign a1730 = ~a1704 & ~i4;
assign a1732 = ~a1730 & ~a1728;
assign a1734 = a1732 & ~l126;
assign a1736 = ~a1734 & a1726;
assign a1738 = a1178 & ~a1170;
assign a1740 = a1088 & ~a1078;
assign a1742 = ~a1740 & ~a1738;
assign a1744 = a1632 & a1094;
assign a1746 = a1744 & ~i4;
assign a1748 = a1298 & i4;
assign a1750 = ~a1748 & ~a1576;
assign a1752 = a1750 & ~a1746;
assign a1754 = ~a1752 & ~l126;
assign a1756 = ~a1754 & a1742;
assign a1758 = a1756 & a1736;
assign a1760 = a1758 & a1720;
assign a1762 = a1760 & a1684;
assign a1764 = a1762 & ~a1560;
assign a1766 = a1764 & ~a1538;
assign a1768 = a1766 & ~a1580;
assign a1770 = a1282 & ~i120;
assign a1772 = a1770 & ~l128;
assign a1774 = ~a1772 & a1768;
assign a1776 = a1774 & ~i2;
assign a1778 = a1776 & i4;
assign a1780 = ~a1778 & a1574;
assign a1782 = a1054 & ~i8;
assign a1784 = ~a1782 & i6;
assign a1786 = ~a1784 & ~l126;
assign a1788 = ~a1786 & ~a238;
assign a1790 = a1788 & i4;
assign a1792 = ~a1556 & ~a1284;
assign a1794 = a1792 & ~a1552;
assign a1796 = a1794 & ~a1544;
assign a1798 = a1748 & l126;
assign a1800 = a250 & ~l146;
assign a1802 = a1800 & l138;
assign a1804 = ~l152 & ~l150;
assign a1806 = a266 & ~l156;
assign a1808 = a1806 & ~l154;
assign a1810 = a1808 & a1804;
assign a1812 = a1810 & ~l148;
assign a1814 = a1812 & a1802;
assign a1816 = a1814 & l158;
assign a1818 = ~l148 & ~l146;
assign a1820 = a1818 & a248;
assign a1822 = a1820 & l140;
assign a1824 = a1822 & a1810;
assign a1826 = a1824 & l160;
assign a1828 = ~a1826 & ~a1816;
assign a1830 = l144 & ~l142;
assign a1832 = a1830 & a1818;
assign a1834 = a1832 & a1810;
assign a1836 = a1834 & l162;
assign a1838 = a416 & a260;
assign a1840 = a1838 & l164;
assign a1842 = ~a1840 & ~a1836;
assign a1844 = a1842 & a1828;
assign a1846 = a424 & a258;
assign a1848 = a1846 & a252;
assign a1850 = a1848 & l166;
assign a1852 = a1810 & l148;
assign a1854 = a1852 & l168;
assign a1856 = ~a1854 & ~a1850;
assign a1858 = ~l152 & l150;
assign a1860 = a1858 & a1808;
assign a1862 = a1860 & l170;
assign a1864 = a1808 & l152;
assign a1866 = a1864 & l172;
assign a1868 = a1806 & l154;
assign a1870 = a1868 & l174;
assign a1872 = ~a1870 & ~a1866;
assign a1874 = a1872 & ~a1862;
assign a1876 = a1874 & a1856;
assign a1878 = a1876 & a1844;
assign a1880 = a276 & l176;
assign a1882 = a300 & l158;
assign a1884 = ~a1882 & ~a1880;
assign a1886 = a316 & l160;
assign a1888 = a336 & l162;
assign a1890 = ~a1888 & ~a1886;
assign a1892 = a1890 & a1884;
assign a1894 = a350 & l164;
assign a1896 = a366 & l166;
assign a1898 = ~a1896 & ~a1894;
assign a1900 = a380 & l172;
assign a1902 = a482 & l174;
assign a1904 = a464 & l176;
assign a1906 = ~a1904 & ~a1902;
assign a1908 = a1906 & ~a1900;
assign a1910 = a1908 & a1898;
assign a1912 = a1910 & a1892;
assign a1914 = a1912 & a1878;
assign a1916 = a406 & l162;
assign a1918 = a418 & l164;
assign a1920 = ~a1918 & ~a1916;
assign a1922 = a426 & l166;
assign a1924 = a432 & l168;
assign a1926 = ~a1924 & ~a1922;
assign a1928 = a446 & l170;
assign a1930 = a454 & l172;
assign a1932 = a476 & l174;
assign a1934 = ~a1932 & ~a1930;
assign a1936 = a1934 & ~a1928;
assign a1938 = a1936 & a1926;
assign a1940 = a1938 & a1920;
assign a1942 = a286 & l176;
assign a1944 = ~a1942 & ~a880;
assign a1946 = a306 & l158;
assign a1948 = a322 & l160;
assign a1950 = a342 & l162;
assign a1952 = ~a1950 & ~a1948;
assign a1954 = a1952 & ~a1946;
assign a1956 = a1954 & a1944;
assign a1958 = a356 & l164;
assign a1960 = a372 & l166;
assign a1962 = ~a1960 & ~a1958;
assign a1964 = a384 & l172;
assign a1966 = a486 & l174;
assign a1968 = a468 & l176;
assign a1970 = ~a1968 & ~a1966;
assign a1972 = a1970 & ~a1964;
assign a1974 = a1972 & a1962;
assign a1976 = a1974 & a1956;
assign a1978 = a1976 & a1940;
assign a1980 = a1978 & a1914;
assign a1982 = ~a1980 & ~i20;
assign a1984 = a1814 & l178;
assign a1986 = a1824 & l158;
assign a1988 = ~a1986 & ~a1984;
assign a1990 = a1834 & l160;
assign a1992 = a1838 & l162;
assign a1994 = ~a1992 & ~a1990;
assign a1996 = a1994 & a1988;
assign a1998 = a1848 & l164;
assign a2000 = a1852 & l166;
assign a2002 = ~a2000 & ~a1998;
assign a2004 = a1860 & l168;
assign a2006 = a1864 & l170;
assign a2008 = a1868 & l172;
assign a2010 = ~a2008 & ~a2006;
assign a2012 = a2010 & ~a2004;
assign a2014 = a2012 & a2002;
assign a2016 = a2014 & a1996;
assign a2018 = a276 & l174;
assign a2020 = a300 & l178;
assign a2022 = ~a2020 & ~a2018;
assign a2024 = a316 & l158;
assign a2026 = a336 & l160;
assign a2028 = ~a2026 & ~a2024;
assign a2030 = a2028 & a2022;
assign a2032 = a350 & l162;
assign a2034 = a366 & l164;
assign a2036 = ~a2034 & ~a2032;
assign a2038 = a380 & l166;
assign a2040 = a482 & l172;
assign a2042 = a464 & l174;
assign a2044 = ~a2042 & ~a2040;
assign a2046 = a2044 & ~a2038;
assign a2048 = a2046 & a2036;
assign a2050 = a2048 & a2030;
assign a2052 = a2050 & a2016;
assign a2054 = a406 & l160;
assign a2056 = a418 & l162;
assign a2058 = ~a2056 & ~a2054;
assign a2060 = a426 & l164;
assign a2062 = a432 & l166;
assign a2064 = ~a2062 & ~a2060;
assign a2066 = a446 & l168;
assign a2068 = a454 & l170;
assign a2070 = a476 & l172;
assign a2072 = ~a2070 & ~a2068;
assign a2074 = a2072 & ~a2066;
assign a2076 = a2074 & a2064;
assign a2078 = a2076 & a2058;
assign a2080 = a286 & l174;
assign a2082 = ~a2080 & ~a656;
assign a2084 = a306 & l178;
assign a2086 = a322 & l158;
assign a2088 = a342 & l160;
assign a2090 = ~a2088 & ~a2086;
assign a2092 = a2090 & ~a2084;
assign a2094 = a2092 & a2082;
assign a2096 = a356 & l162;
assign a2098 = a372 & l164;
assign a2100 = ~a2098 & ~a2096;
assign a2102 = a384 & l166;
assign a2104 = a486 & l172;
assign a2106 = a468 & l174;
assign a2108 = ~a2106 & ~a2104;
assign a2110 = a2108 & ~a2102;
assign a2112 = a2110 & a2100;
assign a2114 = a2112 & a2094;
assign a2116 = a2114 & a2078;
assign a2118 = a2116 & a2052;
assign a2120 = ~a2118 & ~i38;
assign a2122 = ~a2120 & ~a1982;
assign a2124 = a1980 & i20;
assign a2126 = a2118 & i38;
assign a2128 = ~a2126 & ~a2124;
assign a2130 = a2128 & a2122;
assign a2132 = a1814 & l166;
assign a2134 = a1824 & l168;
assign a2136 = ~a2134 & ~a2132;
assign a2138 = a1834 & l170;
assign a2140 = a1838 & l172;
assign a2142 = ~a2140 & ~a2138;
assign a2144 = a2142 & a2136;
assign a2146 = a1848 & l174;
assign a2148 = a1852 & l176;
assign a2150 = ~a2148 & ~a2146;
assign a2152 = a1860 & l186;
assign a2154 = a1864 & l188;
assign a2156 = a1868 & i40;
assign a2158 = ~a2156 & ~a2154;
assign a2160 = a2158 & ~a2152;
assign a2162 = a2160 & a2150;
assign a2164 = a2162 & a2144;
assign a2166 = a276 & i42;
assign a2168 = a300 & l166;
assign a2170 = ~a2168 & ~a2166;
assign a2172 = a316 & l172;
assign a2174 = a336 & l174;
assign a2176 = ~a2174 & ~a2172;
assign a2178 = a2176 & a2170;
assign a2180 = a350 & l176;
assign a2182 = a366 & l186;
assign a2184 = ~a2182 & ~a2180;
assign a2186 = a380 & l188;
assign a2188 = a482 & i40;
assign a2190 = a464 & i42;
assign a2192 = ~a2190 & ~a2188;
assign a2194 = a2192 & ~a2186;
assign a2196 = a2194 & a2184;
assign a2198 = a2196 & a2178;
assign a2200 = a2198 & a2164;
assign a2202 = a406 & l170;
assign a2204 = a418 & l172;
assign a2206 = ~a2204 & ~a2202;
assign a2208 = a426 & l174;
assign a2210 = a432 & l176;
assign a2212 = ~a2210 & ~a2208;
assign a2214 = a446 & l186;
assign a2216 = a454 & l188;
assign a2218 = a476 & i40;
assign a2220 = ~a2218 & ~a2216;
assign a2222 = a2220 & ~a2214;
assign a2224 = a2222 & a2212;
assign a2226 = a2224 & a2206;
assign a2228 = a286 & i42;
assign a2230 = ~a2228 & ~a502;
assign a2232 = a306 & l166;
assign a2234 = a322 & l172;
assign a2236 = a342 & l174;
assign a2238 = ~a2236 & ~a2234;
assign a2240 = a2238 & ~a2232;
assign a2242 = a2240 & a2230;
assign a2244 = a356 & l176;
assign a2246 = a372 & l186;
assign a2248 = ~a2246 & ~a2244;
assign a2250 = a384 & l188;
assign a2252 = a486 & i40;
assign a2254 = a468 & i42;
assign a2256 = ~a2254 & ~a2252;
assign a2258 = a2256 & ~a2250;
assign a2260 = a2258 & a2248;
assign a2262 = a2260 & a2242;
assign a2264 = a2262 & a2226;
assign a2266 = a2264 & a2200;
assign a2268 = ~a2266 & ~i44;
assign a2270 = a1814 & l164;
assign a2272 = a1824 & l166;
assign a2274 = ~a2272 & ~a2270;
assign a2276 = a1834 & l168;
assign a2278 = a1838 & l170;
assign a2280 = ~a2278 & ~a2276;
assign a2282 = a2280 & a2274;
assign a2284 = a1848 & l172;
assign a2286 = a1852 & l174;
assign a2288 = ~a2286 & ~a2284;
assign a2290 = a1860 & l176;
assign a2292 = a1864 & l186;
assign a2294 = a1868 & l188;
assign a2296 = ~a2294 & ~a2292;
assign a2298 = a2296 & ~a2290;
assign a2300 = a2298 & a2288;
assign a2302 = a2300 & a2282;
assign a2304 = a276 & i40;
assign a2306 = a300 & l164;
assign a2308 = ~a2306 & ~a2304;
assign a2310 = a316 & l166;
assign a2312 = a336 & l172;
assign a2314 = ~a2312 & ~a2310;
assign a2316 = a2314 & a2308;
assign a2318 = a350 & l174;
assign a2320 = a366 & l176;
assign a2322 = ~a2320 & ~a2318;
assign a2324 = a380 & l186;
assign a2326 = a482 & l188;
assign a2328 = a464 & i40;
assign a2330 = ~a2328 & ~a2326;
assign a2332 = a2330 & ~a2324;
assign a2334 = a2332 & a2322;
assign a2336 = a2334 & a2316;
assign a2338 = a2336 & a2302;
assign a2340 = a406 & l168;
assign a2342 = a418 & l170;
assign a2344 = ~a2342 & ~a2340;
assign a2346 = a426 & l172;
assign a2348 = a432 & l174;
assign a2350 = ~a2348 & ~a2346;
assign a2352 = a446 & l176;
assign a2354 = a454 & l186;
assign a2356 = a476 & l188;
assign a2358 = ~a2356 & ~a2354;
assign a2360 = a2358 & ~a2352;
assign a2362 = a2360 & a2350;
assign a2364 = a2362 & a2344;
assign a2366 = a286 & i40;
assign a2368 = ~a2366 & ~a738;
assign a2370 = a306 & l164;
assign a2372 = a322 & l166;
assign a2374 = a342 & l172;
assign a2376 = ~a2374 & ~a2372;
assign a2378 = a2376 & ~a2370;
assign a2380 = a2378 & a2368;
assign a2382 = a356 & l174;
assign a2384 = a372 & l176;
assign a2386 = ~a2384 & ~a2382;
assign a2388 = a384 & l186;
assign a2390 = a486 & l188;
assign a2392 = a468 & i40;
assign a2394 = ~a2392 & ~a2390;
assign a2396 = a2394 & ~a2388;
assign a2398 = a2396 & a2386;
assign a2400 = a2398 & a2380;
assign a2402 = a2400 & a2364;
assign a2404 = a2402 & a2338;
assign a2406 = ~a2404 & ~i46;
assign a2408 = ~a2406 & ~a2268;
assign a2410 = a1814 & l162;
assign a2412 = a1824 & l164;
assign a2414 = ~a2412 & ~a2410;
assign a2416 = a1834 & l166;
assign a2418 = a1838 & l168;
assign a2420 = ~a2418 & ~a2416;
assign a2422 = a2420 & a2414;
assign a2424 = a1848 & l170;
assign a2426 = a1852 & l172;
assign a2428 = ~a2426 & ~a2424;
assign a2430 = a1860 & l174;
assign a2432 = a1864 & l176;
assign a2434 = a1868 & l186;
assign a2436 = ~a2434 & ~a2432;
assign a2438 = a2436 & ~a2430;
assign a2440 = a2438 & a2428;
assign a2442 = a2440 & a2422;
assign a2444 = a276 & l188;
assign a2446 = a300 & l162;
assign a2448 = ~a2446 & ~a2444;
assign a2450 = a316 & l164;
assign a2452 = a336 & l166;
assign a2454 = ~a2452 & ~a2450;
assign a2456 = a2454 & a2448;
assign a2458 = a350 & l172;
assign a2460 = a366 & l174;
assign a2462 = ~a2460 & ~a2458;
assign a2464 = a380 & l176;
assign a2466 = a482 & l186;
assign a2468 = a464 & l188;
assign a2470 = ~a2468 & ~a2466;
assign a2472 = a2470 & ~a2464;
assign a2474 = a2472 & a2462;
assign a2476 = a2474 & a2456;
assign a2478 = a2476 & a2442;
assign a2480 = a406 & l166;
assign a2482 = a418 & l168;
assign a2484 = ~a2482 & ~a2480;
assign a2486 = a426 & l170;
assign a2488 = a432 & l172;
assign a2490 = ~a2488 & ~a2486;
assign a2492 = a446 & l174;
assign a2494 = a454 & l176;
assign a2496 = a476 & l186;
assign a2498 = ~a2496 & ~a2494;
assign a2500 = a2498 & ~a2492;
assign a2502 = a2500 & a2490;
assign a2504 = a2502 & a2484;
assign a2506 = a286 & l188;
assign a2508 = ~a2506 & ~a808;
assign a2510 = a306 & l162;
assign a2512 = a322 & l164;
assign a2514 = a342 & l166;
assign a2516 = ~a2514 & ~a2512;
assign a2518 = a2516 & ~a2510;
assign a2520 = a2518 & a2508;
assign a2522 = a356 & l172;
assign a2524 = a372 & l174;
assign a2526 = ~a2524 & ~a2522;
assign a2528 = a384 & l176;
assign a2530 = a486 & l186;
assign a2532 = a468 & l188;
assign a2534 = ~a2532 & ~a2530;
assign a2536 = a2534 & ~a2528;
assign a2538 = a2536 & a2526;
assign a2540 = a2538 & a2520;
assign a2542 = a2540 & a2504;
assign a2544 = a2542 & a2478;
assign a2546 = ~a2544 & ~i48;
assign a2548 = a1814 & l160;
assign a2550 = a1824 & l162;
assign a2552 = ~a2550 & ~a2548;
assign a2554 = a1834 & l164;
assign a2556 = a1838 & l166;
assign a2558 = ~a2556 & ~a2554;
assign a2560 = a2558 & a2552;
assign a2562 = a1848 & l168;
assign a2564 = a1852 & l170;
assign a2566 = ~a2564 & ~a2562;
assign a2568 = a1860 & l172;
assign a2570 = a1864 & l174;
assign a2572 = a1868 & l176;
assign a2574 = ~a2572 & ~a2570;
assign a2576 = a2574 & ~a2568;
assign a2578 = a2576 & a2566;
assign a2580 = a2578 & a2560;
assign a2582 = a276 & l186;
assign a2584 = a300 & l160;
assign a2586 = ~a2584 & ~a2582;
assign a2588 = a316 & l162;
assign a2590 = a336 & l164;
assign a2592 = ~a2590 & ~a2588;
assign a2594 = a2592 & a2586;
assign a2596 = a350 & l166;
assign a2598 = a366 & l172;
assign a2600 = ~a2598 & ~a2596;
assign a2602 = a380 & l174;
assign a2604 = a482 & l176;
assign a2606 = a464 & l186;
assign a2608 = ~a2606 & ~a2604;
assign a2610 = a2608 & ~a2602;
assign a2612 = a2610 & a2600;
assign a2614 = a2612 & a2594;
assign a2616 = a2614 & a2580;
assign a2618 = a406 & l164;
assign a2620 = a418 & l166;
assign a2622 = ~a2620 & ~a2618;
assign a2624 = a426 & l168;
assign a2626 = a432 & l170;
assign a2628 = ~a2626 & ~a2624;
assign a2630 = a446 & l172;
assign a2632 = a454 & l174;
assign a2634 = a476 & l176;
assign a2636 = ~a2634 & ~a2632;
assign a2638 = a2636 & ~a2630;
assign a2640 = a2638 & a2628;
assign a2642 = a2640 & a2622;
assign a2644 = a286 & l186;
assign a2646 = ~a2644 & ~a950;
assign a2648 = a306 & l160;
assign a2650 = a322 & l162;
assign a2652 = a342 & l164;
assign a2654 = ~a2652 & ~a2650;
assign a2656 = a2654 & ~a2648;
assign a2658 = a2656 & a2646;
assign a2660 = a356 & l166;
assign a2662 = a372 & l172;
assign a2664 = ~a2662 & ~a2660;
assign a2666 = a384 & l174;
assign a2668 = a486 & l176;
assign a2670 = a468 & l186;
assign a2672 = ~a2670 & ~a2668;
assign a2674 = a2672 & ~a2666;
assign a2676 = a2674 & a2664;
assign a2678 = a2676 & a2658;
assign a2680 = a2678 & a2642;
assign a2682 = a2680 & a2616;
assign a2684 = ~a2682 & ~i50;
assign a2686 = ~a2684 & ~a2546;
assign a2688 = a2686 & a2408;
assign a2690 = a2688 & a2130;
assign a2692 = a2544 & i48;
assign a2694 = a2682 & i50;
assign a2696 = ~a2694 & ~a2692;
assign a2698 = a2266 & i44;
assign a2700 = a2404 & i46;
assign a2702 = ~a2700 & ~a2698;
assign a2704 = a2702 & a2696;
assign a2706 = a1814 & l168;
assign a2708 = a1824 & l170;
assign a2710 = ~a2708 & ~a2706;
assign a2712 = a1834 & l172;
assign a2714 = a1838 & l174;
assign a2716 = ~a2714 & ~a2712;
assign a2718 = a2716 & a2710;
assign a2720 = a1848 & l176;
assign a2722 = a1852 & l186;
assign a2724 = ~a2722 & ~a2720;
assign a2726 = a1860 & l188;
assign a2728 = a1864 & i40;
assign a2730 = a1868 & i42;
assign a2732 = ~a2730 & ~a2728;
assign a2734 = a2732 & ~a2726;
assign a2736 = a2734 & a2724;
assign a2738 = a2736 & a2718;
assign a2740 = a276 & i52;
assign a2742 = a300 & l172;
assign a2744 = ~a2742 & ~a2740;
assign a2746 = a316 & l174;
assign a2748 = a336 & l176;
assign a2750 = ~a2748 & ~a2746;
assign a2752 = a2750 & a2744;
assign a2754 = a350 & l186;
assign a2756 = a366 & l188;
assign a2758 = ~a2756 & ~a2754;
assign a2760 = a380 & i40;
assign a2762 = a482 & i42;
assign a2764 = a464 & i52;
assign a2766 = ~a2764 & ~a2762;
assign a2768 = a2766 & ~a2760;
assign a2770 = a2768 & a2758;
assign a2772 = a2770 & a2752;
assign a2774 = a2772 & a2738;
assign a2776 = a406 & l172;
assign a2778 = a418 & l174;
assign a2780 = ~a2778 & ~a2776;
assign a2782 = a426 & l176;
assign a2784 = a432 & l186;
assign a2786 = ~a2784 & ~a2782;
assign a2788 = a446 & l188;
assign a2790 = a454 & i40;
assign a2792 = a476 & i42;
assign a2794 = ~a2792 & ~a2790;
assign a2796 = a2794 & ~a2788;
assign a2798 = a2796 & a2786;
assign a2800 = a2798 & a2780;
assign a2802 = a286 & i52;
assign a2804 = ~a2802 & ~a274;
assign a2806 = a306 & l172;
assign a2808 = a322 & l174;
assign a2810 = a342 & l176;
assign a2812 = ~a2810 & ~a2808;
assign a2814 = a2812 & ~a2806;
assign a2816 = a2814 & a2804;
assign a2818 = a356 & l186;
assign a2820 = a372 & l188;
assign a2822 = ~a2820 & ~a2818;
assign a2824 = a384 & i40;
assign a2826 = a486 & i42;
assign a2828 = a468 & i52;
assign a2830 = ~a2828 & ~a2826;
assign a2832 = a2830 & ~a2824;
assign a2834 = a2832 & a2822;
assign a2836 = a2834 & a2816;
assign a2838 = a2836 & a2800;
assign a2840 = a2838 & a2774;
assign a2842 = a2840 & i54;
assign a2844 = ~a2840 & ~i54;
assign a2846 = a1814 & l190;
assign a2848 = a1824 & l192;
assign a2850 = ~a2848 & ~a2846;
assign a2852 = a1834 & l184;
assign a2854 = a1838 & l178;
assign a2856 = a1848 & l158;
assign a2858 = ~a2856 & ~a2854;
assign a2860 = a2858 & ~a2852;
assign a2862 = a2860 & a2850;
assign a2864 = a1852 & l160;
assign a2866 = a1860 & l162;
assign a2868 = ~a2866 & ~a2864;
assign a2870 = a1864 & l164;
assign a2872 = a1868 & l166;
assign a2874 = a276 & l168;
assign a2876 = ~a2874 & ~a2872;
assign a2878 = a2876 & ~a2870;
assign a2880 = a2878 & a2868;
assign a2882 = a2880 & a2862;
assign a2884 = a406 & l184;
assign a2886 = a418 & l178;
assign a2888 = a426 & l158;
assign a2890 = ~a2888 & ~a2886;
assign a2892 = a2890 & ~a2884;
assign a2894 = a432 & l160;
assign a2896 = a446 & l162;
assign a2898 = ~a2896 & ~a2894;
assign a2900 = a454 & l164;
assign a2902 = a476 & l166;
assign a2904 = a286 & l168;
assign a2906 = ~a2904 & ~a2902;
assign a2908 = a2906 & ~a2900;
assign a2910 = a2908 & a2898;
assign a2912 = a2910 & a2892;
assign a2914 = a2912 & a2882;
assign a2916 = ~a2914 & ~i56;
assign a2918 = ~a2916 & ~a2844;
assign a2920 = a2918 & ~a2842;
assign a2922 = a1814 & l184;
assign a2924 = a1824 & l178;
assign a2926 = ~a2924 & ~a2922;
assign a2928 = a1834 & l158;
assign a2930 = a1838 & l160;
assign a2932 = ~a2930 & ~a2928;
assign a2934 = a2932 & a2926;
assign a2936 = a1848 & l162;
assign a2938 = a1852 & l164;
assign a2940 = ~a2938 & ~a2936;
assign a2942 = a1860 & l166;
assign a2944 = a1864 & l168;
assign a2946 = a1868 & l170;
assign a2948 = ~a2946 & ~a2944;
assign a2950 = a2948 & ~a2942;
assign a2952 = a2950 & a2940;
assign a2954 = a2952 & a2934;
assign a2956 = a276 & l172;
assign a2958 = a300 & l184;
assign a2960 = ~a2958 & ~a2956;
assign a2962 = a316 & l178;
assign a2964 = a336 & l158;
assign a2966 = ~a2964 & ~a2962;
assign a2968 = a2966 & a2960;
assign a2970 = a350 & l160;
assign a2972 = a366 & l162;
assign a2974 = ~a2972 & ~a2970;
assign a2976 = a380 & l164;
assign a2978 = a482 & l166;
assign a2980 = a464 & l172;
assign a2982 = ~a2980 & ~a2978;
assign a2984 = a2982 & ~a2976;
assign a2986 = a2984 & a2974;
assign a2988 = a2986 & a2968;
assign a2990 = a2988 & a2954;
assign a2992 = a406 & l158;
assign a2994 = a418 & l160;
assign a2996 = ~a2994 & ~a2992;
assign a2998 = a426 & l162;
assign a3000 = a432 & l164;
assign a3002 = ~a3000 & ~a2998;
assign a3004 = a446 & l166;
assign a3006 = a454 & l168;
assign a3008 = a476 & l170;
assign a3010 = ~a3008 & ~a3006;
assign a3012 = a3010 & ~a3004;
assign a3014 = a3012 & a3002;
assign a3016 = a3014 & a2996;
assign a3018 = a286 & l172;
assign a3020 = ~a3018 & ~a582;
assign a3022 = a306 & l184;
assign a3024 = a322 & l178;
assign a3026 = a342 & l158;
assign a3028 = ~a3026 & ~a3024;
assign a3030 = a3028 & ~a3022;
assign a3032 = a3030 & a3020;
assign a3034 = a356 & l160;
assign a3036 = a372 & l162;
assign a3038 = ~a3036 & ~a3034;
assign a3040 = a384 & l164;
assign a3042 = a486 & l166;
assign a3044 = a468 & l172;
assign a3046 = ~a3044 & ~a3042;
assign a3048 = a3046 & ~a3040;
assign a3050 = a3048 & a3038;
assign a3052 = a3050 & a3032;
assign a3054 = a3052 & a3016;
assign a3056 = a3054 & a2990;
assign a3058 = ~a3056 & ~i58;
assign a3060 = a1814 & l192;
assign a3062 = a1824 & l184;
assign a3064 = ~a3062 & ~a3060;
assign a3066 = a1834 & l178;
assign a3068 = a1838 & l158;
assign a3070 = a1848 & l160;
assign a3072 = ~a3070 & ~a3068;
assign a3074 = a3072 & ~a3066;
assign a3076 = a3074 & a3064;
assign a3078 = a1852 & l162;
assign a3080 = a1860 & l164;
assign a3082 = ~a3080 & ~a3078;
assign a3084 = a1864 & l166;
assign a3086 = a1868 & l168;
assign a3088 = a276 & l170;
assign a3090 = ~a3088 & ~a3086;
assign a3092 = a3090 & ~a3084;
assign a3094 = a3092 & a3082;
assign a3096 = a3094 & a3076;
assign a3098 = a406 & l178;
assign a3100 = a418 & l158;
assign a3102 = a426 & l160;
assign a3104 = ~a3102 & ~a3100;
assign a3106 = a3104 & ~a3098;
assign a3108 = a432 & l162;
assign a3110 = a446 & l164;
assign a3112 = ~a3110 & ~a3108;
assign a3114 = a454 & l166;
assign a3116 = a476 & l168;
assign a3118 = a286 & l170;
assign a3120 = ~a3118 & ~a3116;
assign a3122 = a3120 & ~a3114;
assign a3124 = a3122 & a3112;
assign a3126 = a3124 & a3106;
assign a3128 = a3126 & a3096;
assign a3130 = ~a3128 & ~i60;
assign a3132 = ~a3130 & ~a1304;
assign a3134 = a3132 & ~a3058;
assign a3136 = a3056 & i58;
assign a3138 = a3128 & i60;
assign a3140 = a2914 & i56;
assign a3142 = ~a3140 & ~a3138;
assign a3144 = a3142 & ~a3136;
assign a3146 = a3144 & a3134;
assign a3148 = a3146 & a2920;
assign a3150 = a3148 & a2704;
assign a3152 = a3150 & a2690;
assign a3154 = ~a3152 & ~a1368;
assign a3156 = ~a3154 & a1302;
assign a3158 = a3156 & a1286;
assign a3160 = ~a2682 & ~a1980;
assign a3162 = a2682 & ~i64;
assign a3164 = ~a3162 & ~a3160;
assign a3166 = a2840 & a2266;
assign a3168 = ~a3166 & ~i64;
assign a3170 = ~a3056 & ~a2118;
assign a3172 = ~a3170 & i64;
assign a3174 = ~a3172 & ~a3168;
assign a3176 = a3174 & ~a3164;
assign a3178 = ~a2840 & ~a2266;
assign a3180 = ~a3178 & i64;
assign a3182 = ~a2544 & a2404;
assign a3184 = ~a2404 & ~i64;
assign a3186 = ~a3184 & ~a3182;
assign a3188 = a3186 & ~a3180;
assign a3190 = a2544 & i64;
assign a3192 = a3056 & a2118;
assign a3194 = a3192 & a1980;
assign a3196 = ~a3194 & ~i64;
assign a3198 = ~a3196 & ~a3190;
assign a3200 = a3198 & a3188;
assign a3202 = a3200 & a3176;
assign a3204 = ~a3202 & ~i62;
assign a3206 = ~a3204 & a246;
assign a3208 = ~a3206 & ~a3158;
assign a3210 = a3208 & ~a1798;
assign a3212 = a3210 & a1796;
assign a3214 = a3212 & ~a1790;
assign a3216 = a1578 & ~i66;
assign a3218 = ~a3216 & ~a1294;
assign a3220 = a3166 & a2404;
assign a3222 = a3220 & a2544;
assign a3224 = a3222 & a2682;
assign a3226 = a3224 & a1980;
assign a3228 = a3226 & a2118;
assign a3230 = a3228 & a3056;
assign a3232 = a3230 & a1100;
assign a3234 = a3232 & a1242;
assign a3236 = a3178 & ~a2404;
assign a3238 = a3236 & ~a2544;
assign a3240 = a3238 & a2682;
assign a3242 = a3240 & a3194;
assign a3244 = a3242 & a1100;
assign a3246 = a3244 & a1092;
assign a3248 = a3238 & ~a2682;
assign a3250 = a3248 & a1980;
assign a3252 = a3250 & a1100;
assign a3254 = a3252 & a3192;
assign a3256 = a3254 & a1170;
assign a3258 = a3248 & ~a1980;
assign a3260 = a3258 & a2118;
assign a3262 = a3260 & a1100;
assign a3264 = a3262 & a3056;
assign a3266 = a3264 & a1232;
assign a3268 = ~a3266 & ~a3256;
assign a3270 = a3268 & ~a3246;
assign a3272 = a3236 & a2544;
assign a3274 = a3272 & a3194;
assign a3276 = a3274 & a2682;
assign a3278 = a3276 & a1100;
assign a3280 = a3278 & a1140;
assign a3282 = a2682 & a2544;
assign a3284 = a3178 & a2404;
assign a3286 = a3284 & a1100;
assign a3288 = a3286 & a3282;
assign a3290 = a3288 & a3194;
assign a3292 = a3290 & a1052;
assign a3294 = ~a2840 & a2266;
assign a3296 = a3294 & a3194;
assign a3298 = a3296 & a2404;
assign a3300 = a3298 & a3282;
assign a3302 = a3300 & a1100;
assign a3304 = a3302 & a1122;
assign a3306 = ~a3304 & ~a3292;
assign a3308 = a3306 & ~a3280;
assign a3310 = a3308 & a3270;
assign a3312 = a3310 & ~a3234;
assign a3314 = a3258 & ~a2118;
assign a3316 = a3314 & a1100;
assign a3318 = a3316 & a3056;
assign a3320 = a3318 & a1078;
assign a3322 = a3314 & ~a3056;
assign a3324 = a3322 & a1060;
assign a3326 = a3324 & ~a1242;
assign a3328 = a3230 & a1060;
assign a3330 = ~a3328 & ~a3326;
assign a3332 = a3330 & ~a3320;
assign a3334 = a3332 & a3312;
assign a3336 = a3334 & a3218;
assign a3338 = a3170 & a1060;
assign a3340 = a3338 & ~a1980;
assign a3342 = a3222 & ~a2682;
assign a3344 = a3342 & a3340;
assign a3346 = a3344 & a1092;
assign a3348 = a3340 & a3224;
assign a3350 = a3348 & a1170;
assign a3352 = ~a3350 & ~a3346;
assign a3354 = a2840 & ~a2266;
assign a3356 = ~a2682 & ~a2544;
assign a3358 = a3356 & a3340;
assign a3360 = a3358 & a3354;
assign a3362 = a3360 & ~a2404;
assign a3364 = a3362 & a1122;
assign a3366 = a3166 & ~a2404;
assign a3368 = a3366 & a3358;
assign a3370 = a3368 & a1052;
assign a3372 = a3358 & a3220;
assign a3374 = a3372 & a1140;
assign a3376 = ~a3374 & ~a3370;
assign a3378 = a3376 & ~a3364;
assign a3380 = a3378 & a3352;
assign a3382 = a3324 & a1242;
assign a3384 = ~a3382 & a3380;
assign a3386 = a3338 & a3226;
assign a3388 = a3386 & a1232;
assign a3390 = a3228 & a1060;
assign a3392 = a3390 & ~a3056;
assign a3394 = a3392 & a1078;
assign a3396 = ~a3394 & ~a3388;
assign a3398 = a3230 & a1562;
assign a3400 = ~a3398 & a3396;
assign a3402 = a3400 & a3384;
assign a3404 = a3300 & a1562;
assign a3406 = a3194 & a1562;
assign a3408 = a2404 & a2266;
assign a3410 = a3408 & a2544;
assign a3412 = ~a3410 & a3406;
assign a3414 = a3412 & a2682;
assign a3416 = ~a3414 & ~a3404;
assign a3418 = a3406 & ~a2682;
assign a3420 = a2118 & a1980;
assign a3422 = ~a3420 & a1562;
assign a3424 = a3422 & a3056;
assign a3426 = ~a3424 & ~a3418;
assign a3428 = a3426 & a3416;
assign a3430 = a3428 & a3402;
assign a3432 = a3430 & a3336;
assign a3434 = a3432 & a3214;
assign a3438 = ~a1688 & a238;
assign a3440 = a3438 & ~a1798;
assign a3442 = ~a3440 & l134;
assign a3444 = l136 & ~l134;
assign a3446 = ~l136 & l134;
assign a3448 = ~a3446 & ~a3444;
assign a3450 = ~a3448 & a3156;
assign a3452 = a246 & l134;
assign a3454 = ~a3452 & ~a3450;
assign a3456 = a3454 & ~a3158;
assign a3458 = a3456 & ~a3442;
assign a3460 = a1290 & ~i68;
assign a3462 = a3460 & a1286;
assign a3464 = ~a2840 & ~i46;
assign a3466 = a2840 & i46;
assign a3468 = ~a3466 & ~a3464;
assign a3470 = ~a2266 & ~i48;
assign a3472 = a2266 & i48;
assign a3474 = ~a3472 & ~a3470;
assign a3476 = a3474 & a3468;
assign a3478 = ~a2404 & ~i50;
assign a3480 = a2404 & i50;
assign a3482 = ~a3480 & ~a3478;
assign a3484 = ~a2544 & ~i20;
assign a3486 = a2544 & i20;
assign a3488 = ~a3486 & ~a3484;
assign a3490 = a3488 & a3482;
assign a3492 = a3490 & a3476;
assign a3494 = ~a2682 & ~i38;
assign a3496 = a2682 & i38;
assign a3498 = ~a3496 & ~a3494;
assign a3500 = ~a1980 & ~i58;
assign a3502 = a1980 & i58;
assign a3504 = ~a3502 & ~a3500;
assign a3506 = a3504 & a3498;
assign a3508 = ~a2118 & ~i60;
assign a3510 = a2118 & i60;
assign a3512 = ~a3510 & ~a3508;
assign a3514 = ~a3056 & ~i56;
assign a3516 = a3056 & i56;
assign a3518 = ~a3516 & ~a3514;
assign a3520 = a3518 & a3512;
assign a3522 = a3520 & a3506;
assign a3524 = a3522 & a3492;
assign a3526 = a3524 & ~i64;
assign a3528 = ~a3474 & ~a3468;
assign a3530 = ~a3488 & ~a3482;
assign a3532 = a3530 & a3528;
assign a3534 = ~a3504 & ~a3498;
assign a3536 = ~a3518 & i64;
assign a3538 = a3536 & ~a3512;
assign a3540 = a3538 & a3534;
assign a3542 = a3540 & a3532;
assign a3544 = ~a3542 & ~a3526;
assign a3546 = a3460 & ~a1286;
assign a3548 = a3546 & ~a3544;
assign a3550 = a3548 & ~a3448;
assign a3552 = ~a3550 & ~a1294;
assign a3554 = a3552 & ~a3462;
assign a3556 = ~a1096 & ~a1058;
assign a3558 = ~a3556 & l134;
assign a3560 = a3558 & l126;
assign a3562 = ~a3560 & a3554;
assign a3564 = a3562 & a3458;
assign a3568 = ~a3444 & a3156;
assign a3570 = a3440 & ~a246;
assign a3572 = ~a3570 & l136;
assign a3574 = ~a3572 & ~a3568;
assign a3576 = a3548 & ~l136;
assign a3578 = ~a3576 & ~a1294;
assign a3580 = a3578 & ~a3462;
assign a3582 = ~a3556 & l136;
assign a3584 = a3582 & l126;
assign a3586 = ~a3584 & a3580;
assign a3588 = a3586 & a3574;
assign a3592 = l202 & l200;
assign a3594 = ~l202 & ~l200;
assign a3596 = ~a3594 & ~a3592;
assign a3598 = l206 & l200;
assign a3600 = ~a3598 & l204;
assign a3602 = ~l206 & ~l200;
assign a3604 = ~a3602 & ~l204;
assign a3606 = a3604 & ~l208;
assign a3608 = a3604 & ~a3598;
assign a3610 = ~a3608 & l208;
assign a3612 = ~a3610 & ~a3606;
assign a3614 = a3612 & ~a3600;
assign a3616 = a3614 & a3596;
assign a3618 = l166 & ~l164;
assign a3620 = a3618 & l168;
assign a3622 = ~l166 & l164;
assign a3624 = a3622 & l168;
assign a3626 = ~a3624 & ~a3620;
assign a3628 = ~l176 & ~l174;
assign a3630 = ~l172 & ~l170;
assign a3632 = a3630 & a3628;
assign a3634 = l188 & ~l186;
assign a3636 = a3634 & i40;
assign a3638 = a3636 & a3632;
assign a3640 = a3638 & ~a3626;
assign a3642 = a3622 & ~l168;
assign a3644 = a3618 & ~l168;
assign a3646 = ~a3644 & ~a3642;
assign a3648 = l176 & l174;
assign a3650 = l172 & l170;
assign a3652 = a3650 & a3648;
assign a3654 = ~l188 & l186;
assign a3656 = a3654 & ~i40;
assign a3658 = a3656 & a3652;
assign a3660 = a3658 & ~a3646;
assign a3662 = ~a3660 & ~a3640;
assign a3664 = ~l174 & ~l172;
assign a3666 = ~l170 & ~l168;
assign a3668 = a3666 & a3664;
assign a3670 = l188 & l186;
assign a3672 = a3670 & ~l176;
assign a3674 = a3672 & a3668;
assign a3676 = ~a3674 & l166;
assign a3678 = l174 & l172;
assign a3680 = l170 & l168;
assign a3682 = a3680 & a3678;
assign a3684 = ~l188 & ~l186;
assign a3686 = a3684 & l176;
assign a3688 = a3686 & a3682;
assign a3690 = ~a3688 & ~l166;
assign a3692 = ~a3690 & ~a3676;
assign a3694 = ~l164 & ~l162;
assign a3696 = l164 & l162;
assign a3698 = ~a3696 & ~a3694;
assign a3700 = a3698 & a3692;
assign a3702 = ~l168 & ~l166;
assign a3704 = a3702 & a3630;
assign a3706 = l186 & l176;
assign a3708 = a3706 & ~l174;
assign a3710 = a3708 & a3704;
assign a3712 = ~a3710 & l164;
assign a3714 = l168 & l166;
assign a3716 = a3714 & a3650;
assign a3718 = ~l186 & ~l176;
assign a3720 = a3718 & l174;
assign a3722 = a3720 & a3716;
assign a3724 = ~a3722 & ~l164;
assign a3726 = ~a3724 & ~a3712;
assign a3728 = ~l162 & ~l160;
assign a3730 = l162 & l160;
assign a3732 = ~a3730 & ~a3728;
assign a3734 = a3732 & a3726;
assign a3736 = ~a3734 & ~a3700;
assign a3738 = a3736 & a3662;
assign a3740 = l170 & ~l168;
assign a3742 = a3740 & l172;
assign a3744 = ~l170 & l168;
assign a3746 = a3744 & l172;
assign a3748 = ~a3746 & ~a3742;
assign a3750 = a3684 & a3628;
assign a3752 = i42 & ~i40;
assign a3754 = a3752 & i52;
assign a3756 = a3754 & a3750;
assign a3758 = a3756 & ~a3748;
assign a3760 = a3744 & ~l172;
assign a3762 = a3740 & ~l172;
assign a3764 = ~a3762 & ~a3760;
assign a3766 = a3670 & a3648;
assign a3768 = ~i42 & i40;
assign a3770 = a3768 & ~i52;
assign a3772 = a3770 & a3766;
assign a3774 = a3772 & ~a3764;
assign a3776 = ~a3774 & ~a3758;
assign a3778 = l168 & ~l166;
assign a3780 = a3778 & l170;
assign a3782 = ~l168 & l166;
assign a3784 = a3782 & l170;
assign a3786 = ~a3784 & ~a3780;
assign a3788 = a3718 & a3664;
assign a3790 = ~l188 & i40;
assign a3792 = a3790 & i42;
assign a3794 = a3792 & a3788;
assign a3796 = a3794 & ~a3786;
assign a3798 = a3782 & ~l170;
assign a3800 = a3778 & ~l170;
assign a3802 = ~a3800 & ~a3798;
assign a3804 = a3706 & a3678;
assign a3806 = l188 & ~i40;
assign a3808 = a3806 & ~i42;
assign a3810 = a3808 & a3804;
assign a3812 = a3810 & ~a3802;
assign a3814 = ~a3812 & ~a3796;
assign a3816 = a3814 & a3776;
assign a3818 = a3816 & a3738;
assign a3820 = ~l166 & ~l164;
assign a3822 = a3820 & a3666;
assign a3824 = a3648 & ~l172;
assign a3826 = a3824 & a3822;
assign a3828 = ~a3826 & l162;
assign a3830 = l166 & l164;
assign a3832 = a3830 & a3680;
assign a3834 = a3628 & l172;
assign a3836 = a3834 & a3832;
assign a3838 = ~a3836 & ~l162;
assign a3840 = ~a3838 & ~a3828;
assign a3842 = ~l160 & ~l158;
assign a3844 = l160 & l158;
assign a3846 = ~a3844 & ~a3842;
assign a3848 = a3846 & a3840;
assign a3850 = a3702 & a3694;
assign a3852 = a3678 & ~l170;
assign a3854 = a3852 & a3850;
assign a3856 = ~a3854 & l160;
assign a3858 = a3714 & a3696;
assign a3860 = a3664 & l170;
assign a3862 = a3860 & a3858;
assign a3864 = ~a3862 & ~l160;
assign a3866 = ~a3864 & ~a3856;
assign a3868 = ~l178 & ~l158;
assign a3870 = l178 & l158;
assign a3872 = ~a3870 & ~a3868;
assign a3874 = a3872 & a3866;
assign a3876 = ~a3874 & ~a3848;
assign a3878 = l192 & ~l190;
assign a3880 = ~l192 & l190;
assign a3882 = ~a3880 & ~a3878;
assign a3884 = a3868 & a3728;
assign a3886 = a3884 & a3620;
assign a3888 = ~a3886 & l184;
assign a3890 = a3870 & a3730;
assign a3892 = a3890 & a3642;
assign a3894 = ~a3892 & ~l184;
assign a3896 = ~a3894 & ~a3888;
assign a3898 = a3896 & ~a3882;
assign a3900 = ~l184 & l178;
assign a3902 = l184 & ~l178;
assign a3904 = ~a3902 & ~a3900;
assign a3906 = a3820 & a3728;
assign a3908 = a3906 & a3742;
assign a3910 = ~a3908 & l158;
assign a3912 = a3830 & a3730;
assign a3914 = a3912 & a3760;
assign a3916 = ~a3914 & ~l158;
assign a3918 = ~a3916 & ~a3910;
assign a3920 = a3918 & ~a3904;
assign a3922 = ~l192 & l184;
assign a3924 = l192 & ~l184;
assign a3926 = ~a3924 & ~a3922;
assign a3928 = a3842 & a3694;
assign a3930 = a3928 & a3780;
assign a3932 = ~a3930 & l178;
assign a3934 = a3844 & a3696;
assign a3936 = a3934 & a3798;
assign a3938 = ~a3936 & ~l178;
assign a3940 = ~a3938 & ~a3932;
assign a3942 = a3940 & ~a3926;
assign a3944 = ~a3942 & ~a3920;
assign a3946 = a3944 & ~a3898;
assign a3948 = a3946 & a3876;
assign a3950 = a3948 & ~a3818;
assign a3952 = ~a3948 & a3818;
assign a3954 = ~a3952 & ~a3950;
assign a3956 = ~a3776 & ~l156;
assign a3958 = a3776 & l156;
assign a3960 = ~a3958 & ~a3956;
assign a3962 = ~a3814 & ~l154;
assign a3964 = a3814 & l154;
assign a3966 = ~a3964 & ~a3962;
assign a3968 = a3966 & a3960;
assign a3970 = ~a3662 & ~l152;
assign a3972 = a3662 & l152;
assign a3974 = ~a3972 & ~a3970;
assign a3976 = a3700 & ~l150;
assign a3978 = ~a3700 & l150;
assign a3980 = ~a3978 & ~a3976;
assign a3982 = a3734 & ~l148;
assign a3984 = ~a3734 & l148;
assign a3986 = ~a3984 & ~a3982;
assign a3988 = a3986 & a3980;
assign a3990 = a3988 & a3974;
assign a3992 = a3990 & a3968;
assign a3994 = a3848 & ~l146;
assign a3996 = ~a3848 & l146;
assign a3998 = ~a3996 & ~a3994;
assign a4000 = a3874 & ~l142;
assign a4002 = ~a3874 & l142;
assign a4004 = ~a4002 & ~a4000;
assign a4006 = a4004 & a3998;
assign a4008 = a3920 & ~l144;
assign a4010 = ~a3920 & l144;
assign a4012 = ~a4010 & ~a4008;
assign a4014 = a3942 & ~l140;
assign a4016 = ~a3942 & l140;
assign a4018 = ~a4016 & ~a4014;
assign a4020 = a3898 & ~l138;
assign a4022 = ~a3898 & l138;
assign a4024 = ~a4022 & ~a4020;
assign a4026 = a4024 & a4018;
assign a4028 = a4026 & a4012;
assign a4030 = a4028 & a4006;
assign a4032 = a4030 & a3992;
assign a4034 = a4032 & ~a3954;
assign a4036 = ~a4034 & l212;
assign a4038 = ~a4036 & ~l210;
assign a4040 = ~a4038 & a3616;
assign a4042 = ~a4040 & ~i2;
assign a4044 = a4042 & l138;
assign a4046 = l232 & ~i2;
assign a4048 = a4046 & a4040;
assign a4050 = ~a4048 & ~a4044;
assign a4052 = a4042 & l140;
assign a4054 = l230 & ~i2;
assign a4056 = a4054 & a4040;
assign a4058 = ~a4056 & ~a4052;
assign a4060 = a4042 & l142;
assign a4062 = l226 & ~i2;
assign a4064 = a4062 & a4040;
assign a4066 = ~a4064 & ~a4060;
assign a4068 = a4042 & l144;
assign a4070 = l228 & ~i2;
assign a4072 = a4070 & a4040;
assign a4074 = ~a4072 & ~a4068;
assign a4076 = a4042 & l146;
assign a4078 = l224 & ~i2;
assign a4080 = a4078 & a4040;
assign a4082 = ~a4080 & ~a4076;
assign a4084 = a4042 & l148;
assign a4086 = l222 & ~i2;
assign a4088 = a4086 & a4040;
assign a4090 = ~a4088 & ~a4084;
assign a4092 = a4042 & l150;
assign a4094 = l220 & ~i2;
assign a4096 = a4094 & a4040;
assign a4098 = ~a4096 & ~a4092;
assign a4100 = a4042 & l152;
assign a4102 = l218 & ~i2;
assign a4104 = a4102 & a4040;
assign a4106 = ~a4104 & ~a4100;
assign a4108 = a4042 & l154;
assign a4110 = l216 & ~i2;
assign a4112 = a4110 & a4040;
assign a4114 = ~a4112 & ~a4108;
assign a4116 = a4042 & l156;
assign a4118 = ~l214 & ~i2;
assign a4120 = ~a4118 & ~a4042;
assign a4122 = ~a4120 & ~a4116;
assign a4146 = ~a1098 & ~a1056;
assign a4148 = a3290 & ~a1052;
assign a4150 = a3250 & a3056;
assign a4152 = ~a4150 & ~a3260;
assign a4154 = ~a4152 & ~a3192;
assign a4156 = a3284 & ~a2544;
assign a4158 = a4156 & a2682;
assign a4160 = ~a3294 & ~a2404;
assign a4162 = ~a3354 & a2404;
assign a4164 = ~a4162 & ~a4160;
assign a4166 = a4164 & a3282;
assign a4168 = ~a4166 & ~a4158;
assign a4170 = ~a4168 & a3194;
assign a4172 = a3274 & ~a2682;
assign a4174 = a3240 & ~a3056;
assign a4176 = ~a4174 & ~a4172;
assign a4178 = a4176 & ~a4170;
assign a4180 = a3250 & ~a3056;
assign a4182 = ~a3272 & ~a3192;
assign a4184 = a3284 & ~a1980;
assign a4186 = ~a4184 & a3192;
assign a4188 = ~a4186 & ~a4182;
assign a4190 = ~a4188 & ~a4180;
assign a4192 = a4190 & a4178;
assign a4194 = a4192 & ~a4154;
assign a4196 = a2840 & ~a2404;
assign a4198 = a4196 & a3282;
assign a4200 = ~a3284 & ~a2682;
assign a4202 = a3294 & ~a2544;
assign a4204 = ~a4202 & a2682;
assign a4206 = ~a4204 & ~a4200;
assign a4208 = ~a4206 & ~a4198;
assign a4210 = ~a4208 & a3194;
assign a4212 = ~a4210 & ~a3322;
assign a4214 = ~a3178 & ~a2682;
assign a4216 = a4214 & a3194;
assign a4218 = ~a3356 & a3236;
assign a4220 = a4218 & ~a1980;
assign a4222 = a4220 & a3192;
assign a4224 = ~a4222 & ~a4216;
assign a4226 = a3240 & ~a2118;
assign a4228 = a4226 & a3056;
assign a4230 = a2840 & ~a2544;
assign a4232 = a4230 & a2682;
assign a4234 = a4232 & a3194;
assign a4236 = a3294 & ~a1980;
assign a4238 = a4236 & a3192;
assign a4240 = ~a4238 & ~a4234;
assign a4242 = a2840 & ~a2118;
assign a4244 = a4242 & a3056;
assign a4246 = ~a3294 & ~a3284;
assign a4248 = ~a4246 & ~a3056;
assign a4250 = ~a4248 & ~a4244;
assign a4252 = a4250 & a4240;
assign a4254 = a2118 & ~a1980;
assign a4256 = ~a4254 & a3056;
assign a4258 = ~a4256 & a2840;
assign a4260 = ~a4246 & ~a2118;
assign a4262 = a4260 & a3056;
assign a4264 = ~a4262 & ~a4258;
assign a4266 = a4264 & a4252;
assign a4268 = a4266 & ~a4228;
assign a4270 = a4268 & a4224;
assign a4272 = a4270 & a4212;
assign a4274 = a4272 & a4194;
assign a4276 = ~a4274 & a1100;
assign a4278 = a3232 & ~a1242;
assign a4280 = ~a4278 & ~a4276;
assign a4282 = a3302 & ~a1122;
assign a4284 = ~a4282 & a4280;
assign a4286 = a4284 & ~a1630;
assign a4288 = a4286 & ~a4148;
assign a4290 = a4288 & ~a4146;
assign a4292 = a3278 & ~a1140;
assign a4294 = a3244 & ~a1092;
assign a4296 = ~a4294 & ~a4292;
assign a4298 = a3254 & ~a1170;
assign a4300 = a3264 & ~a1232;
assign a4302 = a3318 & ~a1078;
assign a4304 = ~a4302 & ~a4300;
assign a4306 = a4304 & ~a4298;
assign a4308 = a4306 & a4296;
assign a4310 = a4308 & a4290;
assign a4312 = ~a4310 & l180;
assign a4314 = ~a4312 & a3270;
assign a4316 = a3372 & ~a1140;
assign a4318 = a2404 & ~a2266;
assign a4320 = ~a4318 & ~a3294;
assign a4322 = a4320 & ~a2544;
assign a4324 = a4322 & ~a2682;
assign a4326 = ~a4324 & ~a3222;
assign a4328 = ~a4326 & ~a1980;
assign a4330 = ~a4328 & ~a3226;
assign a4332 = ~a4330 & ~a2118;
assign a4334 = a4332 & a3056;
assign a4336 = a3342 & a1980;
assign a4338 = a4328 & a2118;
assign a4340 = ~a4338 & ~a4336;
assign a4342 = a4340 & ~a4334;
assign a4344 = a4322 & ~a3160;
assign a4346 = a4160 & a2544;
assign a4348 = a4320 & ~a3230;
assign a4350 = a4348 & ~a4346;
assign a4352 = a4350 & ~a4344;
assign a4354 = a4352 & a4342;
assign a4356 = ~a4354 & a1060;
assign a4358 = ~a4356 & ~a1698;
assign a4360 = a3368 & ~a1052;
assign a4362 = a3362 & ~a1122;
assign a4364 = ~a4362 & ~a3326;
assign a4366 = a4364 & ~a4360;
assign a4368 = a4366 & a4358;
assign a4370 = a4368 & ~a4316;
assign a4372 = ~a4370 & l180;
assign a4374 = ~a4372 & ~a3320;
assign a4376 = a3344 & ~a1092;
assign a4378 = a3348 & ~a1170;
assign a4380 = ~a4378 & ~a4376;
assign a4382 = ~a4380 & l180;
assign a4384 = ~a4382 & a3352;
assign a4386 = a3386 & ~a1232;
assign a4388 = a3392 & ~a1078;
assign a4390 = ~a4388 & ~a4386;
assign a4392 = ~a4390 & l180;
assign a4394 = ~a4392 & a3396;
assign a4396 = a4394 & a4384;
assign a4398 = a4396 & a4374;
assign a4400 = a4398 & a4314;
assign a4404 = ~a4290 & l182;
assign a4406 = ~a4404 & ~a3292;
assign a4408 = ~a4296 & l182;
assign a4410 = ~a4408 & ~a3280;
assign a4412 = ~a4306 & l182;
assign a4414 = ~a4412 & ~a3266;
assign a4416 = a4414 & a4410;
assign a4418 = a4416 & a4406;
assign a4420 = ~a4358 & l182;
assign a4422 = ~a4420 & ~a3320;
assign a4424 = ~a4366 & l182;
assign a4426 = ~a4424 & ~a3370;
assign a4428 = a4426 & a4422;
assign a4430 = a4380 & ~a4316;
assign a4432 = ~a4430 & l182;
assign a4434 = ~a4432 & ~a3374;
assign a4436 = ~a4390 & l182;
assign a4438 = ~a4436 & a3396;
assign a4440 = a4438 & a4434;
assign a4442 = a4440 & a4428;
assign a4444 = a4442 & a4418;
assign a4456 = ~a1096 & ~a1056;
assign a4458 = ~a4456 & a3308;
assign a4460 = a4458 & ~a3232;
assign a4462 = ~a4460 & l194;
assign a4464 = a3322 & a1100;
assign a4466 = a4464 & l194;
assign a4468 = a4464 & ~l194;
assign a4470 = l196 & i72;
assign a4472 = a4470 & i70;
assign a4474 = a4472 & ~l194;
assign a4476 = ~a4472 & l194;
assign a4478 = ~a4476 & ~a4474;
assign a4480 = ~a4478 & a4468;
assign a4482 = ~a4480 & ~a4466;
assign a4484 = a4482 & ~a3320;
assign a4486 = a4484 & a3270;
assign a4488 = a4486 & ~a4462;
assign a4490 = a3378 & ~a3324;
assign a4492 = ~a4490 & l194;
assign a4494 = ~a4492 & a3352;
assign a4496 = a3328 & ~l194;
assign a4498 = a4496 & ~a4478;
assign a4500 = ~a4498 & a3396;
assign a4502 = a3328 & l194;
assign a4504 = a1558 & ~a268;
assign a4506 = a4504 & l194;
assign a4508 = ~a4506 & ~a4502;
assign a4510 = a4508 & a4500;
assign a4512 = a4510 & a4494;
assign a4514 = a4512 & a4488;
assign a4518 = a4468 & ~l196;
assign a4520 = a3324 & l196;
assign a4522 = ~a4520 & ~a4466;
assign a4524 = a4522 & ~a4518;
assign a4526 = ~a3280 & ~a3246;
assign a4528 = ~a4456 & ~a3304;
assign a4530 = a4528 & ~a3232;
assign a4532 = a4530 & a4526;
assign a4534 = a4532 & ~a3292;
assign a4536 = ~a3320 & a3268;
assign a4538 = a4536 & a4534;
assign a4540 = ~a4538 & l196;
assign a4542 = ~a4540 & a4524;
assign a4544 = ~a3388 & a3380;
assign a4546 = ~a4544 & l196;
assign a4548 = a3394 & l196;
assign a4550 = a4496 & ~l196;
assign a4552 = ~a4550 & ~a4502;
assign a4554 = a4552 & ~a4548;
assign a4556 = a4504 & l196;
assign a4558 = a3322 & a1562;
assign a4560 = ~a4558 & ~a3398;
assign a4562 = a4560 & ~a4556;
assign a4564 = a4562 & a4554;
assign a4566 = a4564 & ~a4546;
assign a4568 = a4566 & a4542;
assign a4574 = l206 & i104;
assign a4576 = ~a4574 & ~l200;
assign a4578 = a4576 & ~l234;
assign a4580 = ~a3602 & i104;
assign a4582 = a4580 & l234;
assign a4584 = ~a4582 & i106;
assign a4588 = ~a3776 & ~l214;
assign a4590 = a3776 & l214;
assign a4592 = ~a4590 & ~a4588;
assign a4594 = ~a3814 & ~l216;
assign a4596 = a3814 & l216;
assign a4598 = ~a4596 & ~a4594;
assign a4600 = a4598 & a4592;
assign a4602 = ~a3662 & ~l218;
assign a4604 = a3662 & l218;
assign a4606 = ~a4604 & ~a4602;
assign a4608 = a3700 & ~l220;
assign a4610 = ~a3700 & l220;
assign a4612 = ~a4610 & ~a4608;
assign a4614 = a3734 & ~l222;
assign a4616 = ~a3734 & l222;
assign a4618 = ~a4616 & ~a4614;
assign a4620 = a4618 & a4612;
assign a4622 = a4620 & a4606;
assign a4624 = a4622 & a4600;
assign a4626 = a3848 & ~l224;
assign a4628 = ~a3848 & l224;
assign a4630 = ~a4628 & ~a4626;
assign a4632 = a3874 & ~l226;
assign a4634 = ~a3874 & l226;
assign a4636 = ~a4634 & ~a4632;
assign a4638 = a4636 & a4630;
assign a4640 = a3920 & ~l228;
assign a4642 = ~a3920 & l228;
assign a4644 = ~a4642 & ~a4640;
assign a4646 = a3942 & ~l230;
assign a4648 = ~a3942 & l230;
assign a4650 = ~a4648 & ~a4646;
assign a4652 = a3898 & ~l232;
assign a4654 = ~a3898 & l232;
assign a4656 = ~a4654 & ~a4652;
assign a4658 = a4656 & a4650;
assign a4660 = a4658 & a4644;
assign a4662 = a4660 & a4638;
assign a4664 = a4662 & a4624;
assign a4666 = a4664 & ~a3954;
assign a4668 = a4666 & ~a3616;
assign a4670 = ~a4664 & ~a3954;
assign a4672 = ~l212 & ~l210;
assign a4674 = ~a4672 & ~a4670;
assign a4676 = a4674 & ~i2;
assign a4678 = a4676 & a4668;
assign a4680 = a4678 & ~l202;
assign a4682 = a4676 & ~a4668;
assign a4684 = a4682 & l202;
assign a4686 = ~a4684 & ~a4680;
assign a4688 = l208 & l202;
assign a4690 = a4688 & a4668;
assign a4692 = a4690 & l204;
assign a4694 = ~a4690 & ~l204;
assign a4696 = ~a4694 & ~a4692;
assign a4700 = ~l208 & ~l202;
assign a4702 = ~a4700 & ~a4688;
assign a4704 = a4702 & a4678;
assign a4706 = a4682 & l208;
assign a4708 = ~a4706 & ~a4704;
assign a4710 = a3954 & ~i2;
assign a4712 = a4710 & l214;
assign a4714 = a3776 & ~i2;
assign a4716 = ~a4714 & ~a4710;
assign a4718 = ~a4716 & ~a4712;
assign a4720 = ~a3954 & ~i2;
assign a4722 = a4720 & ~a3814;
assign a4724 = a4710 & l216;
assign a4726 = ~a4724 & ~a4722;
assign a4728 = a4720 & ~a3662;
assign a4730 = a4710 & l218;
assign a4732 = ~a4730 & ~a4728;
assign a4734 = a4710 & l220;
assign a4736 = a3700 & ~i2;
assign a4738 = ~a4736 & ~a4734;
assign a4740 = a4710 & l222;
assign a4742 = a3734 & ~i2;
assign a4744 = ~a4742 & ~a4740;
assign a4746 = a4710 & l224;
assign a4748 = a3848 & ~i2;
assign a4750 = ~a4748 & ~a4746;
assign a4752 = a4710 & l226;
assign a4754 = a3874 & ~i2;
assign a4756 = ~a4754 & ~a4752;
assign a4758 = a4720 & a3920;
assign a4760 = a4710 & l228;
assign a4762 = ~a4760 & ~a4758;
assign a4764 = a4720 & a3942;
assign a4766 = a4710 & l230;
assign a4768 = ~a4766 & ~a4764;
assign a4770 = a4720 & a3898;
assign a4772 = a4710 & l232;
assign a4774 = ~a4772 & ~a4770;
assign a4776 = l124 & ~l122;
assign a4778 = ~l124 & l122;
assign a4780 = ~a4778 & ~a4776;
assign p0 = ~a4780;

assert property (~p0);

endmodule
