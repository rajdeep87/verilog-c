module m6s18 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76;

output p0;

wire na1018,na1218,na1236,na1248,na1270,na1288,na1306,na1324,na1352,na1370,na1388,na1406,na1424,na1442,na1460,
na1478,na1496,na1508,na1526,na1538,na1550,na1562,na1574,na1666,na1212,na1692,na1716,na1844,na1878,na1902,
na1914,na1932,na1950,na1968,na1986,na2004,na2016,na2038,na2166,na2182,na2194,na1660,na2188,na2208,na2176,
na2222,na2236,na2202,na2230,na2268,na2286,na2216,na2304,na2326,na2280,na2320,na2344,na2298,na2356,na2368,
na2384,na2396,na2414,na2434,na2446,na2338,na2462,na2440,na2456,na2500,na2428,na2546,na2576,na2602,na2622,
na2638,na2494,na2632,na2616,na2650,na2596,na2644,na2570,na2540,na2408,na2390,na2378,na2362,na2666,na2678,
na2696,na2714,na2732,na2350,na2726,na2708,na2690,na2672,na2746,na2660,na2740,na2262,na2758,na2774,na2786,
na2824,na2160,na2836,na2852,na2818,na2846,na2830,na2780,na2870,na2768,na2892,na2864,na2886,na2752,na2032,
na2010,na1998,na1980,na1962,na1944,na1926,na1908,na2926,na2956,na2982,na3008,na3038,na3060,na3082,na3100,
na3122,na1896,na3116,na3094,na3076,na3054,na3032,na3002,na2976,na2950,na2920,na1872,na1838,na1710,na1686,
na3134,na1568,na3146,na3128,na3158,na3140,na3170,na3152,na3182,na3164,na3194,na3176,na3208,na3188,na3220,
na3202,na3232,na3214,na3244,na3226,na3256,na3238,na3250,na1556,na1544,na1532,na1520,na1502,na1490,na1472,
na1454,na1436,na1418,na1400,na1382,na1364,na1346,na1318,na1300,na1282,na1264,na1242,a1230,na3264,na3258,
na3282,na3300,na3318,na3336,na3354,na3372,na3390,na3408,na3426,na3444,na3462,na3480,na3498,na3502,na3520,
na3526,na3532,na3538,na3550,na3638,na1012,na3650,na3674,na3786,na3820,na3844,na3856,na3874,na3892,na3910,
na3928,na3946,na3968,na4084,na4100,na4106,na4126,na3632,na4132,na4120,na4146,na4094,na4160,na4174,na4140,
na4168,na4202,na4220,na4154,na4238,na4260,na4214,na4254,na4278,na4232,na4290,na4302,na4318,na4338,na4350,
na4272,na4366,na4344,na4360,na4400,na4332,na4438,na4466,na4492,na4512,na4528,na4394,na4522,na4506,na4534,
na4486,na4460,na4432,na4312,na4296,na4550,na4556,na4574,na4592,na4610,na4284,na4604,na4586,na4568,na4624,
na4544,na4618,na4196,na4636,na4652,na4658,na4696,na4078,na4712,na4690,na4706,na4730,na4646,na4752,na4724,
na4746,na4630,na3962,na3940,na3922,na3904,na3886,na3868,na3850,na4786,na4816,na4842,na4868,na4898,na4920,
na4942,na4960,na4982,na3838,na4976,na4954,na4936,na4914,na4892,na4862,na4836,na4810,na4780,na3814,na3780,
na3668,na3644,na4994,na3544,na5006,na4988,na5018,na5000,na5030,na5012,na5042,na5024,na5054,na5036,na5066,
na5048,na5078,na5060,na5090,na5072,na5102,na5084,na5114,na5096,na5108,na3514,na3492,na3474,na3456,na3438,
na3420,na3402,na3384,na3366,na3348,na3330,na3312,na3294,a3276,na5120,c1,a822,a824,a826,a828,
a830,a832,a834,a836,a838,a840,a842,a844,a846,a848,a850,a852,a854,a856,a858,
a860,a862,a864,a866,a868,a870,a872,a874,a876,a878,a880,a882,a884,a886,a888,
a890,a892,a894,a896,a898,a900,a902,a904,a906,a908,a910,a912,a914,a916,a918,
a920,a922,a924,a926,a928,a930,a932,a934,a936,a938,a940,a942,a944,a946,a948,
a950,a952,a954,a956,a958,a960,a962,a964,a966,a968,a970,a972,a974,a976,a978,
a980,a982,a984,a986,a988,a990,a992,a994,a996,a998,a1000,a1002,a1004,a1006,a1008,
a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,a1038,
a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,a1062,a1064,a1066,a1068,
a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,a1092,a1094,a1096,a1098,
a1100,a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,a1124,a1126,a1128,
a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,a1154,a1156,a1158,
a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,a1178,a1180,a1182,a1184,a1186,a1188,
a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,a1218,
a1220,a1222,a1224,a1226,a1228,a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,a1248,a1250,
a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,a1268,a1270,a1272,a1274,a1276,a1278,a1280,
a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,a1310,
a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,a1334,a1336,a1338,a1340,
a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,a1368,a1370,
a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,a1388,a1390,a1392,a1394,a1396,a1398,a1400,
a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1426,a1428,a1430,
a1432,a1434,a1436,a1438,a1440,a1442,a1444,a1446,a1448,a1450,a1452,a1454,a1456,a1458,a1460,
a1462,a1464,a1466,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1482,a1484,a1486,a1488,a1490,
a1492,a1494,a1496,a1498,a1500,a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,a1518,a1520,
a1522,a1524,a1526,a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,a1548,a1550,
a1552,a1554,a1556,a1558,a1560,a1562,a1564,a1566,a1568,a1570,a1572,a1574,a1576,a1578,a1580,
a1582,a1584,a1586,a1588,a1590,a1592,a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,a1610,
a1612,a1614,a1616,a1618,a1620,a1622,a1624,a1626,a1628,a1630,a1632,a1634,a1636,a1638,a1640,
a1642,a1644,a1646,a1648,a1650,a1652,a1654,a1656,a1658,a1660,a1662,a1664,a1666,a1668,a1670,
a1672,a1674,a1676,a1678,a1680,a1682,a1684,a1686,a1688,a1690,a1692,a1694,a1696,a1698,a1700,
a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,
a1732,a1734,a1736,a1738,a1740,a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,a1758,a1760,
a1762,a1764,a1766,a1768,a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,a1790,
a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,
a1822,a1824,a1826,a1828,a1830,a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,a1848,a1850,
a1852,a1854,a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,
a1882,a1884,a1886,a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,a1910,
a1912,a1914,a1916,a1918,a1920,a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,a1938,a1940,
a1942,a1944,a1946,a1948,a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,
a1972,a1974,a1976,a1978,a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,a1998,a2000,
a2002,a2004,a2006,a2008,a2010,a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,a2030,
a2032,a2034,a2036,a2038,a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,a2058,a2060,
a2062,a2064,a2066,a2068,a2070,a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,a2090,
a2092,a2094,a2096,a2098,a2100,a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,a2120,
a2122,a2124,a2126,a2128,a2130,a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,
a2152,a2154,a2156,a2158,a2160,a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,a2178,a2180,
a2182,a2184,a2186,a2188,a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,a2208,a2210,
a2212,a2214,a2216,a2218,a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,a2238,a2240,
a2242,a2244,a2246,a2248,a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,a2268,a2270,
a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,a2298,a2300,
a2302,a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,a2328,a2330,
a2332,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,a2358,a2360,
a2362,a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,a2388,a2390,
a2392,a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,a2420,
a2422,a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,a2448,a2450,
a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,a2478,a2480,
a2482,a2484,a2486,a2488,a2490,a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,a2508,a2510,
a2512,a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,a2540,
a2542,a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,
a2572,a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,
a2602,a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,a2630,
a2632,a2634,a2636,a2638,a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,
a2662,a2664,a2666,a2668,a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,
a2692,a2694,a2696,a2698,a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,a2718,a2720,
a2722,a2724,a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,
a2752,a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,
a2782,a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,a2810,
a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,a2840,
a2842,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,a2870,
a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,a2900,
a2902,a2904,a2906,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2930,
a2932,a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,a2960,
a2962,a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,a2988,a2990,
a2992,a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,
a3022,a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,a3048,a3050,
a3052,a3054,a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,a3078,a3080,
a3082,a3084,a3086,a3088,a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,
a3112,a3114,a3116,a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,
a3142,a3144,a3146,a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,
a3172,a3174,a3176,a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3200,
a3202,a3204,a3206,a3208,a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,a3228,a3230,
a3232,a3234,a3236,a3238,a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,
a3262,a3264,a3266,a3268,a3270,a3272,a3274,a3278,a3280,a3282,a3284,a3286,a3288,a3290,a3292,
a3294,a3296,a3298,a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,
a3324,a3326,a3328,a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,
a3354,a3356,a3358,a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3382,
a3384,a3386,a3388,a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,a3408,a3410,a3412,
a3414,a3416,a3418,a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,a3438,a3440,a3442,
a3444,a3446,a3448,a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,a3468,a3470,a3472,
a3474,a3476,a3478,a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,a3498,a3500,a3502,
a3504,a3506,a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,a3528,a3530,a3532,
a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,a3558,a3560,a3562,
a3564,a3566,a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,a3588,a3590,a3592,
a3594,a3596,a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,a3618,a3620,a3622,
a3624,a3626,a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3648,a3650,a3652,
a3654,a3656,a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,a3678,a3680,a3682,
a3684,a3686,a3688,a3690,a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,a3712,
a3714,a3716,a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,a3738,a3740,a3742,
a3744,a3746,a3748,a3750,a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,a3768,a3770,a3772,
a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,a3798,a3800,a3802,
a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,a3828,a3830,a3832,
a3834,a3836,a3838,a3840,a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,a3858,a3860,a3862,
a3864,a3866,a3868,a3870,a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,a3888,a3890,a3892,
a3894,a3896,a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,a3918,a3920,a3922,
a3924,a3926,a3928,a3930,a3932,a3934,a3936,a3938,a3940,a3942,a3944,a3946,a3948,a3950,a3952,
a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,a3978,a3980,a3982,
a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,a4008,a4010,a4012,
a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,a4038,a4040,a4042,
a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,a4068,a4070,a4072,
a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,a4096,a4098,a4100,a4102,
a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4124,a4126,a4128,a4130,a4132,
a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,a4152,a4154,a4156,a4158,a4160,a4162,
a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,a4184,a4186,a4188,a4190,a4192,
a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,a4214,a4216,a4218,a4220,a4222,
a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,a4244,a4246,a4248,a4250,a4252,
a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,a4274,a4276,a4278,a4280,a4282,
a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,a4306,a4308,a4310,a4312,
a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,a4334,a4336,a4338,a4340,a4342,
a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,a4368,a4370,a4372,
a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,a4394,a4396,a4398,a4400,a4402,
a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,a4432,
a4434,a4436,a4438,a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,a4458,a4460,a4462,
a4464,a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4482,a4484,a4486,a4488,a4490,a4492,
a4494,a4496,a4498,a4500,a4502,a4504,a4506,a4508,a4510,a4512,a4514,a4516,a4518,a4520,a4522,
a4524,a4526,a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,
a4554,a4556,a4558,a4560,a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,a4578,a4580,a4582,
a4584,a4586,a4588,a4590,a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,a4612,
a4614,a4616,a4618,a4620,a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,a4642,
a4644,a4646,a4648,a4650,a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,a4672,
a4674,a4676,a4678,a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,a4696,a4698,a4700,a4702,
a4704,a4706,a4708,a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,a4726,a4728,a4730,a4732,
a4734,a4736,a4738,a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,a4756,a4758,a4760,a4762,
a4764,a4766,a4768,a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4784,a4786,a4788,a4790,a4792,
a4794,a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,a4818,a4820,a4822,
a4824,a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,a4844,a4846,a4848,a4850,a4852,
a4854,a4856,a4858,a4860,a4862,a4864,a4866,a4868,a4870,a4872,a4874,a4876,a4878,a4880,a4882,
a4884,a4886,a4888,a4890,a4892,a4894,a4896,a4898,a4900,a4902,a4904,a4906,a4908,a4910,a4912,
a4914,a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,a4938,a4940,a4942,
a4944,a4946,a4948,a4950,a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,a4968,a4970,a4972,
a4974,a4976,a4978,a4980,a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,a4998,a5000,a5002,
a5004,a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,a5028,a5030,a5032,
a5034,a5036,a5038,a5040,a5042,a5044,a5046,a5048,a5050,a5052,a5054,a5056,a5058,a5060,a5062,
a5064,a5066,a5068,a5070,a5072,a5074,a5076,a5078,a5080,a5082,a5084,a5086,a5088,a5090,a5092,
a5094,a5096,a5098,a5100,a5102,a5104,a5106,a5108,a5110,a5112,a5114,a5116,a5118,a5120,p0;

reg l78,l80,l82,l84,l86,l88,l90,l92,l94,l96,l98,l100,l102,l104,l106,
l108,l110,l112,l114,l116,l118,l120,l122,l124,l126,l128,l130,l132,l134,l136,
l138,l140,l142,l144,l146,l148,l150,l152,l154,l156,l158,l160,l162,l164,l166,
l168,l170,l172,l174,l176,l178,l180,l182,l184,l186,l188,l190,l192,l194,l196,
l198,l200,l202,l204,l206,l208,l210,l212,l214,l216,l218,l220,l222,l224,l226,
l228,l230,l232,l234,l236,l238,l240,l242,l244,l246,l248,l250,l252,l254,l256,
l258,l260,l262,l264,l266,l268,l270,l272,l274,l276,l278,l280,l282,l284,l286,
l288,l290,l292,l294,l296,l298,l300,l302,l304,l306,l308,l310,l312,l314,l316,
l318,l320,l322,l324,l326,l328,l330,l332,l334,l336,l338,l340,l342,l344,l346,
l348,l350,l352,l354,l356,l358,l360,l362,l364,l366,l368,l370,l372,l374,l376,
l378,l380,l382,l384,l386,l388,l390,l392,l394,l396,l398,l400,l402,l404,l406,
l408,l410,l412,l414,l416,l418,l420,l422,l424,l426,l428,l430,l432,l434,l436,
l438,l440,l442,l444,l446,l448,l450,l452,l454,l456,l458,l460,l462,l464,l466,
l468,l470,l472,l474,l476,l478,l480,l482,l484,l486,l488,l490,l492,l494,l496,
l498,l500,l502,l504,l506,l508,l510,l512,l514,l516,l518,l520,l522,l524,l526,
l528,l530,l532,l534,l536,l538,l540,l542,l544,l546,l548,l550,l552,l554,l556,
l558,l560,l562,l564,l566,l568,l570,l572,l574,l576,l578,l580,l582,l584,l586,
l588,l590,l592,l594,l596,l598,l600,l602,l604,l606,l608,l610,l612,l614,l616,
l618,l620,l622,l624,l626,l628,l630,l632,l634,l636,l638,l640,l642,l644,l646,
l648,l650,l652,l654,l656,l658,l660,l662,l664,l666,l668,l670,l672,l674,l676,
l678,l680,l682,l684,l686,l688,l690,l692,l694,l696,l698,l700,l702,l704,l706,
l708,l710,l712,l714,l716,l718,l720,l722,l724,l726,l728,l730,l732,l734,l736,
l738,l740,l742,l744,l746,l748,l750,l752,l754,l756,l758,l760,l762,l764,l766,
l768,l770,l772,l774,l776,l778,l780,l782,l784,l786,l788,l790,l792,l794,l796,
l798,l800,l802,l804,l806,l808,l810,l812,l814,l816,l818,l820;

initial
begin
   l78 = 0;
   l80 = 0;
   l82 = 0;
   l84 = 0;
   l86 = 0;
   l88 = 0;
   l90 = 0;
   l92 = 0;
   l94 = 0;
   l96 = 0;
   l98 = 0;
   l100 = 0;
   l102 = 0;
   l104 = 0;
   l106 = 0;
   l108 = 0;
   l110 = 0;
   l112 = 0;
   l114 = 0;
   l116 = 0;
   l118 = 0;
   l120 = 0;
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
   l392 = 0;
   l394 = 0;
   l396 = 0;
   l398 = 0;
   l400 = 0;
   l402 = 0;
   l404 = 0;
   l406 = 0;
   l408 = 0;
   l410 = 0;
   l412 = 0;
   l414 = 0;
   l416 = 0;
   l418 = 0;
   l420 = 0;
   l422 = 0;
   l424 = 0;
   l426 = 0;
   l428 = 0;
   l430 = 0;
   l432 = 0;
   l434 = 0;
   l436 = 0;
   l438 = 0;
   l440 = 0;
   l442 = 0;
   l444 = 0;
   l446 = 0;
   l448 = 0;
   l450 = 0;
   l452 = 0;
   l454 = 0;
   l456 = 0;
   l458 = 0;
   l460 = 0;
   l462 = 0;
   l464 = 0;
   l466 = 0;
   l468 = 0;
   l470 = 0;
   l472 = 0;
   l474 = 0;
   l476 = 0;
   l478 = 0;
   l480 = 0;
   l482 = 0;
   l484 = 0;
   l486 = 0;
   l488 = 0;
   l490 = 0;
   l492 = 0;
   l494 = 0;
   l496 = 0;
   l498 = 0;
   l500 = 0;
   l502 = 0;
   l504 = 0;
   l506 = 0;
   l508 = 0;
   l510 = 0;
   l512 = 0;
   l514 = 0;
   l516 = 0;
   l518 = 0;
   l520 = 0;
   l522 = 0;
   l524 = 0;
   l526 = 0;
   l528 = 0;
   l530 = 0;
   l532 = 0;
   l534 = 0;
   l536 = 0;
   l538 = 0;
   l540 = 0;
   l542 = 0;
   l544 = 0;
   l546 = 0;
   l548 = 0;
   l550 = 0;
   l552 = 0;
   l554 = 0;
   l556 = 0;
   l558 = 0;
   l560 = 0;
   l562 = 0;
   l564 = 0;
   l566 = 0;
   l568 = 0;
   l570 = 0;
   l572 = 0;
   l574 = 0;
   l576 = 0;
   l578 = 0;
   l580 = 0;
   l582 = 0;
   l584 = 0;
   l586 = 0;
   l588 = 0;
   l590 = 0;
   l592 = 0;
   l594 = 0;
   l596 = 0;
   l598 = 0;
   l600 = 0;
   l602 = 0;
   l604 = 0;
   l606 = 0;
   l608 = 0;
   l610 = 0;
   l612 = 0;
   l614 = 0;
   l616 = 0;
   l618 = 0;
   l620 = 0;
   l622 = 0;
   l624 = 0;
   l626 = 0;
   l628 = 0;
   l630 = 0;
   l632 = 0;
   l634 = 0;
   l636 = 0;
   l638 = 0;
   l640 = 0;
   l642 = 0;
   l644 = 0;
   l646 = 0;
   l648 = 0;
   l650 = 0;
   l652 = 0;
   l654 = 0;
   l656 = 0;
   l658 = 0;
   l660 = 0;
   l662 = 0;
   l664 = 0;
   l666 = 0;
   l668 = 0;
   l670 = 0;
   l672 = 0;
   l674 = 0;
   l676 = 0;
   l678 = 0;
   l680 = 0;
   l682 = 0;
   l684 = 0;
   l686 = 0;
   l688 = 0;
   l690 = 0;
   l692 = 0;
   l694 = 0;
   l696 = 0;
   l698 = 0;
   l700 = 0;
   l702 = 0;
   l704 = 0;
   l706 = 0;
   l708 = 0;
   l710 = 0;
   l712 = 0;
   l714 = 0;
   l716 = 0;
   l718 = 0;
   l720 = 0;
   l722 = 0;
   l724 = 0;
   l726 = 0;
   l728 = 0;
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
   l802 = 0;
   l804 = 0;
   l806 = 0;
   l808 = 0;
   l810 = 0;
   l812 = 0;
   l814 = 0;
   l816 = 0;
   l818 = 0;
   l820 = 0;
end

always @(posedge na1018)
   l78 <= na1018;

always @(posedge na1218)
   l80 <= na1218;

always @(posedge na1236)
   l82 <= na1236;

always @(posedge na1248)
   l84 <= na1248;

always @(posedge i2)
   l86 <= i2;

always @(posedge na1270)
   l88 <= na1270;

always @(posedge na1288)
   l90 <= na1288;

always @(posedge na1306)
   l92 <= na1306;

always @(posedge na1324)
   l94 <= na1324;

always @(posedge na1352)
   l96 <= na1352;

always @(posedge na1370)
   l98 <= na1370;

always @(posedge na1388)
   l100 <= na1388;

always @(posedge na1406)
   l102 <= na1406;

always @(posedge na1424)
   l104 <= na1424;

always @(posedge na1442)
   l106 <= na1442;

always @(posedge na1460)
   l108 <= na1460;

always @(posedge na1478)
   l110 <= na1478;

always @(posedge na1496)
   l112 <= na1496;

always @(posedge na1508)
   l114 <= na1508;

always @(posedge na1526)
   l116 <= na1526;

always @(posedge na1538)
   l118 <= na1538;

always @(posedge na1550)
   l120 <= na1550;

always @(posedge na1562)
   l122 <= na1562;

always @(posedge na1574)
   l124 <= na1574;

always @(posedge na1666)
   l126 <= na1666;

always @(posedge na1212)
   l128 <= na1212;

always @(posedge na1692)
   l130 <= na1692;

always @(posedge na1716)
   l132 <= na1716;

always @(posedge na1844)
   l134 <= na1844;

always @(posedge na1878)
   l136 <= na1878;

always @(posedge na1902)
   l138 <= na1902;

always @(posedge na1914)
   l140 <= na1914;

always @(posedge na1932)
   l142 <= na1932;

always @(posedge na1950)
   l144 <= na1950;

always @(posedge na1968)
   l146 <= na1968;

always @(posedge na1986)
   l148 <= na1986;

always @(posedge na2004)
   l150 <= na2004;

always @(posedge na2016)
   l152 <= na2016;

always @(posedge na2038)
   l154 <= na2038;

always @(posedge na2166)
   l156 <= na2166;

always @(posedge na2182)
   l158 <= na2182;

always @(posedge na2194)
   l160 <= na2194;

always @(posedge na1660)
   l162 <= na1660;

always @(posedge na2188)
   l164 <= na2188;

always @(posedge na2208)
   l166 <= na2208;

always @(posedge na2176)
   l168 <= na2176;

always @(posedge na2222)
   l170 <= na2222;

always @(posedge na2236)
   l172 <= na2236;

always @(posedge na2202)
   l174 <= na2202;

always @(posedge na2230)
   l176 <= na2230;

always @(posedge na2268)
   l178 <= na2268;

always @(posedge na2286)
   l180 <= na2286;

always @(posedge na2216)
   l182 <= na2216;

always @(posedge na2304)
   l184 <= na2304;

always @(posedge na2326)
   l186 <= na2326;

always @(posedge na2280)
   l188 <= na2280;

always @(posedge na2320)
   l190 <= na2320;

always @(posedge na2344)
   l192 <= na2344;

always @(posedge na2298)
   l194 <= na2298;

always @(posedge na2356)
   l196 <= na2356;

always @(posedge na2368)
   l198 <= na2368;

always @(posedge na2384)
   l200 <= na2384;

always @(posedge na2396)
   l202 <= na2396;

always @(posedge na2414)
   l204 <= na2414;

always @(posedge na2434)
   l206 <= na2434;

always @(posedge na2446)
   l208 <= na2446;

always @(posedge na2338)
   l210 <= na2338;

always @(posedge na2462)
   l212 <= na2462;

always @(posedge na2440)
   l214 <= na2440;

always @(posedge na2456)
   l216 <= na2456;

always @(posedge na2500)
   l218 <= na2500;

always @(posedge na2428)
   l220 <= na2428;

always @(posedge na2546)
   l222 <= na2546;

always @(posedge na2576)
   l224 <= na2576;

always @(posedge na2602)
   l226 <= na2602;

always @(posedge na2622)
   l228 <= na2622;

always @(posedge na2638)
   l230 <= na2638;

always @(posedge na2494)
   l232 <= na2494;

always @(posedge na2632)
   l234 <= na2632;

always @(posedge na2616)
   l236 <= na2616;

always @(posedge na2650)
   l238 <= na2650;

always @(posedge na2596)
   l240 <= na2596;

always @(posedge na2644)
   l242 <= na2644;

always @(posedge na2570)
   l244 <= na2570;

always @(posedge na2540)
   l246 <= na2540;

always @(posedge na2408)
   l248 <= na2408;

always @(posedge na2390)
   l250 <= na2390;

always @(posedge na2378)
   l252 <= na2378;

always @(posedge na2362)
   l254 <= na2362;

always @(posedge na2666)
   l256 <= na2666;

always @(posedge na2678)
   l258 <= na2678;

always @(posedge na2696)
   l260 <= na2696;

always @(posedge na2714)
   l262 <= na2714;

always @(posedge na2732)
   l264 <= na2732;

always @(posedge na2350)
   l266 <= na2350;

always @(posedge na2726)
   l268 <= na2726;

always @(posedge na2708)
   l270 <= na2708;

always @(posedge na2690)
   l272 <= na2690;

always @(posedge na2672)
   l274 <= na2672;

always @(posedge na2746)
   l276 <= na2746;

always @(posedge na2660)
   l278 <= na2660;

always @(posedge na2740)
   l280 <= na2740;

always @(posedge na2262)
   l282 <= na2262;

always @(posedge na2758)
   l284 <= na2758;

always @(posedge na2774)
   l286 <= na2774;

always @(posedge na2786)
   l288 <= na2786;

always @(posedge na2824)
   l290 <= na2824;

always @(posedge na2160)
   l292 <= na2160;

always @(posedge na2836)
   l294 <= na2836;

always @(posedge na2852)
   l296 <= na2852;

always @(posedge na2818)
   l298 <= na2818;

always @(posedge na2846)
   l300 <= na2846;

always @(posedge na2830)
   l302 <= na2830;

always @(posedge na2780)
   l304 <= na2780;

always @(posedge na2870)
   l306 <= na2870;

always @(posedge na2768)
   l308 <= na2768;

always @(posedge na2892)
   l310 <= na2892;

always @(posedge na2864)
   l312 <= na2864;

always @(posedge na2886)
   l314 <= na2886;

always @(posedge na2752)
   l316 <= na2752;

always @(posedge na2032)
   l318 <= na2032;

always @(posedge na2010)
   l320 <= na2010;

always @(posedge na1998)
   l322 <= na1998;

always @(posedge na1980)
   l324 <= na1980;

always @(posedge na1962)
   l326 <= na1962;

always @(posedge na1944)
   l328 <= na1944;

always @(posedge na1926)
   l330 <= na1926;

always @(posedge na1908)
   l332 <= na1908;

always @(posedge na2926)
   l334 <= na2926;

always @(posedge na2956)
   l336 <= na2956;

always @(posedge na2982)
   l338 <= na2982;

always @(posedge na3008)
   l340 <= na3008;

always @(posedge na3038)
   l342 <= na3038;

always @(posedge na3060)
   l344 <= na3060;

always @(posedge na3082)
   l346 <= na3082;

always @(posedge na3100)
   l348 <= na3100;

always @(posedge na3122)
   l350 <= na3122;

always @(posedge na1896)
   l352 <= na1896;

always @(posedge na3116)
   l354 <= na3116;

always @(posedge na3094)
   l356 <= na3094;

always @(posedge na3076)
   l358 <= na3076;

always @(posedge na3054)
   l360 <= na3054;

always @(posedge na3032)
   l362 <= na3032;

always @(posedge na3002)
   l364 <= na3002;

always @(posedge na2976)
   l366 <= na2976;

always @(posedge na2950)
   l368 <= na2950;

always @(posedge na2920)
   l370 <= na2920;

always @(posedge na1872)
   l372 <= na1872;

always @(posedge na1838)
   l374 <= na1838;

always @(posedge na1710)
   l376 <= na1710;

always @(posedge na1686)
   l378 <= na1686;

always @(posedge na3134)
   l380 <= na3134;

always @(posedge na1568)
   l382 <= na1568;

always @(posedge na3146)
   l384 <= na3146;

always @(posedge na3128)
   l386 <= na3128;

always @(posedge na3158)
   l388 <= na3158;

always @(posedge na3140)
   l390 <= na3140;

always @(posedge na3170)
   l392 <= na3170;

always @(posedge na3152)
   l394 <= na3152;

always @(posedge na3182)
   l396 <= na3182;

always @(posedge na3164)
   l398 <= na3164;

always @(posedge na3194)
   l400 <= na3194;

always @(posedge na3176)
   l402 <= na3176;

always @(posedge na3208)
   l404 <= na3208;

always @(posedge na3188)
   l406 <= na3188;

always @(posedge na3220)
   l408 <= na3220;

always @(posedge na3202)
   l410 <= na3202;

always @(posedge na3232)
   l412 <= na3232;

always @(posedge na3214)
   l414 <= na3214;

always @(posedge na3244)
   l416 <= na3244;

always @(posedge na3226)
   l418 <= na3226;

always @(posedge na3256)
   l420 <= na3256;

always @(posedge na3238)
   l422 <= na3238;

always @(posedge na3250)
   l424 <= na3250;

always @(posedge na1556)
   l426 <= na1556;

always @(posedge na1544)
   l428 <= na1544;

always @(posedge na1532)
   l430 <= na1532;

always @(posedge na1520)
   l432 <= na1520;

always @(posedge na1502)
   l434 <= na1502;

always @(posedge na1490)
   l436 <= na1490;

always @(posedge na1472)
   l438 <= na1472;

always @(posedge na1454)
   l440 <= na1454;

always @(posedge na1436)
   l442 <= na1436;

always @(posedge na1418)
   l444 <= na1418;

always @(posedge na1400)
   l446 <= na1400;

always @(posedge na1382)
   l448 <= na1382;

always @(posedge na1364)
   l450 <= na1364;

always @(posedge na1346)
   l452 <= na1346;

always @(posedge na1318)
   l454 <= na1318;

always @(posedge na1300)
   l456 <= na1300;

always @(posedge na1282)
   l458 <= na1282;

always @(posedge na1264)
   l460 <= na1264;

always @(posedge na1242)
   l462 <= na1242;

always @(posedge a1230)
   l464 <= a1230;

always @(posedge na3264)
   l466 <= na3264;

always @(posedge na3258)
   l468 <= na3258;

always @(posedge na3282)
   l470 <= na3282;

always @(posedge na3300)
   l472 <= na3300;

always @(posedge na3318)
   l474 <= na3318;

always @(posedge na3336)
   l476 <= na3336;

always @(posedge na3354)
   l478 <= na3354;

always @(posedge na3372)
   l480 <= na3372;

always @(posedge na3390)
   l482 <= na3390;

always @(posedge na3408)
   l484 <= na3408;

always @(posedge na3426)
   l486 <= na3426;

always @(posedge na3444)
   l488 <= na3444;

always @(posedge na3462)
   l490 <= na3462;

always @(posedge na3480)
   l492 <= na3480;

always @(posedge na3498)
   l494 <= na3498;

always @(posedge na3502)
   l496 <= na3502;

always @(posedge na3520)
   l498 <= na3520;

always @(posedge na3526)
   l500 <= na3526;

always @(posedge na3532)
   l502 <= na3532;

always @(posedge na3538)
   l504 <= na3538;

always @(posedge na3550)
   l506 <= na3550;

always @(posedge na3638)
   l508 <= na3638;

always @(posedge na1012)
   l510 <= na1012;

always @(posedge na3650)
   l512 <= na3650;

always @(posedge na3674)
   l514 <= na3674;

always @(posedge na3786)
   l516 <= na3786;

always @(posedge na3820)
   l518 <= na3820;

always @(posedge na3844)
   l520 <= na3844;

always @(posedge na3856)
   l522 <= na3856;

always @(posedge na3874)
   l524 <= na3874;

always @(posedge na3892)
   l526 <= na3892;

always @(posedge na3910)
   l528 <= na3910;

always @(posedge na3928)
   l530 <= na3928;

always @(posedge na3946)
   l532 <= na3946;

always @(posedge na3968)
   l534 <= na3968;

always @(posedge na4084)
   l536 <= na4084;

always @(posedge na4100)
   l538 <= na4100;

always @(posedge na4106)
   l540 <= na4106;

always @(posedge na4126)
   l542 <= na4126;

always @(posedge na3632)
   l544 <= na3632;

always @(posedge na4132)
   l546 <= na4132;

always @(posedge na4120)
   l548 <= na4120;

always @(posedge na4146)
   l550 <= na4146;

always @(posedge na4094)
   l552 <= na4094;

always @(posedge na4160)
   l554 <= na4160;

always @(posedge na4174)
   l556 <= na4174;

always @(posedge na4140)
   l558 <= na4140;

always @(posedge na4168)
   l560 <= na4168;

always @(posedge na4202)
   l562 <= na4202;

always @(posedge na4220)
   l564 <= na4220;

always @(posedge na4154)
   l566 <= na4154;

always @(posedge na4238)
   l568 <= na4238;

always @(posedge na4260)
   l570 <= na4260;

always @(posedge na4214)
   l572 <= na4214;

always @(posedge na4254)
   l574 <= na4254;

always @(posedge na4278)
   l576 <= na4278;

always @(posedge na4232)
   l578 <= na4232;

always @(posedge na4290)
   l580 <= na4290;

always @(posedge na4302)
   l582 <= na4302;

always @(posedge na4318)
   l584 <= na4318;

always @(posedge na4338)
   l586 <= na4338;

always @(posedge na4350)
   l588 <= na4350;

always @(posedge na4272)
   l590 <= na4272;

always @(posedge na4366)
   l592 <= na4366;

always @(posedge na4344)
   l594 <= na4344;

always @(posedge na4360)
   l596 <= na4360;

always @(posedge na4400)
   l598 <= na4400;

always @(posedge na4332)
   l600 <= na4332;

always @(posedge na4438)
   l602 <= na4438;

always @(posedge na4466)
   l604 <= na4466;

always @(posedge na4492)
   l606 <= na4492;

always @(posedge na4512)
   l608 <= na4512;

always @(posedge na4528)
   l610 <= na4528;

always @(posedge na4394)
   l612 <= na4394;

always @(posedge na4522)
   l614 <= na4522;

always @(posedge na4506)
   l616 <= na4506;

always @(posedge na4534)
   l618 <= na4534;

always @(posedge na4486)
   l620 <= na4486;

always @(posedge na4460)
   l622 <= na4460;

always @(posedge na4432)
   l624 <= na4432;

always @(posedge na4312)
   l626 <= na4312;

always @(posedge na4296)
   l628 <= na4296;

always @(posedge na4550)
   l630 <= na4550;

always @(posedge na4556)
   l632 <= na4556;

always @(posedge na4574)
   l634 <= na4574;

always @(posedge na4592)
   l636 <= na4592;

always @(posedge na4610)
   l638 <= na4610;

always @(posedge na4284)
   l640 <= na4284;

always @(posedge na4604)
   l642 <= na4604;

always @(posedge na4586)
   l644 <= na4586;

always @(posedge na4568)
   l646 <= na4568;

always @(posedge na4624)
   l648 <= na4624;

always @(posedge na4544)
   l650 <= na4544;

always @(posedge na4618)
   l652 <= na4618;

always @(posedge na4196)
   l654 <= na4196;

always @(posedge na4636)
   l656 <= na4636;

always @(posedge na4652)
   l658 <= na4652;

always @(posedge na4658)
   l660 <= na4658;

always @(posedge na4696)
   l662 <= na4696;

always @(posedge na4078)
   l664 <= na4078;

always @(posedge na4712)
   l666 <= na4712;

always @(posedge na4690)
   l668 <= na4690;

always @(posedge na4706)
   l670 <= na4706;

always @(posedge na4730)
   l672 <= na4730;

always @(posedge na4646)
   l674 <= na4646;

always @(posedge na4752)
   l676 <= na4752;

always @(posedge na4724)
   l678 <= na4724;

always @(posedge na4746)
   l680 <= na4746;

always @(posedge na4630)
   l682 <= na4630;

always @(posedge na3962)
   l684 <= na3962;

always @(posedge na3940)
   l686 <= na3940;

always @(posedge na3922)
   l688 <= na3922;

always @(posedge na3904)
   l690 <= na3904;

always @(posedge na3886)
   l692 <= na3886;

always @(posedge na3868)
   l694 <= na3868;

always @(posedge na3850)
   l696 <= na3850;

always @(posedge na4786)
   l698 <= na4786;

always @(posedge na4816)
   l700 <= na4816;

always @(posedge na4842)
   l702 <= na4842;

always @(posedge na4868)
   l704 <= na4868;

always @(posedge na4898)
   l706 <= na4898;

always @(posedge na4920)
   l708 <= na4920;

always @(posedge na4942)
   l710 <= na4942;

always @(posedge na4960)
   l712 <= na4960;

always @(posedge na4982)
   l714 <= na4982;

always @(posedge na3838)
   l716 <= na3838;

always @(posedge na4976)
   l718 <= na4976;

always @(posedge na4954)
   l720 <= na4954;

always @(posedge na4936)
   l722 <= na4936;

always @(posedge na4914)
   l724 <= na4914;

always @(posedge na4892)
   l726 <= na4892;

always @(posedge na4862)
   l728 <= na4862;

always @(posedge na4836)
   l730 <= na4836;

always @(posedge na4810)
   l732 <= na4810;

always @(posedge na4780)
   l734 <= na4780;

always @(posedge na3814)
   l736 <= na3814;

always @(posedge na3780)
   l738 <= na3780;

always @(posedge na3668)
   l740 <= na3668;

always @(posedge na3644)
   l742 <= na3644;

always @(posedge na4994)
   l744 <= na4994;

always @(posedge na3544)
   l746 <= na3544;

always @(posedge na5006)
   l748 <= na5006;

always @(posedge na4988)
   l750 <= na4988;

always @(posedge na5018)
   l752 <= na5018;

always @(posedge na5000)
   l754 <= na5000;

always @(posedge na5030)
   l756 <= na5030;

always @(posedge na5012)
   l758 <= na5012;

always @(posedge na5042)
   l760 <= na5042;

always @(posedge na5024)
   l762 <= na5024;

always @(posedge na5054)
   l764 <= na5054;

always @(posedge na5036)
   l766 <= na5036;

always @(posedge na5066)
   l768 <= na5066;

always @(posedge na5048)
   l770 <= na5048;

always @(posedge na5078)
   l772 <= na5078;

always @(posedge na5060)
   l774 <= na5060;

always @(posedge na5090)
   l776 <= na5090;

always @(posedge na5072)
   l778 <= na5072;

always @(posedge na5102)
   l780 <= na5102;

always @(posedge na5084)
   l782 <= na5084;

always @(posedge na5114)
   l784 <= na5114;

always @(posedge na5096)
   l786 <= na5096;

always @(posedge na5108)
   l788 <= na5108;

always @(posedge na3514)
   l790 <= na3514;

always @(posedge na3492)
   l792 <= na3492;

always @(posedge na3474)
   l794 <= na3474;

always @(posedge na3456)
   l796 <= na3456;

always @(posedge na3438)
   l798 <= na3438;

always @(posedge na3420)
   l800 <= na3420;

always @(posedge na3402)
   l802 <= na3402;

always @(posedge na3384)
   l804 <= na3384;

always @(posedge na3366)
   l806 <= na3366;

always @(posedge na3348)
   l808 <= na3348;

always @(posedge na3330)
   l810 <= na3330;

always @(posedge na3312)
   l812 <= na3312;

always @(posedge na3294)
   l814 <= na3294;

always @(posedge a3276)
   l816 <= a3276;

always @(posedge na5120)
   l818 <= na5120;

always @(posedge c1)
   l820 <= c1;


assign na1018 = ~a1018;
assign na1218 = ~a1218;
assign na1236 = ~a1236;
assign na1248 = ~a1248;
assign na1270 = ~a1270;
assign na1288 = ~a1288;
assign na1306 = ~a1306;
assign na1324 = ~a1324;
assign na1352 = ~a1352;
assign na1370 = ~a1370;
assign na1388 = ~a1388;
assign na1406 = ~a1406;
assign na1424 = ~a1424;
assign na1442 = ~a1442;
assign na1460 = ~a1460;
assign na1478 = ~a1478;
assign na1496 = ~a1496;
assign na1508 = ~a1508;
assign na1526 = ~a1526;
assign na1538 = ~a1538;
assign na1550 = ~a1550;
assign na1562 = ~a1562;
assign na1574 = ~a1574;
assign na1666 = ~a1666;
assign na1212 = ~a1212;
assign na1692 = ~a1692;
assign na1716 = ~a1716;
assign na1844 = ~a1844;
assign na1878 = ~a1878;
assign na1902 = ~a1902;
assign na1914 = ~a1914;
assign na1932 = ~a1932;
assign na1950 = ~a1950;
assign na1968 = ~a1968;
assign na1986 = ~a1986;
assign na2004 = ~a2004;
assign na2016 = ~a2016;
assign na2038 = ~a2038;
assign na2166 = ~a2166;
assign na2182 = ~a2182;
assign na2194 = ~a2194;
assign na1660 = ~a1660;
assign na2188 = ~a2188;
assign na2208 = ~a2208;
assign na2176 = ~a2176;
assign na2222 = ~a2222;
assign na2236 = ~a2236;
assign na2202 = ~a2202;
assign na2230 = ~a2230;
assign na2268 = ~a2268;
assign na2286 = ~a2286;
assign na2216 = ~a2216;
assign na2304 = ~a2304;
assign na2326 = ~a2326;
assign na2280 = ~a2280;
assign na2320 = ~a2320;
assign na2344 = ~a2344;
assign na2298 = ~a2298;
assign na2356 = ~a2356;
assign na2368 = ~a2368;
assign na2384 = ~a2384;
assign na2396 = ~a2396;
assign na2414 = ~a2414;
assign na2434 = ~a2434;
assign na2446 = ~a2446;
assign na2338 = ~a2338;
assign na2462 = ~a2462;
assign na2440 = ~a2440;
assign na2456 = ~a2456;
assign na2500 = ~a2500;
assign na2428 = ~a2428;
assign na2546 = ~a2546;
assign na2576 = ~a2576;
assign na2602 = ~a2602;
assign na2622 = ~a2622;
assign na2638 = ~a2638;
assign na2494 = ~a2494;
assign na2632 = ~a2632;
assign na2616 = ~a2616;
assign na2650 = ~a2650;
assign na2596 = ~a2596;
assign na2644 = ~a2644;
assign na2570 = ~a2570;
assign na2540 = ~a2540;
assign na2408 = ~a2408;
assign na2390 = ~a2390;
assign na2378 = ~a2378;
assign na2362 = ~a2362;
assign na2666 = ~a2666;
assign na2678 = ~a2678;
assign na2696 = ~a2696;
assign na2714 = ~a2714;
assign na2732 = ~a2732;
assign na2350 = ~a2350;
assign na2726 = ~a2726;
assign na2708 = ~a2708;
assign na2690 = ~a2690;
assign na2672 = ~a2672;
assign na2746 = ~a2746;
assign na2660 = ~a2660;
assign na2740 = ~a2740;
assign na2262 = ~a2262;
assign na2758 = ~a2758;
assign na2774 = ~a2774;
assign na2786 = ~a2786;
assign na2824 = ~a2824;
assign na2160 = ~a2160;
assign na2836 = ~a2836;
assign na2852 = ~a2852;
assign na2818 = ~a2818;
assign na2846 = ~a2846;
assign na2830 = ~a2830;
assign na2780 = ~a2780;
assign na2870 = ~a2870;
assign na2768 = ~a2768;
assign na2892 = ~a2892;
assign na2864 = ~a2864;
assign na2886 = ~a2886;
assign na2752 = ~a2752;
assign na2032 = ~a2032;
assign na2010 = ~a2010;
assign na1998 = ~a1998;
assign na1980 = ~a1980;
assign na1962 = ~a1962;
assign na1944 = ~a1944;
assign na1926 = ~a1926;
assign na1908 = ~a1908;
assign na2926 = ~a2926;
assign na2956 = ~a2956;
assign na2982 = ~a2982;
assign na3008 = ~a3008;
assign na3038 = ~a3038;
assign na3060 = ~a3060;
assign na3082 = ~a3082;
assign na3100 = ~a3100;
assign na3122 = ~a3122;
assign na1896 = ~a1896;
assign na3116 = ~a3116;
assign na3094 = ~a3094;
assign na3076 = ~a3076;
assign na3054 = ~a3054;
assign na3032 = ~a3032;
assign na3002 = ~a3002;
assign na2976 = ~a2976;
assign na2950 = ~a2950;
assign na2920 = ~a2920;
assign na1872 = ~a1872;
assign na1838 = ~a1838;
assign na1710 = ~a1710;
assign na1686 = ~a1686;
assign na3134 = ~a3134;
assign na1568 = ~a1568;
assign na3146 = ~a3146;
assign na3128 = ~a3128;
assign na3158 = ~a3158;
assign na3140 = ~a3140;
assign na3170 = ~a3170;
assign na3152 = ~a3152;
assign na3182 = ~a3182;
assign na3164 = ~a3164;
assign na3194 = ~a3194;
assign na3176 = ~a3176;
assign na3208 = ~a3208;
assign na3188 = ~a3188;
assign na3220 = ~a3220;
assign na3202 = ~a3202;
assign na3232 = ~a3232;
assign na3214 = ~a3214;
assign na3244 = ~a3244;
assign na3226 = ~a3226;
assign na3256 = ~a3256;
assign na3238 = ~a3238;
assign na3250 = ~a3250;
assign na1556 = ~a1556;
assign na1544 = ~a1544;
assign na1532 = ~a1532;
assign na1520 = ~a1520;
assign na1502 = ~a1502;
assign na1490 = ~a1490;
assign na1472 = ~a1472;
assign na1454 = ~a1454;
assign na1436 = ~a1436;
assign na1418 = ~a1418;
assign na1400 = ~a1400;
assign na1382 = ~a1382;
assign na1364 = ~a1364;
assign na1346 = ~a1346;
assign na1318 = ~a1318;
assign na1300 = ~a1300;
assign na1282 = ~a1282;
assign na1264 = ~a1264;
assign na1242 = ~a1242;
assign a1230 = ~a1228 & ~a1220;
assign na3264 = ~a3264;
assign na3258 = ~a3258;
assign na3282 = ~a3282;
assign na3300 = ~a3300;
assign na3318 = ~a3318;
assign na3336 = ~a3336;
assign na3354 = ~a3354;
assign na3372 = ~a3372;
assign na3390 = ~a3390;
assign na3408 = ~a3408;
assign na3426 = ~a3426;
assign na3444 = ~a3444;
assign na3462 = ~a3462;
assign na3480 = ~a3480;
assign na3498 = ~a3498;
assign na3502 = ~a3502;
assign na3520 = ~a3520;
assign na3526 = ~a3526;
assign na3532 = ~a3532;
assign na3538 = ~a3538;
assign na3550 = ~a3550;
assign na3638 = ~a3638;
assign na1012 = ~a1012;
assign na3650 = ~a3650;
assign na3674 = ~a3674;
assign na3786 = ~a3786;
assign na3820 = ~a3820;
assign na3844 = ~a3844;
assign na3856 = ~a3856;
assign na3874 = ~a3874;
assign na3892 = ~a3892;
assign na3910 = ~a3910;
assign na3928 = ~a3928;
assign na3946 = ~a3946;
assign na3968 = ~a3968;
assign na4084 = ~a4084;
assign na4100 = ~a4100;
assign na4106 = ~a4106;
assign na4126 = ~a4126;
assign na3632 = ~a3632;
assign na4132 = ~a4132;
assign na4120 = ~a4120;
assign na4146 = ~a4146;
assign na4094 = ~a4094;
assign na4160 = ~a4160;
assign na4174 = ~a4174;
assign na4140 = ~a4140;
assign na4168 = ~a4168;
assign na4202 = ~a4202;
assign na4220 = ~a4220;
assign na4154 = ~a4154;
assign na4238 = ~a4238;
assign na4260 = ~a4260;
assign na4214 = ~a4214;
assign na4254 = ~a4254;
assign na4278 = ~a4278;
assign na4232 = ~a4232;
assign na4290 = ~a4290;
assign na4302 = ~a4302;
assign na4318 = ~a4318;
assign na4338 = ~a4338;
assign na4350 = ~a4350;
assign na4272 = ~a4272;
assign na4366 = ~a4366;
assign na4344 = ~a4344;
assign na4360 = ~a4360;
assign na4400 = ~a4400;
assign na4332 = ~a4332;
assign na4438 = ~a4438;
assign na4466 = ~a4466;
assign na4492 = ~a4492;
assign na4512 = ~a4512;
assign na4528 = ~a4528;
assign na4394 = ~a4394;
assign na4522 = ~a4522;
assign na4506 = ~a4506;
assign na4534 = ~a4534;
assign na4486 = ~a4486;
assign na4460 = ~a4460;
assign na4432 = ~a4432;
assign na4312 = ~a4312;
assign na4296 = ~a4296;
assign na4550 = ~a4550;
assign na4556 = ~a4556;
assign na4574 = ~a4574;
assign na4592 = ~a4592;
assign na4610 = ~a4610;
assign na4284 = ~a4284;
assign na4604 = ~a4604;
assign na4586 = ~a4586;
assign na4568 = ~a4568;
assign na4624 = ~a4624;
assign na4544 = ~a4544;
assign na4618 = ~a4618;
assign na4196 = ~a4196;
assign na4636 = ~a4636;
assign na4652 = ~a4652;
assign na4658 = ~a4658;
assign na4696 = ~a4696;
assign na4078 = ~a4078;
assign na4712 = ~a4712;
assign na4690 = ~a4690;
assign na4706 = ~a4706;
assign na4730 = ~a4730;
assign na4646 = ~a4646;
assign na4752 = ~a4752;
assign na4724 = ~a4724;
assign na4746 = ~a4746;
assign na4630 = ~a4630;
assign na3962 = ~a3962;
assign na3940 = ~a3940;
assign na3922 = ~a3922;
assign na3904 = ~a3904;
assign na3886 = ~a3886;
assign na3868 = ~a3868;
assign na3850 = ~a3850;
assign na4786 = ~a4786;
assign na4816 = ~a4816;
assign na4842 = ~a4842;
assign na4868 = ~a4868;
assign na4898 = ~a4898;
assign na4920 = ~a4920;
assign na4942 = ~a4942;
assign na4960 = ~a4960;
assign na4982 = ~a4982;
assign na3838 = ~a3838;
assign na4976 = ~a4976;
assign na4954 = ~a4954;
assign na4936 = ~a4936;
assign na4914 = ~a4914;
assign na4892 = ~a4892;
assign na4862 = ~a4862;
assign na4836 = ~a4836;
assign na4810 = ~a4810;
assign na4780 = ~a4780;
assign na3814 = ~a3814;
assign na3780 = ~a3780;
assign na3668 = ~a3668;
assign na3644 = ~a3644;
assign na4994 = ~a4994;
assign na3544 = ~a3544;
assign na5006 = ~a5006;
assign na4988 = ~a4988;
assign na5018 = ~a5018;
assign na5000 = ~a5000;
assign na5030 = ~a5030;
assign na5012 = ~a5012;
assign na5042 = ~a5042;
assign na5024 = ~a5024;
assign na5054 = ~a5054;
assign na5036 = ~a5036;
assign na5066 = ~a5066;
assign na5048 = ~a5048;
assign na5078 = ~a5078;
assign na5060 = ~a5060;
assign na5090 = ~a5090;
assign na5072 = ~a5072;
assign na5102 = ~a5102;
assign na5084 = ~a5084;
assign na5114 = ~a5114;
assign na5096 = ~a5096;
assign na5108 = ~a5108;
assign na3514 = ~a3514;
assign na3492 = ~a3492;
assign na3474 = ~a3474;
assign na3456 = ~a3456;
assign na3438 = ~a3438;
assign na3420 = ~a3420;
assign na3402 = ~a3402;
assign na3384 = ~a3384;
assign na3366 = ~a3366;
assign na3348 = ~a3348;
assign na3330 = ~a3330;
assign na3312 = ~a3312;
assign na3294 = ~a3294;
assign a3276 = ~a3274 & ~a3266;
assign na5120 = ~a5120;
assign c1 = 1;
assign a822 = l80 & ~l78;
assign a824 = ~l80 & l78;
assign a826 = ~a824 & ~a822;
assign a828 = l470 & ~l84;
assign a830 = a828 & l86;
assign a832 = ~a830 & i2;
assign a834 = ~l474 & ~l472;
assign a836 = ~l478 & l476;
assign a838 = a836 & a834;
assign a840 = l482 & l480;
assign a842 = ~l486 & ~l484;
assign a844 = l490 & l488;
assign a846 = a844 & a842;
assign a848 = a846 & a840;
assign a850 = ~l488 & l486;
assign a852 = a850 & ~l484;
assign a854 = a852 & l490;
assign a856 = a854 & ~a840;
assign a858 = ~a856 & ~a848;
assign a860 = ~a858 & a838;
assign a862 = a850 & l484;
assign a864 = a862 & ~l480;
assign a866 = a864 & ~l490;
assign a868 = a840 & ~l490;
assign a870 = a868 & a852;
assign a872 = ~a870 & ~a866;
assign a874 = a872 & ~a860;
assign a876 = l474 & l472;
assign a878 = a876 & ~l476;
assign a880 = a878 & ~l478;
assign a882 = a842 & ~l480;
assign a884 = ~l490 & ~l488;
assign a886 = a884 & l482;
assign a888 = a886 & a882;
assign a890 = a888 & ~l108;
assign a892 = a890 & a880;
assign a894 = a840 & l490;
assign a896 = a894 & a862;
assign a898 = a882 & ~l482;
assign a900 = a898 & l488;
assign a902 = a838 & l482;
assign a904 = a846 & l480;
assign a906 = a904 & ~a902;
assign a908 = ~a906 & ~a900;
assign a910 = a908 & ~a896;
assign a912 = a854 & ~a838;
assign a914 = ~a912 & a910;
assign a916 = a914 & ~a892;
assign a918 = ~l492 & ~l482;
assign a920 = ~a918 & l490;
assign a922 = a920 & a864;
assign a924 = ~a922 & ~a866;
assign a926 = a924 & a916;
assign a928 = l474 & ~l472;
assign a930 = a928 & l494;
assign a932 = a930 & ~a926;
assign a934 = ~a932 & a874;
assign a936 = ~l474 & l472;
assign a938 = a876 & l498;
assign a940 = ~a938 & ~a936;
assign a942 = ~a940 & a836;
assign a944 = a936 & ~l476;
assign a946 = ~a944 & ~a880;
assign a948 = a946 & ~a942;
assign a950 = ~a922 & ~a854;
assign a952 = a950 & ~a866;
assign a954 = ~a952 & ~a948;
assign a956 = ~a954 & ~a860;
assign a958 = ~a956 & l500;
assign a960 = a842 & l480;
assign a962 = a960 & a884;
assign a964 = a898 & ~l488;
assign a966 = ~a964 & ~a888;
assign a968 = a966 & ~a962;
assign a970 = a900 & ~l490;
assign a972 = a928 & ~l476;
assign a974 = a972 & l478;
assign a976 = a974 & ~l494;
assign a978 = ~a976 & ~l472;
assign a980 = ~a978 & a970;
assign a982 = ~a980 & a968;
assign a984 = ~l504 & ~l500;
assign a986 = a984 & ~l502;
assign a988 = ~a986 & ~a982;
assign a990 = ~a988 & ~a958;
assign a992 = l508 & l506;
assign a994 = a992 & ~a990;
assign a996 = ~a994 & l496;
assign a998 = a996 & ~a922;
assign a1000 = a998 & a934;
assign a1002 = ~a994 & ~l496;
assign a1004 = a1002 & l78;
assign a1006 = ~a1004 & ~a1000;
assign a1008 = ~a1006 & l86;
assign a1010 = l510 & ~l86;
assign a1012 = ~a1010 & ~a1008;
assign a1014 = ~a1012 & a832;
assign a1016 = ~a832 & l78;
assign a1018 = ~a1016 & ~a1014;
assign a1020 = ~l84 & l82;
assign a1022 = a1020 & l86;
assign a1024 = ~a1022 & i2;
assign a1026 = ~l90 & ~l88;
assign a1028 = ~l94 & l92;
assign a1030 = a1028 & a1026;
assign a1032 = l98 & l96;
assign a1034 = ~l102 & ~l100;
assign a1036 = l106 & l104;
assign a1038 = a1036 & a1034;
assign a1040 = a1038 & a1032;
assign a1042 = ~l104 & l102;
assign a1044 = a1042 & ~l100;
assign a1046 = a1044 & l106;
assign a1048 = a1046 & ~a1032;
assign a1050 = ~a1048 & ~a1040;
assign a1052 = ~a1050 & a1030;
assign a1054 = a1042 & l100;
assign a1056 = a1054 & ~l96;
assign a1058 = a1056 & ~l106;
assign a1060 = a1032 & ~l106;
assign a1062 = a1060 & a1044;
assign a1064 = ~a1062 & ~a1058;
assign a1066 = a1064 & ~a1052;
assign a1068 = l90 & l88;
assign a1070 = ~l94 & ~l92;
assign a1072 = a1070 & a1068;
assign a1074 = a1034 & ~l96;
assign a1076 = ~l106 & ~l104;
assign a1078 = a1076 & l98;
assign a1080 = a1078 & a1074;
assign a1082 = a1080 & ~l108;
assign a1084 = a1082 & a1072;
assign a1086 = a1032 & l106;
assign a1088 = a1086 & a1054;
assign a1090 = a1074 & ~l98;
assign a1092 = a1090 & l104;
assign a1094 = a1030 & l98;
assign a1096 = a1038 & l96;
assign a1098 = a1096 & ~a1094;
assign a1100 = ~a1098 & ~a1092;
assign a1102 = a1100 & ~a1088;
assign a1104 = a1046 & ~a1030;
assign a1106 = ~a1104 & a1102;
assign a1108 = a1106 & ~a1084;
assign a1110 = ~l110 & ~l98;
assign a1112 = ~a1110 & l106;
assign a1114 = a1112 & a1056;
assign a1116 = ~a1114 & ~a1058;
assign a1118 = a1116 & a1108;
assign a1120 = l90 & ~l88;
assign a1122 = a1120 & l112;
assign a1124 = a1122 & ~a1118;
assign a1126 = ~a1124 & a1066;
assign a1128 = ~l90 & l88;
assign a1130 = a1128 & ~l92;
assign a1132 = a1068 & l116;
assign a1134 = ~a1132 & ~a1128;
assign a1136 = ~a1134 & a1028;
assign a1138 = ~a1136 & ~a1072;
assign a1140 = a1138 & ~a1130;
assign a1142 = ~a1114 & ~a1046;
assign a1144 = a1142 & ~a1058;
assign a1146 = ~a1144 & ~a1140;
assign a1148 = ~a1146 & ~a1052;
assign a1150 = ~a1148 & l118;
assign a1152 = ~l122 & ~l118;
assign a1154 = a1152 & ~l120;
assign a1156 = a1092 & ~l106;
assign a1158 = l94 & ~l92;
assign a1160 = a1158 & a1120;
assign a1162 = a1160 & ~l112;
assign a1164 = ~a1162 & ~l88;
assign a1166 = ~a1164 & a1156;
assign a1168 = a1034 & l96;
assign a1170 = a1168 & a1076;
assign a1172 = a1090 & ~l104;
assign a1174 = ~a1172 & ~a1080;
assign a1176 = a1174 & ~a1170;
assign a1178 = l102 & l100;
assign a1180 = a1036 & a1032;
assign a1182 = a1180 & a1178;
assign a1184 = ~a1182 & a1176;
assign a1186 = a1184 & ~a1166;
assign a1188 = ~a1186 & ~a1154;
assign a1190 = ~a1188 & ~a1150;
assign a1192 = l126 & l124;
assign a1194 = a1192 & ~a1190;
assign a1196 = ~a1194 & l114;
assign a1198 = a1196 & ~a1114;
assign a1200 = a1198 & a1126;
assign a1202 = ~a1194 & ~l114;
assign a1204 = a1202 & l80;
assign a1206 = ~a1204 & ~a1200;
assign a1208 = ~a1206 & l86;
assign a1210 = l128 & ~l86;
assign a1212 = ~a1210 & ~a1208;
assign a1214 = ~a1212 & a1024;
assign a1216 = ~a1024 & l80;
assign a1218 = ~a1216 & ~a1214;
assign a1220 = ~l464 & ~l86;
assign a1222 = l230 & l156;
assign a1224 = ~a1222 & l86;
assign a1226 = ~a1020 & l466;
assign a1228 = a1226 & a1224;
assign a1232 = a1230 & a1024;
assign a1234 = ~a1024 & l82;
assign a1236 = ~a1234 & ~a1232;
assign a1238 = l86 & i76;
assign a1240 = l462 & ~l86;
assign a1242 = ~a1240 & ~a1238;
assign a1244 = ~a1242 & i2;
assign a1246 = l84 & ~i2;
assign a1248 = ~a1246 & ~a1244;
assign a1250 = l86 & i18;
assign a1252 = ~a1250 & i2;
assign a1254 = a1020 & i74;
assign a1256 = ~a1020 & l88;
assign a1258 = ~a1256 & ~a1254;
assign a1260 = ~a1258 & l86;
assign a1262 = l460 & ~l86;
assign a1264 = ~a1262 & ~a1260;
assign a1266 = ~a1264 & a1252;
assign a1268 = ~a1252 & l88;
assign a1270 = ~a1268 & ~a1266;
assign a1272 = a1020 & i72;
assign a1274 = ~a1020 & l90;
assign a1276 = ~a1274 & ~a1272;
assign a1278 = ~a1276 & l86;
assign a1280 = l458 & ~l86;
assign a1282 = ~a1280 & ~a1278;
assign a1284 = ~a1282 & a1252;
assign a1286 = ~a1252 & l90;
assign a1288 = ~a1286 & ~a1284;
assign a1290 = a1020 & i70;
assign a1292 = ~a1020 & l92;
assign a1294 = ~a1292 & ~a1290;
assign a1296 = ~a1294 & l86;
assign a1298 = l456 & ~l86;
assign a1300 = ~a1298 & ~a1296;
assign a1302 = ~a1300 & a1252;
assign a1304 = ~a1252 & l92;
assign a1306 = ~a1304 & ~a1302;
assign a1308 = a1020 & i68;
assign a1310 = ~a1020 & l94;
assign a1312 = ~a1310 & ~a1308;
assign a1314 = ~a1312 & l86;
assign a1316 = l454 & ~l86;
assign a1318 = ~a1316 & ~a1314;
assign a1320 = ~a1318 & a1252;
assign a1322 = ~a1252 & l94;
assign a1324 = ~a1322 & ~a1320;
assign a1326 = i58 & i56;
assign a1328 = a1326 & i62;
assign a1330 = a1328 & i60;
assign a1332 = a1330 & i64;
assign a1334 = ~a1332 & i66;
assign a1336 = a1334 & a1020;
assign a1338 = ~a1020 & l96;
assign a1340 = ~a1338 & ~a1336;
assign a1342 = ~a1340 & l86;
assign a1344 = l452 & ~l86;
assign a1346 = ~a1344 & ~a1342;
assign a1348 = ~a1346 & a1252;
assign a1350 = ~a1252 & l96;
assign a1352 = ~a1350 & ~a1348;
assign a1354 = a1020 & i64;
assign a1356 = ~a1020 & l98;
assign a1358 = ~a1356 & ~a1354;
assign a1360 = ~a1358 & l86;
assign a1362 = l450 & ~l86;
assign a1364 = ~a1362 & ~a1360;
assign a1366 = ~a1364 & a1252;
assign a1368 = ~a1252 & l98;
assign a1370 = ~a1368 & ~a1366;
assign a1372 = a1020 & i62;
assign a1374 = ~a1020 & l100;
assign a1376 = ~a1374 & ~a1372;
assign a1378 = ~a1376 & l86;
assign a1380 = l448 & ~l86;
assign a1382 = ~a1380 & ~a1378;
assign a1384 = ~a1382 & a1252;
assign a1386 = ~a1252 & l100;
assign a1388 = ~a1386 & ~a1384;
assign a1390 = a1020 & i60;
assign a1392 = ~a1020 & l102;
assign a1394 = ~a1392 & ~a1390;
assign a1396 = ~a1394 & l86;
assign a1398 = l446 & ~l86;
assign a1400 = ~a1398 & ~a1396;
assign a1402 = ~a1400 & a1252;
assign a1404 = ~a1252 & l102;
assign a1406 = ~a1404 & ~a1402;
assign a1408 = a1020 & i58;
assign a1410 = ~a1020 & l104;
assign a1412 = ~a1410 & ~a1408;
assign a1414 = ~a1412 & l86;
assign a1416 = l444 & ~l86;
assign a1418 = ~a1416 & ~a1414;
assign a1420 = ~a1418 & a1252;
assign a1422 = ~a1252 & l104;
assign a1424 = ~a1422 & ~a1420;
assign a1426 = a1020 & i56;
assign a1428 = ~a1020 & l106;
assign a1430 = ~a1428 & ~a1426;
assign a1432 = ~a1430 & l86;
assign a1434 = l442 & ~l86;
assign a1436 = ~a1434 & ~a1432;
assign a1438 = ~a1436 & a1252;
assign a1440 = ~a1252 & l106;
assign a1442 = ~a1440 & ~a1438;
assign a1444 = l84 & i54;
assign a1446 = l108 & ~l84;
assign a1448 = ~a1446 & ~a1444;
assign a1450 = ~a1448 & l86;
assign a1452 = l440 & ~l86;
assign a1454 = ~a1452 & ~a1450;
assign a1456 = ~a1454 & a1024;
assign a1458 = ~a1024 & l108;
assign a1460 = ~a1458 & ~a1456;
assign a1462 = a1020 & i52;
assign a1464 = ~a1020 & l110;
assign a1466 = ~a1464 & ~a1462;
assign a1468 = ~a1466 & l86;
assign a1470 = l438 & ~l86;
assign a1472 = ~a1470 & ~a1468;
assign a1474 = ~a1472 & a1252;
assign a1476 = ~a1252 & l110;
assign a1478 = ~a1476 & ~a1474;
assign a1480 = a1020 & i50;
assign a1482 = ~a1020 & l112;
assign a1484 = ~a1482 & ~a1480;
assign a1486 = ~a1484 & l86;
assign a1488 = l436 & ~l86;
assign a1490 = ~a1488 & ~a1486;
assign a1492 = ~a1490 & a1252;
assign a1494 = ~a1252 & l112;
assign a1496 = ~a1494 & ~a1492;
assign a1498 = l86 & l84;
assign a1500 = l434 & ~l86;
assign a1502 = ~a1500 & ~a1498;
assign a1504 = ~a1502 & a1024;
assign a1506 = ~a1024 & l114;
assign a1508 = ~a1506 & ~a1504;
assign a1510 = a1020 & i48;
assign a1512 = ~a1020 & l116;
assign a1514 = ~a1512 & ~a1510;
assign a1516 = ~a1514 & l86;
assign a1518 = l432 & ~l86;
assign a1520 = ~a1518 & ~a1516;
assign a1522 = ~a1520 & a1252;
assign a1524 = ~a1252 & l116;
assign a1526 = ~a1524 & ~a1522;
assign a1528 = l86 & i46;
assign a1530 = l430 & ~l86;
assign a1532 = ~a1530 & ~a1528;
assign a1534 = ~a1532 & a1024;
assign a1536 = ~a1024 & l118;
assign a1538 = ~a1536 & ~a1534;
assign a1540 = l86 & i44;
assign a1542 = l428 & ~l86;
assign a1544 = ~a1542 & ~a1540;
assign a1546 = ~a1544 & a1024;
assign a1548 = ~a1024 & l120;
assign a1550 = ~a1548 & ~a1546;
assign a1552 = l86 & i42;
assign a1554 = l426 & ~l86;
assign a1556 = ~a1554 & ~a1552;
assign a1558 = ~a1556 & a1024;
assign a1560 = ~a1024 & l122;
assign a1562 = ~a1560 & ~a1558;
assign a1564 = l380 & l86;
assign a1566 = l382 & ~l86;
assign a1568 = ~a1566 & ~a1564;
assign a1570 = ~a1568 & a1024;
assign a1572 = ~a1024 & l124;
assign a1574 = ~a1572 & ~a1570;
assign a1576 = ~l140 & ~l138;
assign a1578 = a1576 & ~l136;
assign a1580 = ~a1578 & ~l134;
assign a1582 = ~l148 & ~l146;
assign a1584 = a1582 & l144;
assign a1586 = a1584 & ~l142;
assign a1588 = l150 & l142;
assign a1590 = a1582 & ~l144;
assign a1592 = a1590 & a1588;
assign a1594 = ~a1592 & ~a1586;
assign a1596 = ~a1594 & a1156;
assign a1598 = ~l150 & l142;
assign a1600 = ~l148 & l146;
assign a1602 = a1600 & ~l144;
assign a1604 = ~a1602 & ~a1584;
assign a1606 = ~a1604 & a1598;
assign a1608 = a1606 & ~a1176;
assign a1610 = ~a1608 & ~a1596;
assign a1612 = a1610 & a1580;
assign a1614 = a1176 & ~a1156;
assign a1616 = ~a1614 & a1128;
assign a1618 = a1616 & a1612;
assign a1620 = a1618 & l132;
assign a1622 = a1620 & l154;
assign a1624 = ~l156 & l152;
assign a1626 = l160 & l158;
assign a1628 = ~a1626 & ~a1624;
assign a1630 = a1176 & ~a1166;
assign a1632 = a1630 & l114;
assign a1634 = a1130 & l94;
assign a1636 = ~a1634 & a1146;
assign a1638 = ~a1636 & a1632;
assign a1640 = ~a1638 & a1628;
assign a1642 = a1640 & ~a1622;
assign a1644 = a1642 & ~l152;
assign a1646 = ~a1644 & ~a1620;
assign a1648 = ~a1646 & ~a1182;
assign a1650 = ~a1648 & l130;
assign a1652 = l126 & ~l124;
assign a1654 = ~a1652 & ~a1650;
assign a1656 = ~a1654 & l86;
assign a1658 = l162 & ~l86;
assign a1660 = ~a1658 & ~a1656;
assign a1662 = ~a1660 & a1024;
assign a1664 = ~a1024 & l126;
assign a1666 = ~a1664 & ~a1662;
assign a1668 = ~a1636 & a1630;
assign a1670 = a1668 & ~a1182;
assign a1672 = ~a1670 & l294;
assign a1674 = a1672 & l114;
assign a1676 = ~a1620 & l130;
assign a1678 = a1676 & a1648;
assign a1680 = ~a1678 & ~a1674;
assign a1682 = ~a1680 & l86;
assign a1684 = l378 & ~l86;
assign a1686 = ~a1684 & ~a1682;
assign a1688 = ~a1686 & a1024;
assign a1690 = ~a1024 & l130;
assign a1692 = ~a1690 & ~a1688;
assign a1694 = ~a1630 & l114;
assign a1696 = ~a1610 & a1580;
assign a1698 = ~a1696 & a1616;
assign a1700 = a1698 & l132;
assign a1702 = a1700 & ~a1618;
assign a1704 = ~a1702 & ~a1694;
assign a1706 = ~a1704 & l86;
assign a1708 = l376 & ~l86;
assign a1710 = ~a1708 & ~a1706;
assign a1712 = ~a1710 & a1024;
assign a1714 = ~a1024 & l132;
assign a1716 = ~a1714 & ~a1712;
assign a1718 = a1600 & l144;
assign a1720 = l112 & l88;
assign a1722 = a1720 & ~a1108;
assign a1724 = a1128 & l94;
assign a1726 = ~a1184 & ~l92;
assign a1728 = a1726 & a1724;
assign a1730 = a1724 & l92;
assign a1732 = a1158 & a1068;
assign a1734 = ~a1732 & ~a1730;
assign a1736 = ~a1734 & ~a1176;
assign a1738 = a1736 & l112;
assign a1740 = ~a1738 & ~a1728;
assign a1742 = a1740 & ~a1722;
assign a1744 = ~a1742 & l178;
assign a1746 = ~a1634 & ~a1052;
assign a1748 = ~a1746 & ~l178;
assign a1750 = ~a1748 & ~a1744;
assign a1752 = a1750 & l150;
assign a1754 = ~a1752 & ~l142;
assign a1756 = ~a1754 & ~a1588;
assign a1758 = a1756 & a1718;
assign a1760 = a1758 & a1580;
assign a1762 = a1760 & l180;
assign a1764 = a1762 & l140;
assign a1766 = l198 & ~l156;
assign a1768 = l200 & i10;
assign a1770 = ~a1768 & ~a1766;
assign a1772 = a1770 & ~a1632;
assign a1774 = a1772 & ~a1620;
assign a1776 = a1774 & ~l198;
assign a1778 = ~a1182 & l114;
assign a1780 = l202 & ~l156;
assign a1782 = l204 & i12;
assign a1784 = ~a1782 & ~a1780;
assign a1786 = a1784 & ~a1778;
assign a1788 = a1786 & ~l202;
assign a1790 = ~a1788 & l138;
assign a1792 = a1790 & ~a1776;
assign a1794 = a1792 & l196;
assign a1796 = l206 & l178;
assign a1798 = a1796 & a1794;
assign a1800 = l134 & i30;
assign a1802 = ~l184 & ~l170;
assign a1804 = a1802 & ~l212;
assign a1806 = a1804 & ~l192;
assign a1808 = ~a1806 & ~l180;
assign a1810 = ~a1808 & a1800;
assign a1812 = ~a1810 & l134;
assign a1814 = l106 & l90;
assign a1816 = ~a1814 & a1092;
assign a1818 = ~a1816 & ~a1098;
assign a1820 = ~a1818 & l88;
assign a1822 = ~a1820 & a1176;
assign a1824 = a1822 & a1148;
assign a1826 = ~a1824 & l114;
assign a1828 = ~a1826 & ~a1812;
assign a1830 = a1828 & ~a1798;
assign a1832 = a1830 & ~a1764;
assign a1834 = ~a1832 & l86;
assign a1836 = l374 & ~l86;
assign a1838 = ~a1836 & ~a1834;
assign a1840 = ~a1838 & a1024;
assign a1842 = ~a1024 & l134;
assign a1844 = ~a1842 & ~a1840;
assign a1846 = ~a1762 & l140;
assign a1848 = ~l336 & ~l334;
assign a1850 = ~l340 & ~l338;
assign a1852 = a1850 & a1848;
assign a1854 = ~l344 & ~l342;
assign a1856 = ~l348 & ~l346;
assign a1858 = a1856 & ~l350;
assign a1860 = a1858 & a1854;
assign a1862 = a1860 & a1852;
assign a1864 = ~a1862 & l136;
assign a1866 = ~a1864 & ~a1846;
assign a1868 = ~a1866 & l86;
assign a1870 = l372 & ~l86;
assign a1872 = ~a1870 & ~a1868;
assign a1874 = ~a1872 & a1024;
assign a1876 = ~a1024 & l136;
assign a1878 = ~a1876 & ~a1874;
assign a1880 = ~a1798 & ~l156;
assign a1882 = a1880 & l138;
assign a1884 = a1862 & l136;
assign a1886 = a1824 & l114;
assign a1888 = ~a1886 & ~a1884;
assign a1890 = a1888 & ~a1882;
assign a1892 = ~a1890 & l86;
assign a1894 = l352 & ~l86;
assign a1896 = ~a1894 & ~a1892;
assign a1898 = ~a1896 & a1024;
assign a1900 = ~a1024 & l138;
assign a1902 = ~a1900 & ~a1898;
assign a1904 = a1810 & l86;
assign a1906 = l332 & ~l86;
assign a1908 = ~a1906 & ~a1904;
assign a1910 = ~a1908 & a1024;
assign a1912 = ~a1024 & l140;
assign a1914 = ~a1912 & ~a1910;
assign a1916 = a1810 & i40;
assign a1918 = ~a1810 & l142;
assign a1920 = ~a1918 & ~a1916;
assign a1922 = ~a1920 & l86;
assign a1924 = l330 & ~l86;
assign a1926 = ~a1924 & ~a1922;
assign a1928 = ~a1926 & a1024;
assign a1930 = ~a1024 & l142;
assign a1932 = ~a1930 & ~a1928;
assign a1934 = a1810 & i38;
assign a1936 = ~a1810 & l144;
assign a1938 = ~a1936 & ~a1934;
assign a1940 = ~a1938 & l86;
assign a1942 = l328 & ~l86;
assign a1944 = ~a1942 & ~a1940;
assign a1946 = ~a1944 & a1024;
assign a1948 = ~a1024 & l144;
assign a1950 = ~a1948 & ~a1946;
assign a1952 = a1810 & i36;
assign a1954 = ~a1810 & l146;
assign a1956 = ~a1954 & ~a1952;
assign a1958 = ~a1956 & l86;
assign a1960 = l326 & ~l86;
assign a1962 = ~a1960 & ~a1958;
assign a1964 = ~a1962 & a1024;
assign a1966 = ~a1024 & l146;
assign a1968 = ~a1966 & ~a1964;
assign a1970 = a1810 & i34;
assign a1972 = ~a1810 & l148;
assign a1974 = ~a1972 & ~a1970;
assign a1976 = ~a1974 & l86;
assign a1978 = l324 & ~l86;
assign a1980 = ~a1978 & ~a1976;
assign a1982 = ~a1980 & a1024;
assign a1984 = ~a1024 & l148;
assign a1986 = ~a1984 & ~a1982;
assign a1988 = a1810 & i32;
assign a1990 = ~a1810 & l150;
assign a1992 = ~a1990 & ~a1988;
assign a1994 = ~a1992 & l86;
assign a1996 = l322 & ~l86;
assign a1998 = ~a1996 & ~a1994;
assign a2000 = ~a1998 & a1024;
assign a2002 = ~a1024 & l150;
assign a2004 = ~a2002 & ~a2000;
assign a2006 = ~a1642 & l86;
assign a2008 = l320 & ~l86;
assign a2010 = ~a2008 & ~a2006;
assign a2012 = ~a2010 & a1024;
assign a2014 = ~a1024 & l152;
assign a2016 = ~a2014 & ~a2012;
assign a2018 = ~a1668 & l84;
assign a2020 = ~l172 & ~l170;
assign a2022 = a2020 & l154;
assign a2024 = a2022 & ~a1620;
assign a2026 = ~a2024 & ~a2018;
assign a2028 = ~a2026 & l86;
assign a2030 = l318 & ~l86;
assign a2032 = ~a2030 & ~a2028;
assign a2034 = ~a2032 & a1024;
assign a2036 = ~a1024 & l154;
assign a2038 = ~a2036 & ~a2034;
assign a2040 = l112 & l92;
assign a2042 = ~a2040 & a1128;
assign a2044 = a2042 & ~a1176;
assign a2046 = a1182 & ~a1068;
assign a2048 = a1170 & a1160;
assign a2050 = a2048 & ~l112;
assign a2052 = ~a2050 & ~a2046;
assign a2054 = a2052 & ~a2044;
assign a2056 = l218 & l206;
assign a2058 = a2056 & a1794;
assign a2060 = ~a2058 & ~a1798;
assign a2062 = ~a2060 & ~a2054;
assign a2064 = l284 & ~l156;
assign a2066 = a2064 & ~a2062;
assign a2068 = l288 & l286;
assign a2070 = a2040 & a1128;
assign a2072 = ~a2070 & ~a1068;
assign a2074 = a2072 & ~a1160;
assign a2076 = ~a2074 & ~a1174;
assign a2078 = a1182 & a1068;
assign a2080 = ~a2072 & a1170;
assign a2082 = ~a2080 & ~a2078;
assign a2084 = a2082 & ~a2076;
assign a2086 = a1142 & a1102;
assign a2088 = a2086 & a1066;
assign a2090 = a2088 & a2084;
assign a2092 = a2090 & l114;
assign a2094 = ~a2092 & ~a2068;
assign a2096 = a2094 & ~a2066;
assign a2098 = a2096 & ~l284;
assign a2100 = l290 & l86;
assign a2102 = a2100 & a1792;
assign a2104 = a2102 & ~a2098;
assign a2106 = a1580 & l180;
assign a2108 = a2106 & ~a1758;
assign a2110 = a2108 & ~a1750;
assign a2112 = a1880 & l208;
assign a2114 = l212 & i14;
assign a2116 = a1148 & l114;
assign a2118 = ~a2116 & ~a2114;
assign a2120 = a2118 & ~a2112;
assign a2122 = a2120 & ~a2110;
assign a2124 = a2122 & ~l208;
assign a2126 = ~a1750 & a1722;
assign a2128 = ~a2126 & a1798;
assign a2130 = ~a2128 & ~a2058;
assign a2132 = l196 & ~l156;
assign a2134 = a2132 & a2130;
assign a2136 = l258 & l256;
assign a2138 = ~l264 & ~l262;
assign a2140 = a2138 & l260;
assign a2142 = ~a2140 & ~a2136;
assign a2144 = a1118 & l114;
assign a2146 = ~a2144 & a2142;
assign a2148 = a2146 & ~a2134;
assign a2150 = a2148 & ~l196;
assign a2152 = ~a2150 & ~a1644;
assign a2154 = a2152 & ~a2124;
assign a2156 = a2154 & a2104;
assign a2158 = l292 & ~l86;
assign a2160 = ~a2158 & ~a2156;
assign a2162 = ~a2160 & a1024;
assign a2164 = ~a1024 & l156;
assign a2166 = ~a2164 & ~a2162;
assign a2168 = ~l160 & l158;
assign a2170 = ~a2168 & ~l166;
assign a2172 = ~a2170 & l86;
assign a2174 = l168 & ~l86;
assign a2176 = ~a2174 & ~a2172;
assign a2178 = ~a2176 & a1024;
assign a2180 = ~a1024 & l158;
assign a2182 = ~a2180 & ~a2178;
assign a2184 = l86 & i4;
assign a2186 = l164 & ~l86;
assign a2188 = ~a2186 & ~a2184;
assign a2190 = ~a2188 & a1024;
assign a2192 = ~a1024 & l160;
assign a2194 = ~a2192 & ~a2190;
assign a2196 = l154 & l86;
assign a2198 = a2196 & ~a2020;
assign a2200 = l174 & ~l86;
assign a2202 = ~a2200 & ~a2198;
assign a2204 = ~a2202 & a1024;
assign a2206 = ~a1024 & l166;
assign a2208 = ~a2206 & ~a2204;
assign a2210 = a1750 & l86;
assign a2212 = a2210 & a2108;
assign a2214 = l182 & ~l86;
assign a2216 = ~a2214 & ~a2212;
assign a2218 = ~a2216 & a1024;
assign a2220 = ~a1024 & l170;
assign a2222 = ~a2220 & ~a2218;
assign a2224 = l132 & l86;
assign a2226 = a2224 & ~a1698;
assign a2228 = l176 & ~l86;
assign a2230 = ~a2228 & ~a2226;
assign a2232 = ~a2230 & a1024;
assign a2234 = ~a1024 & l172;
assign a2236 = ~a2234 & ~a2232;
assign a2238 = l226 & l222;
assign a2240 = ~l224 & ~l222;
assign a2242 = ~a2240 & ~l228;
assign a2244 = a2242 & ~a2238;
assign a2246 = a2244 & ~a1630;
assign a2248 = a1182 & ~a1140;
assign a2250 = ~a2248 & l124;
assign a2252 = a2250 & ~a2246;
assign a2254 = ~l178 & ~l124;
assign a2256 = ~a2254 & a1224;
assign a2258 = a2256 & ~a2252;
assign a2260 = l282 & ~l86;
assign a2262 = ~a2260 & ~a2258;
assign a2264 = ~a2262 & a1024;
assign a2266 = ~a1024 & l178;
assign a2268 = ~a2266 & ~a2264;
assign a2270 = ~l186 & l184;
assign a2272 = ~a1580 & l180;
assign a2274 = ~a2272 & ~a2270;
assign a2276 = ~a2274 & l86;
assign a2278 = l188 & ~l86;
assign a2280 = ~a2278 & ~a2276;
assign a2282 = ~a2280 & a1024;
assign a2284 = ~a1024 & l180;
assign a2286 = ~a2284 & ~a2282;
assign a2288 = l186 & l184;
assign a2290 = ~a2288 & ~l192;
assign a2292 = a2290 & ~a1762;
assign a2294 = ~a2292 & l86;
assign a2296 = l194 & ~l86;
assign a2298 = ~a2296 & ~a2294;
assign a2300 = ~a2298 & a1024;
assign a2302 = ~a1024 & l184;
assign a2304 = ~a2302 & ~a2300;
assign a2306 = a1760 & i6;
assign a2308 = ~a2306 & ~l186;
assign a2310 = ~a1760 & i8;
assign a2312 = l86 & ~l82;
assign a2314 = a2312 & ~a2310;
assign a2316 = a2314 & ~a2308;
assign a2318 = l190 & ~l86;
assign a2320 = ~a2318 & ~a2316;
assign a2322 = ~a2320 & a1024;
assign a2324 = ~a1024 & l186;
assign a2326 = ~a2324 & ~a2322;
assign a2328 = a1798 & l208;
assign a2330 = ~a1148 & l114;
assign a2332 = ~a2330 & ~a2328;
assign a2334 = ~a2332 & l86;
assign a2336 = l210 & ~l86;
assign a2338 = ~a2336 & ~a2334;
assign a2340 = ~a2338 & a1024;
assign a2342 = ~a1024 & l192;
assign a2344 = ~a2342 & ~a2340;
assign a2346 = ~a2148 & l86;
assign a2348 = l266 & ~l86;
assign a2350 = ~a2348 & ~a2346;
assign a2352 = ~a2350 & a1024;
assign a2354 = ~a1024 & l196;
assign a2356 = ~a2354 & ~a2352;
assign a2358 = ~a1774 & l86;
assign a2360 = l254 & ~l86;
assign a2362 = ~a2360 & ~a2358;
assign a2364 = ~a2362 & a1024;
assign a2366 = ~a1024 & l198;
assign a2368 = ~a2366 & ~a2364;
assign a2370 = l200 & ~i10;
assign a2372 = ~a2370 & ~l172;
assign a2374 = ~a2372 & l86;
assign a2376 = l252 & ~l86;
assign a2378 = ~a2376 & ~a2374;
assign a2380 = ~a2378 & a1024;
assign a2382 = ~a1024 & l200;
assign a2384 = ~a2382 & ~a2380;
assign a2386 = ~a1786 & l86;
assign a2388 = l250 & ~l86;
assign a2390 = ~a2388 & ~a2386;
assign a2392 = ~a2390 & a1024;
assign a2394 = ~a1024 & l202;
assign a2396 = ~a2394 & ~a2392;
assign a2398 = a1182 & l114;
assign a2400 = l204 & ~i12;
assign a2402 = ~a2400 & ~a2398;
assign a2404 = ~a2402 & l86;
assign a2406 = l248 & ~l86;
assign a2408 = ~a2406 & ~a2404;
assign a2410 = ~a2408 & a1024;
assign a2412 = ~a1024 & l204;
assign a2414 = ~a2412 & ~a2410;
assign a2416 = ~l218 & ~l178;
assign a2418 = ~a2416 & l206;
assign a2420 = a2418 & ~a1794;
assign a2422 = ~a2420 & ~a1194;
assign a2424 = ~a2422 & l86;
assign a2426 = l220 & ~l86;
assign a2428 = ~a2426 & ~a2424;
assign a2430 = ~a2428 & a1024;
assign a2432 = ~a1024 & l206;
assign a2434 = ~a2432 & ~a2430;
assign a2436 = ~a2122 & l86;
assign a2438 = l214 & ~l86;
assign a2440 = ~a2438 & ~a2436;
assign a2442 = ~a2440 & a1024;
assign a2444 = ~a1024 & l208;
assign a2446 = ~a2444 & ~a2442;
assign a2448 = l212 & ~i14;
assign a2450 = ~a2448 & ~l170;
assign a2452 = ~a2450 & l86;
assign a2454 = l216 & ~l86;
assign a2456 = ~a2454 & ~a2452;
assign a2458 = ~a2456 & a1024;
assign a2460 = ~a1024 & l212;
assign a2462 = ~a2460 & ~a2458;
assign a2464 = l228 & ~l226;
assign a2466 = a2464 & a2240;
assign a2468 = ~l228 & l224;
assign a2470 = a2468 & a2238;
assign a2472 = ~a2470 & ~a2466;
assign a2474 = ~a2472 & ~a1630;
assign a2476 = a1734 & ~a1120;
assign a2478 = ~a2476 & a1182;
assign a2480 = ~a2048 & l124;
assign a2482 = a2480 & ~a2478;
assign a2484 = a2482 & ~a2474;
assign a2486 = ~l218 & ~l124;
assign a2488 = ~a2486 & a1224;
assign a2490 = a2488 & ~a2484;
assign a2492 = l232 & ~l86;
assign a2494 = ~a2492 & ~a2490;
assign a2496 = ~a2494 & a1024;
assign a2498 = ~a1024 & l218;
assign a2500 = ~a2498 & ~a2496;
assign a2502 = ~a1026 & ~l112;
assign a2504 = a2502 & ~a1108;
assign a2506 = ~a2504 & ~a1722;
assign a2508 = ~a1734 & a1182;
assign a2510 = a1736 & ~l112;
assign a2512 = ~a2510 & ~a2508;
assign a2514 = a1182 & ~a1138;
assign a2516 = ~a1082 & a1072;
assign a2518 = ~a2516 & ~a1136;
assign a2520 = ~a2518 & ~a1176;
assign a2522 = a2520 & ~l112;
assign a2524 = ~a2522 & ~a2514;
assign a2526 = a2524 & a2512;
assign a2528 = a2526 & a2506;
assign a2530 = ~a2528 & a1196;
assign a2532 = a1202 & l222;
assign a2534 = ~a2532 & ~a2530;
assign a2536 = ~a2534 & l86;
assign a2538 = l246 & ~l86;
assign a2540 = ~a2538 & ~a2536;
assign a2542 = ~a2540 & a1024;
assign a2544 = ~a1024 & l222;
assign a2546 = ~a2544 & ~a2542;
assign a2548 = a2512 & a1740;
assign a2550 = a1128 & ~l94;
assign a2552 = a2550 & a1726;
assign a2554 = ~a2552 & ~a2520;
assign a2556 = a2554 & ~a2514;
assign a2558 = a2556 & a2548;
assign a2560 = ~a2558 & a1196;
assign a2562 = a1202 & l224;
assign a2564 = ~a2562 & ~a2560;
assign a2566 = ~a2564 & l86;
assign a2568 = l244 & ~l86;
assign a2570 = ~a2568 & ~a2566;
assign a2572 = ~a2570 & a1024;
assign a2574 = ~a1024 & l224;
assign a2576 = ~a2574 & ~a2572;
assign a2578 = l238 & l118;
assign a2580 = a2578 & a1194;
assign a2582 = a2548 & ~a2504;
assign a2584 = ~a2582 & a1196;
assign a2586 = ~a2584 & ~a2580;
assign a2588 = a1202 & l226;
assign a2590 = ~a2588 & a2586;
assign a2592 = ~a2590 & l86;
assign a2594 = l240 & ~l86;
assign a2596 = ~a2594 & ~a2592;
assign a2598 = ~a2596 & a1024;
assign a2600 = ~a1024 & l226;
assign a2602 = ~a2600 & ~a2598;
assign a2604 = ~a1176 & a1160;
assign a2606 = a2604 & a1196;
assign a2608 = a1202 & l228;
assign a2610 = ~a2608 & ~a2606;
assign a2612 = ~a2610 & l86;
assign a2614 = l236 & ~l86;
assign a2616 = ~a2614 & ~a2612;
assign a2618 = ~a2616 & a1024;
assign a2620 = ~a1024 & l228;
assign a2622 = ~a2620 & ~a2618;
assign a2624 = l230 & ~l156;
assign a2626 = ~a2624 & ~l114;
assign a2628 = ~a2626 & l86;
assign a2630 = l234 & ~l86;
assign a2632 = ~a2630 & ~a2628;
assign a2634 = ~a2632 & a1024;
assign a2636 = ~a1024 & l230;
assign a2638 = ~a2636 & ~a2634;
assign a2640 = l86 & i16;
assign a2642 = l242 & ~l86;
assign a2644 = ~a2642 & ~a2640;
assign a2646 = ~a2644 & a1024;
assign a2648 = ~a1024 & l238;
assign a2650 = ~a2648 & ~a2646;
assign a2652 = ~l258 & l256;
assign a2654 = ~a2652 & ~l276;
assign a2656 = ~a2654 & l86;
assign a2658 = l278 & ~l86;
assign a2660 = ~a2658 & ~a2656;
assign a2662 = ~a2660 & a1024;
assign a2664 = ~a1024 & l256;
assign a2666 = ~a2664 & ~a2662;
assign a2668 = l86 & i24;
assign a2670 = l274 & ~l86;
assign a2672 = ~a2670 & ~a2668;
assign a2674 = ~a2672 & a1024;
assign a2676 = ~a1024 & l258;
assign a2678 = ~a2676 & ~a2674;
assign a2680 = ~a1118 & l114;
assign a2682 = ~a2130 & l196;
assign a2684 = ~a2682 & ~a2680;
assign a2686 = ~a2684 & l86;
assign a2688 = l272 & ~l86;
assign a2690 = ~a2688 & ~a2686;
assign a2692 = ~a2690 & a1024;
assign a2694 = ~a1024 & l260;
assign a2696 = ~a2694 & ~a2692;
assign a2698 = a1020 & i22;
assign a2700 = ~a1020 & l262;
assign a2702 = ~a2700 & ~a2698;
assign a2704 = ~a2702 & l86;
assign a2706 = l270 & ~l86;
assign a2708 = ~a2706 & ~a2704;
assign a2710 = ~a2708 & a1252;
assign a2712 = ~a1252 & l262;
assign a2714 = ~a2712 & ~a2710;
assign a2716 = a1020 & i20;
assign a2718 = ~a1020 & l264;
assign a2720 = ~a2718 & ~a2716;
assign a2722 = ~a2720 & l86;
assign a2724 = l268 & ~l86;
assign a2726 = ~a2724 & ~a2722;
assign a2728 = ~a2726 & a1252;
assign a2730 = ~a1252 & l264;
assign a2732 = ~a2730 & ~a2728;
assign a2734 = l260 & l86;
assign a2736 = a2734 & ~a2138;
assign a2738 = l280 & ~l86;
assign a2740 = ~a2738 & ~a2736;
assign a2742 = ~a2740 & a1024;
assign a2744 = ~a1024 & l276;
assign a2746 = ~a2744 & ~a2742;
assign a2748 = ~a2096 & l86;
assign a2750 = l316 & ~l86;
assign a2752 = ~a2750 & ~a2748;
assign a2754 = ~a2752 & a1024;
assign a2756 = ~a1024 & l284;
assign a2758 = ~a2756 & ~a2754;
assign a2760 = ~l288 & l286;
assign a2762 = ~a2760 & ~l306;
assign a2764 = ~a2762 & l86;
assign a2766 = l308 & ~l86;
assign a2768 = ~a2766 & ~a2764;
assign a2770 = ~a2768 & a1024;
assign a2772 = ~a1024 & l286;
assign a2774 = ~a2772 & ~a2770;
assign a2776 = l86 & i28;
assign a2778 = l304 & ~l86;
assign a2780 = ~a2778 & ~a2776;
assign a2782 = ~a2780 & a1024;
assign a2784 = ~a1024 & l288;
assign a2786 = ~a2784 & ~a2782;
assign a2788 = a1620 & l130;
assign a2790 = ~a1672 & l114;
assign a2792 = ~a2790 & ~a2788;
assign a2794 = a1192 & a1190;
assign a2796 = ~l212 & ~l208;
assign a2798 = ~a2796 & l196;
assign a2800 = a2798 & l296;
assign a2802 = l290 & ~l156;
assign a2804 = a2416 & l206;
assign a2806 = ~a2804 & ~a2802;
assign a2808 = a2806 & ~a2800;
assign a2810 = a2808 & ~a2794;
assign a2812 = a2810 & a2792;
assign a2814 = ~a2812 & l86;
assign a2816 = l298 & ~l86;
assign a2818 = ~a2816 & ~a2814;
assign a2820 = ~a2818 & a1024;
assign a2822 = ~a1024 & l290;
assign a2824 = ~a2822 & ~a2820;
assign a2826 = l86 & i26;
assign a2828 = l302 & ~l86;
assign a2830 = ~a2828 & ~a2826;
assign a2832 = ~a2830 & a1024;
assign a2834 = ~a1024 & l294;
assign a2836 = ~a2834 & ~a2832;
assign a2838 = ~a2798 & l296;
assign a2840 = ~a2838 & a2060;
assign a2842 = ~a2840 & l86;
assign a2844 = l300 & ~l86;
assign a2846 = ~a2844 & ~a2842;
assign a2848 = ~a2846 & a1024;
assign a2850 = ~a1024 & l296;
assign a2852 = ~a2850 & ~a2848;
assign a2854 = ~l296 & ~l290;
assign a2856 = ~a2854 & a2152;
assign a2858 = l310 & l86;
assign a2860 = a2858 & a2856;
assign a2862 = l312 & ~l86;
assign a2864 = ~a2862 & ~a2860;
assign a2866 = ~a2864 & a1024;
assign a2868 = ~a1024 & l306;
assign a2870 = ~a2868 & ~a2866;
assign a2872 = ~a2856 & l310;
assign a2874 = a2062 & l284;
assign a2876 = ~a2090 & l114;
assign a2878 = ~a2876 & ~a2874;
assign a2880 = a2878 & ~a2872;
assign a2882 = ~a2880 & l86;
assign a2884 = l314 & ~l86;
assign a2886 = ~a2884 & ~a2882;
assign a2888 = ~a2886 & a1024;
assign a2890 = ~a1024 & l310;
assign a2892 = ~a2890 & ~a2888;
assign a2894 = ~a1846 & ~l136;
assign a2896 = a2894 & l334;
assign a2898 = l334 & ~l140;
assign a2900 = l346 & ~l140;
assign a2902 = l348 & ~l140;
assign a2904 = ~a2902 & ~a2900;
assign a2906 = a2904 & ~a2898;
assign a2908 = ~a2904 & a2898;
assign a2910 = ~a2908 & ~a2906;
assign a2912 = ~a2910 & ~a2894;
assign a2914 = ~a2912 & ~a2896;
assign a2916 = ~a2914 & l86;
assign a2918 = l370 & ~l86;
assign a2920 = ~a2918 & ~a2916;
assign a2922 = ~a2920 & a1024;
assign a2924 = ~a1024 & l334;
assign a2926 = ~a2924 & ~a2922;
assign a2928 = a2894 & l336;
assign a2930 = l350 & ~l140;
assign a2932 = ~a2930 & a2906;
assign a2934 = l336 & ~l140;
assign a2936 = ~a2934 & a2932;
assign a2938 = a2934 & ~a2932;
assign a2940 = ~a2938 & ~a2936;
assign a2942 = ~a2940 & ~a2894;
assign a2944 = ~a2942 & ~a2928;
assign a2946 = ~a2944 & l86;
assign a2948 = l368 & ~l86;
assign a2950 = ~a2948 & ~a2946;
assign a2952 = ~a2950 & a1024;
assign a2954 = ~a1024 & l336;
assign a2956 = ~a2954 & ~a2952;
assign a2958 = a2894 & l338;
assign a2960 = l338 & ~l140;
assign a2962 = ~a2960 & a2936;
assign a2964 = a2960 & ~a2936;
assign a2966 = ~a2964 & ~a2962;
assign a2968 = ~a2966 & ~a2894;
assign a2970 = ~a2968 & ~a2958;
assign a2972 = ~a2970 & l86;
assign a2974 = l366 & ~l86;
assign a2976 = ~a2974 & ~a2972;
assign a2978 = ~a2976 & a1024;
assign a2980 = ~a1024 & l338;
assign a2982 = ~a2980 & ~a2978;
assign a2984 = a2894 & l340;
assign a2986 = l340 & ~l140;
assign a2988 = ~a2986 & a2962;
assign a2990 = a2986 & ~a2962;
assign a2992 = ~a2990 & ~a2988;
assign a2994 = ~a2992 & ~a2894;
assign a2996 = ~a2994 & ~a2984;
assign a2998 = ~a2996 & l86;
assign a3000 = l364 & ~l86;
assign a3002 = ~a3000 & ~a2998;
assign a3004 = ~a3002 & a1024;
assign a3006 = ~a1024 & l340;
assign a3008 = ~a3006 & ~a3004;
assign a3010 = a2894 & l342;
assign a3012 = l344 & ~l140;
assign a3014 = ~a3012 & a2988;
assign a3016 = l342 & ~l140;
assign a3018 = a3016 & ~a3014;
assign a3020 = ~a3016 & a3014;
assign a3022 = ~a3020 & ~a3018;
assign a3024 = ~a3022 & ~a2894;
assign a3026 = ~a3024 & ~a3010;
assign a3028 = ~a3026 & l86;
assign a3030 = l362 & ~l86;
assign a3032 = ~a3030 & ~a3028;
assign a3034 = ~a3032 & a1024;
assign a3036 = ~a1024 & l342;
assign a3038 = ~a3036 & ~a3034;
assign a3040 = a2894 & l344;
assign a3042 = a3012 & ~a2988;
assign a3044 = ~a3042 & ~a3014;
assign a3046 = ~a3044 & ~a2894;
assign a3048 = ~a3046 & ~a3040;
assign a3050 = ~a3048 & l86;
assign a3052 = l360 & ~l86;
assign a3054 = ~a3052 & ~a3050;
assign a3056 = ~a3054 & a1024;
assign a3058 = ~a1024 & l344;
assign a3060 = ~a3058 & ~a3056;
assign a3062 = a2894 & l346;
assign a3064 = a2900 & l348;
assign a3066 = ~a3064 & ~a2904;
assign a3068 = ~a3066 & ~a2894;
assign a3070 = ~a3068 & ~a3062;
assign a3072 = ~a3070 & l86;
assign a3074 = l358 & ~l86;
assign a3076 = ~a3074 & ~a3072;
assign a3078 = ~a3076 & a1024;
assign a3080 = ~a1024 & l346;
assign a3082 = ~a3080 & ~a3078;
assign a3084 = a2894 & l348;
assign a3086 = ~a2902 & ~a2894;
assign a3088 = ~a3086 & ~a3084;
assign a3090 = ~a3088 & l86;
assign a3092 = l356 & ~l86;
assign a3094 = ~a3092 & ~a3090;
assign a3096 = ~a3094 & a1024;
assign a3098 = ~a1024 & l348;
assign a3100 = ~a3098 & ~a3096;
assign a3102 = a2894 & l350;
assign a3104 = a2930 & ~a2906;
assign a3106 = ~a3104 & ~a2932;
assign a3108 = ~a3106 & ~a2894;
assign a3110 = ~a3108 & ~a3102;
assign a3112 = ~a3110 & l86;
assign a3114 = l354 & ~l86;
assign a3116 = ~a3114 & ~a3112;
assign a3118 = ~a3116 & a1024;
assign a3120 = ~a1024 & l350;
assign a3122 = ~a3120 & ~a3118;
assign a3124 = l384 & l86;
assign a3126 = l386 & ~l86;
assign a3128 = ~a3126 & ~a3124;
assign a3130 = ~a3128 & a1024;
assign a3132 = ~a1024 & l380;
assign a3134 = ~a3132 & ~a3130;
assign a3136 = l388 & l86;
assign a3138 = l390 & ~l86;
assign a3140 = ~a3138 & ~a3136;
assign a3142 = ~a3140 & a1024;
assign a3144 = ~a1024 & l384;
assign a3146 = ~a3144 & ~a3142;
assign a3148 = l392 & l86;
assign a3150 = l394 & ~l86;
assign a3152 = ~a3150 & ~a3148;
assign a3154 = ~a3152 & a1024;
assign a3156 = ~a1024 & l388;
assign a3158 = ~a3156 & ~a3154;
assign a3160 = l396 & l86;
assign a3162 = l398 & ~l86;
assign a3164 = ~a3162 & ~a3160;
assign a3166 = ~a3164 & a1024;
assign a3168 = ~a1024 & l392;
assign a3170 = ~a3168 & ~a3166;
assign a3172 = l400 & l86;
assign a3174 = l402 & ~l86;
assign a3176 = ~a3174 & ~a3172;
assign a3178 = ~a3176 & a1024;
assign a3180 = ~a1024 & l396;
assign a3182 = ~a3180 & ~a3178;
assign a3184 = l404 & l86;
assign a3186 = l406 & ~l86;
assign a3188 = ~a3186 & ~a3184;
assign a3190 = ~a3188 & a1024;
assign a3192 = ~a1024 & l400;
assign a3194 = ~a3192 & ~a3190;
assign a3196 = ~a2398 & ~l408;
assign a3198 = ~a3196 & l86;
assign a3200 = l410 & ~l86;
assign a3202 = ~a3200 & ~a3198;
assign a3204 = ~a3202 & a1024;
assign a3206 = ~a1024 & l404;
assign a3208 = ~a3206 & ~a3204;
assign a3210 = l412 & l86;
assign a3212 = l414 & ~l86;
assign a3214 = ~a3212 & ~a3210;
assign a3216 = ~a3214 & a1024;
assign a3218 = ~a1024 & l408;
assign a3220 = ~a3218 & ~a3216;
assign a3222 = l416 & l86;
assign a3224 = l418 & ~l86;
assign a3226 = ~a3224 & ~a3222;
assign a3228 = ~a3226 & a1024;
assign a3230 = ~a1024 & l412;
assign a3232 = ~a3230 & ~a3228;
assign a3234 = l420 & l86;
assign a3236 = l422 & ~l86;
assign a3238 = ~a3236 & ~a3234;
assign a3240 = ~a3238 & a1024;
assign a3242 = ~a1024 & l416;
assign a3244 = ~a3242 & ~a3240;
assign a3246 = a1650 & l86;
assign a3248 = l424 & ~l86;
assign a3250 = ~a3248 & ~a3246;
assign a3252 = ~a3250 & a1024;
assign a3254 = ~a1024 & l420;
assign a3256 = ~a3254 & ~a3252;
assign a3258 = ~l468 & ~l86;
assign a3260 = ~a3258 & a1024;
assign a3262 = ~a1024 & l466;
assign a3264 = ~a3262 & ~a3260;
assign a3266 = ~l816 & ~l86;
assign a3268 = l610 & l536;
assign a3270 = ~a3268 & l86;
assign a3272 = ~a828 & l818;
assign a3274 = a3272 & a3270;
assign a3278 = a3276 & a832;
assign a3280 = ~a832 & l470;
assign a3282 = ~a3280 & ~a3278;
assign a3284 = a828 & i74;
assign a3286 = ~a828 & l472;
assign a3288 = ~a3286 & ~a3284;
assign a3290 = ~a3288 & l86;
assign a3292 = l814 & ~l86;
assign a3294 = ~a3292 & ~a3290;
assign a3296 = ~a3294 & a1252;
assign a3298 = ~a1252 & l472;
assign a3300 = ~a3298 & ~a3296;
assign a3302 = a828 & i72;
assign a3304 = ~a828 & l474;
assign a3306 = ~a3304 & ~a3302;
assign a3308 = ~a3306 & l86;
assign a3310 = l812 & ~l86;
assign a3312 = ~a3310 & ~a3308;
assign a3314 = ~a3312 & a1252;
assign a3316 = ~a1252 & l474;
assign a3318 = ~a3316 & ~a3314;
assign a3320 = a828 & i70;
assign a3322 = ~a828 & l476;
assign a3324 = ~a3322 & ~a3320;
assign a3326 = ~a3324 & l86;
assign a3328 = l810 & ~l86;
assign a3330 = ~a3328 & ~a3326;
assign a3332 = ~a3330 & a1252;
assign a3334 = ~a1252 & l476;
assign a3336 = ~a3334 & ~a3332;
assign a3338 = a828 & i68;
assign a3340 = ~a828 & l478;
assign a3342 = ~a3340 & ~a3338;
assign a3344 = ~a3342 & l86;
assign a3346 = l808 & ~l86;
assign a3348 = ~a3346 & ~a3344;
assign a3350 = ~a3348 & a1252;
assign a3352 = ~a1252 & l478;
assign a3354 = ~a3352 & ~a3350;
assign a3356 = a1334 & a828;
assign a3358 = ~a828 & l480;
assign a3360 = ~a3358 & ~a3356;
assign a3362 = ~a3360 & l86;
assign a3364 = l806 & ~l86;
assign a3366 = ~a3364 & ~a3362;
assign a3368 = ~a3366 & a1252;
assign a3370 = ~a1252 & l480;
assign a3372 = ~a3370 & ~a3368;
assign a3374 = a828 & i64;
assign a3376 = ~a828 & l482;
assign a3378 = ~a3376 & ~a3374;
assign a3380 = ~a3378 & l86;
assign a3382 = l804 & ~l86;
assign a3384 = ~a3382 & ~a3380;
assign a3386 = ~a3384 & a1252;
assign a3388 = ~a1252 & l482;
assign a3390 = ~a3388 & ~a3386;
assign a3392 = a828 & i62;
assign a3394 = ~a828 & l484;
assign a3396 = ~a3394 & ~a3392;
assign a3398 = ~a3396 & l86;
assign a3400 = l802 & ~l86;
assign a3402 = ~a3400 & ~a3398;
assign a3404 = ~a3402 & a1252;
assign a3406 = ~a1252 & l484;
assign a3408 = ~a3406 & ~a3404;
assign a3410 = a828 & i60;
assign a3412 = ~a828 & l486;
assign a3414 = ~a3412 & ~a3410;
assign a3416 = ~a3414 & l86;
assign a3418 = l800 & ~l86;
assign a3420 = ~a3418 & ~a3416;
assign a3422 = ~a3420 & a1252;
assign a3424 = ~a1252 & l486;
assign a3426 = ~a3424 & ~a3422;
assign a3428 = a828 & i58;
assign a3430 = ~a828 & l488;
assign a3432 = ~a3430 & ~a3428;
assign a3434 = ~a3432 & l86;
assign a3436 = l798 & ~l86;
assign a3438 = ~a3436 & ~a3434;
assign a3440 = ~a3438 & a1252;
assign a3442 = ~a1252 & l488;
assign a3444 = ~a3442 & ~a3440;
assign a3446 = a828 & i56;
assign a3448 = ~a828 & l490;
assign a3450 = ~a3448 & ~a3446;
assign a3452 = ~a3450 & l86;
assign a3454 = l796 & ~l86;
assign a3456 = ~a3454 & ~a3452;
assign a3458 = ~a3456 & a1252;
assign a3460 = ~a1252 & l490;
assign a3462 = ~a3460 & ~a3458;
assign a3464 = a828 & i52;
assign a3466 = ~a828 & l492;
assign a3468 = ~a3466 & ~a3464;
assign a3470 = ~a3468 & l86;
assign a3472 = l794 & ~l86;
assign a3474 = ~a3472 & ~a3470;
assign a3476 = ~a3474 & a1252;
assign a3478 = ~a1252 & l492;
assign a3480 = ~a3478 & ~a3476;
assign a3482 = a828 & i50;
assign a3484 = ~a828 & l494;
assign a3486 = ~a3484 & ~a3482;
assign a3488 = ~a3486 & l86;
assign a3490 = l792 & ~l86;
assign a3492 = ~a3490 & ~a3488;
assign a3494 = ~a3492 & a1252;
assign a3496 = ~a1252 & l494;
assign a3498 = ~a3496 & ~a3494;
assign a3500 = ~a832 & l496;
assign a3502 = ~a3500 & ~a1504;
assign a3504 = a828 & i48;
assign a3506 = ~a828 & l498;
assign a3508 = ~a3506 & ~a3504;
assign a3510 = ~a3508 & l86;
assign a3512 = l790 & ~l86;
assign a3514 = ~a3512 & ~a3510;
assign a3516 = ~a3514 & a1252;
assign a3518 = ~a1252 & l498;
assign a3520 = ~a3518 & ~a3516;
assign a3522 = ~a1532 & a832;
assign a3524 = ~a832 & l500;
assign a3526 = ~a3524 & ~a3522;
assign a3528 = ~a1544 & a832;
assign a3530 = ~a832 & l502;
assign a3532 = ~a3530 & ~a3528;
assign a3534 = ~a1556 & a832;
assign a3536 = ~a832 & l504;
assign a3538 = ~a3536 & ~a3534;
assign a3540 = l744 & l86;
assign a3542 = l746 & ~l86;
assign a3544 = ~a3542 & ~a3540;
assign a3546 = ~a3544 & a832;
assign a3548 = ~a832 & l506;
assign a3550 = ~a3548 & ~a3546;
assign a3552 = ~l522 & ~l520;
assign a3554 = a3552 & ~l518;
assign a3556 = ~a3554 & ~l516;
assign a3558 = ~l530 & ~l528;
assign a3560 = a3558 & l526;
assign a3562 = a3560 & ~l524;
assign a3564 = l532 & l524;
assign a3566 = a3558 & ~l526;
assign a3568 = a3566 & a3564;
assign a3570 = ~a3568 & ~a3562;
assign a3572 = ~a3570 & a970;
assign a3574 = ~l532 & l524;
assign a3576 = ~l530 & l528;
assign a3578 = a3576 & ~l526;
assign a3580 = ~a3578 & ~a3560;
assign a3582 = ~a3580 & a3574;
assign a3584 = a3582 & ~a968;
assign a3586 = ~a3584 & ~a3572;
assign a3588 = a3586 & a3556;
assign a3590 = ~a970 & a968;
assign a3592 = ~a3590 & a936;
assign a3594 = a3592 & a3588;
assign a3596 = a3594 & l514;
assign a3598 = a3596 & l534;
assign a3600 = ~l536 & l512;
assign a3602 = l540 & l538;
assign a3604 = ~a3602 & ~a3600;
assign a3606 = a944 & l478;
assign a3608 = ~a3606 & a954;
assign a3610 = ~a3608 & a982;
assign a3612 = a3610 & l496;
assign a3614 = ~a3612 & a3604;
assign a3616 = a3614 & ~a3598;
assign a3618 = a3616 & ~l512;
assign a3620 = ~a3596 & l542;
assign a3622 = a3620 & ~a3618;
assign a3624 = l508 & ~l506;
assign a3626 = ~a3624 & ~a3622;
assign a3628 = ~a3626 & l86;
assign a3630 = l544 & ~l86;
assign a3632 = ~a3630 & ~a3628;
assign a3634 = ~a3632 & a832;
assign a3636 = ~a832 & l508;
assign a3638 = ~a3636 & ~a3634;
assign a3640 = ~a3616 & l86;
assign a3642 = l742 & ~l86;
assign a3644 = ~a3642 & ~a3640;
assign a3646 = ~a3644 & a832;
assign a3648 = ~a832 & l512;
assign a3650 = ~a3648 & ~a3646;
assign a3652 = ~a982 & l496;
assign a3654 = ~a3586 & a3556;
assign a3656 = ~a3654 & a3592;
assign a3658 = a3656 & l514;
assign a3660 = a3658 & ~a3594;
assign a3662 = ~a3660 & ~a3652;
assign a3664 = ~a3662 & l86;
assign a3666 = l740 & ~l86;
assign a3668 = ~a3666 & ~a3664;
assign a3670 = ~a3668 & a832;
assign a3672 = ~a832 & l514;
assign a3674 = ~a3672 & ~a3670;
assign a3676 = a3576 & l526;
assign a3678 = l494 & l472;
assign a3680 = a3678 & ~a916;
assign a3682 = ~a968 & l478;
assign a3684 = a3682 & a944;
assign a3686 = a936 & l476;
assign a3688 = ~a3686 & ~a878;
assign a3690 = ~a3688 & a3682;
assign a3692 = a3690 & l494;
assign a3694 = ~a3692 & ~a3684;
assign a3696 = a3694 & ~a3680;
assign a3698 = ~a3696 & l562;
assign a3700 = ~a3606 & ~a860;
assign a3702 = ~a3700 & ~l562;
assign a3704 = ~a3702 & ~a3698;
assign a3706 = a3704 & l532;
assign a3708 = ~a3706 & ~l524;
assign a3710 = ~a3708 & ~a3564;
assign a3712 = a3710 & a3676;
assign a3714 = a3712 & a3556;
assign a3716 = a3714 & l564;
assign a3718 = a3716 & l522;
assign a3720 = l582 & ~l536;
assign a3722 = l584 & i10;
assign a3724 = ~a3722 & ~a3720;
assign a3726 = a982 & l496;
assign a3728 = ~a3726 & a3724;
assign a3730 = a3728 & ~a3596;
assign a3732 = a3730 & ~l582;
assign a3734 = ~a3732 & l520;
assign a3736 = a3734 & l580;
assign a3738 = l586 & l562;
assign a3740 = a3738 & a3736;
assign a3742 = l516 & i30;
assign a3744 = ~l568 & ~l554;
assign a3746 = a3744 & ~l592;
assign a3748 = a3746 & ~l576;
assign a3750 = ~a3748 & ~l564;
assign a3752 = ~a3750 & a3742;
assign a3754 = ~a3752 & l516;
assign a3756 = l490 & l474;
assign a3758 = ~a3756 & a900;
assign a3760 = ~a3758 & ~a906;
assign a3762 = ~a3760 & l472;
assign a3764 = ~a3762 & a968;
assign a3766 = a3764 & a956;
assign a3768 = ~a3766 & l496;
assign a3770 = ~a3768 & ~a3754;
assign a3772 = a3770 & ~a3740;
assign a3774 = a3772 & ~a3718;
assign a3776 = ~a3774 & l86;
assign a3778 = l738 & ~l86;
assign a3780 = ~a3778 & ~a3776;
assign a3782 = ~a3780 & a832;
assign a3784 = ~a832 & l516;
assign a3786 = ~a3784 & ~a3782;
assign a3788 = ~a3716 & l522;
assign a3790 = ~l700 & ~l698;
assign a3792 = ~l704 & ~l702;
assign a3794 = a3792 & a3790;
assign a3796 = ~l708 & ~l706;
assign a3798 = ~l712 & ~l710;
assign a3800 = a3798 & ~l714;
assign a3802 = a3800 & a3796;
assign a3804 = a3802 & a3794;
assign a3806 = ~a3804 & l518;
assign a3808 = ~a3806 & ~a3788;
assign a3810 = ~a3808 & l86;
assign a3812 = l736 & ~l86;
assign a3814 = ~a3812 & ~a3810;
assign a3816 = ~a3814 & a832;
assign a3818 = ~a832 & l518;
assign a3820 = ~a3818 & ~a3816;
assign a3822 = ~a3740 & ~l536;
assign a3824 = a3822 & l520;
assign a3826 = a3804 & l518;
assign a3828 = a3766 & l496;
assign a3830 = ~a3828 & ~a3826;
assign a3832 = a3830 & ~a3824;
assign a3834 = ~a3832 & l86;
assign a3836 = l716 & ~l86;
assign a3838 = ~a3836 & ~a3834;
assign a3840 = ~a3838 & a832;
assign a3842 = ~a832 & l520;
assign a3844 = ~a3842 & ~a3840;
assign a3846 = a3752 & l86;
assign a3848 = l696 & ~l86;
assign a3850 = ~a3848 & ~a3846;
assign a3852 = ~a3850 & a832;
assign a3854 = ~a832 & l522;
assign a3856 = ~a3854 & ~a3852;
assign a3858 = a3752 & i40;
assign a3860 = ~a3752 & l524;
assign a3862 = ~a3860 & ~a3858;
assign a3864 = ~a3862 & l86;
assign a3866 = l694 & ~l86;
assign a3868 = ~a3866 & ~a3864;
assign a3870 = ~a3868 & a832;
assign a3872 = ~a832 & l524;
assign a3874 = ~a3872 & ~a3870;
assign a3876 = a3752 & i38;
assign a3878 = ~a3752 & l526;
assign a3880 = ~a3878 & ~a3876;
assign a3882 = ~a3880 & l86;
assign a3884 = l692 & ~l86;
assign a3886 = ~a3884 & ~a3882;
assign a3888 = ~a3886 & a832;
assign a3890 = ~a832 & l526;
assign a3892 = ~a3890 & ~a3888;
assign a3894 = a3752 & i36;
assign a3896 = ~a3752 & l528;
assign a3898 = ~a3896 & ~a3894;
assign a3900 = ~a3898 & l86;
assign a3902 = l690 & ~l86;
assign a3904 = ~a3902 & ~a3900;
assign a3906 = ~a3904 & a832;
assign a3908 = ~a832 & l528;
assign a3910 = ~a3908 & ~a3906;
assign a3912 = a3752 & i34;
assign a3914 = ~a3752 & l530;
assign a3916 = ~a3914 & ~a3912;
assign a3918 = ~a3916 & l86;
assign a3920 = l688 & ~l86;
assign a3922 = ~a3920 & ~a3918;
assign a3924 = ~a3922 & a832;
assign a3926 = ~a832 & l530;
assign a3928 = ~a3926 & ~a3924;
assign a3930 = a3752 & i32;
assign a3932 = ~a3752 & l532;
assign a3934 = ~a3932 & ~a3930;
assign a3936 = ~a3934 & l86;
assign a3938 = l686 & ~l86;
assign a3940 = ~a3938 & ~a3936;
assign a3942 = ~a3940 & a832;
assign a3944 = ~a832 & l532;
assign a3946 = ~a3944 & ~a3942;
assign a3948 = ~a3610 & l84;
assign a3950 = ~l556 & ~l554;
assign a3952 = a3950 & l534;
assign a3954 = a3952 & ~a3596;
assign a3956 = ~a3954 & ~a3948;
assign a3958 = ~a3956 & l86;
assign a3960 = l684 & ~l86;
assign a3962 = ~a3960 & ~a3958;
assign a3964 = ~a3962 & a832;
assign a3966 = ~a832 & l534;
assign a3968 = ~a3966 & ~a3964;
assign a3970 = ~a968 & a936;
assign a3972 = l494 & l476;
assign a3974 = ~a3972 & a3970;
assign a3976 = a976 & a962;
assign a3978 = ~a3976 & ~a3974;
assign a3980 = l598 & l586;
assign a3982 = a3980 & a3736;
assign a3984 = ~a3982 & ~a3740;
assign a3986 = ~a3984 & ~a3978;
assign a3988 = l656 & ~l536;
assign a3990 = a3988 & ~a3986;
assign a3992 = l660 & l658;
assign a3994 = a3972 & a936;
assign a3996 = ~a3994 & ~a876;
assign a3998 = a974 & ~a966;
assign a4000 = ~a3998 & a3996;
assign a4002 = ~a4000 & ~a968;
assign a4004 = a950 & a910;
assign a4006 = a4004 & a874;
assign a4008 = a4006 & ~a4002;
assign a4010 = a4008 & l496;
assign a4012 = ~a4010 & ~a3992;
assign a4014 = a4012 & ~a3990;
assign a4016 = a4014 & ~l656;
assign a4018 = l662 & l86;
assign a4020 = a4018 & a3734;
assign a4022 = a4020 & ~a4016;
assign a4024 = a3556 & l564;
assign a4026 = a4024 & ~a3712;
assign a4028 = a4026 & ~a3704;
assign a4030 = a3822 & l588;
assign a4032 = l592 & i14;
assign a4034 = a956 & l496;
assign a4036 = ~a4034 & ~a4032;
assign a4038 = a4036 & ~a4030;
assign a4040 = a4038 & ~a4028;
assign a4042 = a4040 & ~l588;
assign a4044 = ~a3704 & a3680;
assign a4046 = ~a4044 & a3740;
assign a4048 = ~a4046 & ~a3982;
assign a4050 = l580 & ~l536;
assign a4052 = a4050 & a4048;
assign a4054 = l632 & l630;
assign a4056 = ~l638 & ~l636;
assign a4058 = a4056 & l634;
assign a4060 = ~a4058 & ~a4054;
assign a4062 = a926 & l496;
assign a4064 = ~a4062 & a4060;
assign a4066 = a4064 & ~a4052;
assign a4068 = a4066 & ~l580;
assign a4070 = ~a4068 & ~a3618;
assign a4072 = a4070 & ~a4042;
assign a4074 = a4072 & a4022;
assign a4076 = l664 & ~l86;
assign a4078 = ~a4076 & ~a4074;
assign a4080 = ~a4078 & a832;
assign a4082 = ~a832 & l536;
assign a4084 = ~a4082 & ~a4080;
assign a4086 = ~l540 & l538;
assign a4088 = ~a4086 & ~l550;
assign a4090 = ~a4088 & l86;
assign a4092 = l552 & ~l86;
assign a4094 = ~a4092 & ~a4090;
assign a4096 = ~a4094 & a832;
assign a4098 = ~a832 & l538;
assign a4100 = ~a4098 & ~a4096;
assign a4102 = ~a2188 & a832;
assign a4104 = ~a832 & l540;
assign a4106 = ~a4104 & ~a4102;
assign a4108 = ~a3610 & l546;
assign a4110 = a4108 & l496;
assign a4112 = a3620 & a3618;
assign a4114 = ~a4112 & ~a4110;
assign a4116 = ~a4114 & l86;
assign a4118 = l548 & ~l86;
assign a4120 = ~a4118 & ~a4116;
assign a4122 = ~a4120 & a832;
assign a4124 = ~a832 & l542;
assign a4126 = ~a4124 & ~a4122;
assign a4128 = ~a2830 & a832;
assign a4130 = ~a832 & l546;
assign a4132 = ~a4130 & ~a4128;
assign a4134 = l534 & l86;
assign a4136 = a4134 & ~a3950;
assign a4138 = l558 & ~l86;
assign a4140 = ~a4138 & ~a4136;
assign a4142 = ~a4140 & a832;
assign a4144 = ~a832 & l550;
assign a4146 = ~a4144 & ~a4142;
assign a4148 = a3704 & l86;
assign a4150 = a4148 & a4026;
assign a4152 = l566 & ~l86;
assign a4154 = ~a4152 & ~a4150;
assign a4156 = ~a4154 & a832;
assign a4158 = ~a832 & l554;
assign a4160 = ~a4158 & ~a4156;
assign a4162 = l514 & l86;
assign a4164 = a4162 & ~a3656;
assign a4166 = l560 & ~l86;
assign a4168 = ~a4166 & ~a4164;
assign a4170 = ~a4168 & a832;
assign a4172 = ~a832 & l556;
assign a4174 = ~a4172 & ~a4170;
assign a4176 = l606 & l602;
assign a4178 = ~l604 & ~l602;
assign a4180 = ~a4178 & ~l608;
assign a4182 = a4180 & ~a4176;
assign a4184 = a4182 & ~a982;
assign a4186 = ~a4184 & l506;
assign a4188 = ~l562 & ~l506;
assign a4190 = ~a4188 & a3270;
assign a4192 = a4190 & ~a4186;
assign a4194 = l654 & ~l86;
assign a4196 = ~a4194 & ~a4192;
assign a4198 = ~a4196 & a832;
assign a4200 = ~a832 & l562;
assign a4202 = ~a4200 & ~a4198;
assign a4204 = ~l570 & l568;
assign a4206 = ~a3556 & l564;
assign a4208 = ~a4206 & ~a4204;
assign a4210 = ~a4208 & l86;
assign a4212 = l572 & ~l86;
assign a4214 = ~a4212 & ~a4210;
assign a4216 = ~a4214 & a832;
assign a4218 = ~a832 & l564;
assign a4220 = ~a4218 & ~a4216;
assign a4222 = l570 & l568;
assign a4224 = ~a4222 & ~l576;
assign a4226 = a4224 & ~a3716;
assign a4228 = ~a4226 & l86;
assign a4230 = l578 & ~l86;
assign a4232 = ~a4230 & ~a4228;
assign a4234 = ~a4232 & a832;
assign a4236 = ~a832 & l568;
assign a4238 = ~a4236 & ~a4234;
assign a4240 = a3714 & i6;
assign a4242 = ~a4240 & ~l570;
assign a4244 = ~a3714 & i8;
assign a4246 = ~l470 & l86;
assign a4248 = a4246 & ~a4244;
assign a4250 = a4248 & ~a4242;
assign a4252 = l574 & ~l86;
assign a4254 = ~a4252 & ~a4250;
assign a4256 = ~a4254 & a832;
assign a4258 = ~a832 & l570;
assign a4260 = ~a4258 & ~a4256;
assign a4262 = a3740 & l588;
assign a4264 = ~a956 & l496;
assign a4266 = ~a4264 & ~a4262;
assign a4268 = ~a4266 & l86;
assign a4270 = l590 & ~l86;
assign a4272 = ~a4270 & ~a4268;
assign a4274 = ~a4272 & a832;
assign a4276 = ~a832 & l576;
assign a4278 = ~a4276 & ~a4274;
assign a4280 = ~a4066 & l86;
assign a4282 = l640 & ~l86;
assign a4284 = ~a4282 & ~a4280;
assign a4286 = ~a4284 & a832;
assign a4288 = ~a832 & l580;
assign a4290 = ~a4288 & ~a4286;
assign a4292 = ~a3730 & l86;
assign a4294 = l628 & ~l86;
assign a4296 = ~a4294 & ~a4292;
assign a4298 = ~a4296 & a832;
assign a4300 = ~a832 & l582;
assign a4302 = ~a4300 & ~a4298;
assign a4304 = l584 & ~i10;
assign a4306 = ~a4304 & ~l556;
assign a4308 = ~a4306 & l86;
assign a4310 = l626 & ~l86;
assign a4312 = ~a4310 & ~a4308;
assign a4314 = ~a4312 & a832;
assign a4316 = ~a832 & l584;
assign a4318 = ~a4316 & ~a4314;
assign a4320 = ~l598 & ~l562;
assign a4322 = ~a4320 & l586;
assign a4324 = a4322 & ~a3736;
assign a4326 = ~a4324 & ~a994;
assign a4328 = ~a4326 & l86;
assign a4330 = l600 & ~l86;
assign a4332 = ~a4330 & ~a4328;
assign a4334 = ~a4332 & a832;
assign a4336 = ~a832 & l586;
assign a4338 = ~a4336 & ~a4334;
assign a4340 = ~a4040 & l86;
assign a4342 = l594 & ~l86;
assign a4344 = ~a4342 & ~a4340;
assign a4346 = ~a4344 & a832;
assign a4348 = ~a832 & l588;
assign a4350 = ~a4348 & ~a4346;
assign a4352 = l592 & ~i14;
assign a4354 = ~a4352 & ~l554;
assign a4356 = ~a4354 & l86;
assign a4358 = l596 & ~l86;
assign a4360 = ~a4358 & ~a4356;
assign a4362 = ~a4360 & a832;
assign a4364 = ~a832 & l592;
assign a4366 = ~a4364 & ~a4362;
assign a4368 = l608 & ~l606;
assign a4370 = a4368 & a4178;
assign a4372 = ~l608 & l604;
assign a4374 = a4372 & a4176;
assign a4376 = ~a4374 & ~a4370;
assign a4378 = ~a4376 & ~a982;
assign a4380 = a974 & a962;
assign a4382 = ~a4380 & l506;
assign a4384 = a4382 & ~a4378;
assign a4386 = ~l598 & ~l506;
assign a4388 = ~a4386 & a3270;
assign a4390 = a4388 & ~a4384;
assign a4392 = l612 & ~l86;
assign a4394 = ~a4392 & ~a4390;
assign a4396 = ~a4394 & a832;
assign a4398 = ~a832 & l598;
assign a4400 = ~a4398 & ~a4396;
assign a4402 = ~a890 & a880;
assign a4404 = ~a4402 & ~a942;
assign a4406 = ~a4404 & ~a968;
assign a4408 = a4406 & ~l494;
assign a4410 = ~a4408 & ~a3680;
assign a4412 = ~a834 & ~l494;
assign a4414 = a4412 & ~a916;
assign a4416 = a3690 & ~l494;
assign a4418 = ~a4416 & ~a4414;
assign a4420 = a4418 & a4410;
assign a4422 = ~a4420 & a996;
assign a4424 = a1002 & l602;
assign a4426 = ~a4424 & ~a4422;
assign a4428 = ~a4426 & l86;
assign a4430 = l624 & ~l86;
assign a4432 = ~a4430 & ~a4428;
assign a4434 = ~a4432 & a832;
assign a4436 = ~a832 & l602;
assign a4438 = ~a4436 & ~a4434;
assign a4440 = ~a4416 & a3694;
assign a4442 = ~l478 & ~l476;
assign a4444 = a4442 & a3970;
assign a4446 = ~a4444 & ~a4406;
assign a4448 = a4446 & a4440;
assign a4450 = ~a4448 & a996;
assign a4452 = a1002 & l604;
assign a4454 = ~a4452 & ~a4450;
assign a4456 = ~a4454 & l86;
assign a4458 = l622 & ~l86;
assign a4460 = ~a4458 & ~a4456;
assign a4462 = ~a4460 & a832;
assign a4464 = ~a832 & l604;
assign a4466 = ~a4464 & ~a4462;
assign a4468 = l618 & l500;
assign a4470 = a4468 & a994;
assign a4472 = a4440 & ~a4414;
assign a4474 = ~a4472 & a996;
assign a4476 = ~a4474 & ~a4470;
assign a4478 = a1002 & l606;
assign a4480 = ~a4478 & a4476;
assign a4482 = ~a4480 & l86;
assign a4484 = l620 & ~l86;
assign a4486 = ~a4484 & ~a4482;
assign a4488 = ~a4486 & a832;
assign a4490 = ~a832 & l606;
assign a4492 = ~a4490 & ~a4488;
assign a4494 = a3682 & a972;
assign a4496 = a4494 & a996;
assign a4498 = a1002 & l608;
assign a4500 = ~a4498 & ~a4496;
assign a4502 = ~a4500 & l86;
assign a4504 = l616 & ~l86;
assign a4506 = ~a4504 & ~a4502;
assign a4508 = ~a4506 & a832;
assign a4510 = ~a832 & l608;
assign a4512 = ~a4510 & ~a4508;
assign a4514 = l610 & ~l536;
assign a4516 = ~a4514 & ~l496;
assign a4518 = ~a4516 & l86;
assign a4520 = l614 & ~l86;
assign a4522 = ~a4520 & ~a4518;
assign a4524 = ~a4522 & a832;
assign a4526 = ~a832 & l610;
assign a4528 = ~a4526 & ~a4524;
assign a4530 = ~a2644 & a832;
assign a4532 = ~a832 & l618;
assign a4534 = ~a4532 & ~a4530;
assign a4536 = ~l632 & l630;
assign a4538 = ~a4536 & ~l648;
assign a4540 = ~a4538 & l86;
assign a4542 = l650 & ~l86;
assign a4544 = ~a4542 & ~a4540;
assign a4546 = ~a4544 & a832;
assign a4548 = ~a832 & l630;
assign a4550 = ~a4548 & ~a4546;
assign a4552 = ~a2672 & a832;
assign a4554 = ~a832 & l632;
assign a4556 = ~a4554 & ~a4552;
assign a4558 = ~a926 & l496;
assign a4560 = ~a4048 & l580;
assign a4562 = ~a4560 & ~a4558;
assign a4564 = ~a4562 & l86;
assign a4566 = l646 & ~l86;
assign a4568 = ~a4566 & ~a4564;
assign a4570 = ~a4568 & a832;
assign a4572 = ~a832 & l634;
assign a4574 = ~a4572 & ~a4570;
assign a4576 = a828 & i22;
assign a4578 = ~a828 & l636;
assign a4580 = ~a4578 & ~a4576;
assign a4582 = ~a4580 & l86;
assign a4584 = l644 & ~l86;
assign a4586 = ~a4584 & ~a4582;
assign a4588 = ~a4586 & a1252;
assign a4590 = ~a1252 & l636;
assign a4592 = ~a4590 & ~a4588;
assign a4594 = a828 & i20;
assign a4596 = ~a828 & l638;
assign a4598 = ~a4596 & ~a4594;
assign a4600 = ~a4598 & l86;
assign a4602 = l642 & ~l86;
assign a4604 = ~a4602 & ~a4600;
assign a4606 = ~a4604 & a1252;
assign a4608 = ~a1252 & l638;
assign a4610 = ~a4608 & ~a4606;
assign a4612 = l634 & l86;
assign a4614 = a4612 & ~a4056;
assign a4616 = l652 & ~l86;
assign a4618 = ~a4616 & ~a4614;
assign a4620 = ~a4618 & a832;
assign a4622 = ~a832 & l648;
assign a4624 = ~a4622 & ~a4620;
assign a4626 = ~a4014 & l86;
assign a4628 = l682 & ~l86;
assign a4630 = ~a4628 & ~a4626;
assign a4632 = ~a4630 & a832;
assign a4634 = ~a832 & l656;
assign a4636 = ~a4634 & ~a4632;
assign a4638 = ~l660 & l658;
assign a4640 = ~a4638 & ~l672;
assign a4642 = ~a4640 & l86;
assign a4644 = l674 & ~l86;
assign a4646 = ~a4644 & ~a4642;
assign a4648 = ~a4646 & a832;
assign a4650 = ~a832 & l658;
assign a4652 = ~a4650 & ~a4648;
assign a4654 = ~a2780 & a832;
assign a4656 = ~a832 & l660;
assign a4658 = ~a4656 & ~a4654;
assign a4660 = ~a4108 & l496;
assign a4662 = ~l592 & ~l588;
assign a4664 = ~a4662 & l580;
assign a4666 = a4664 & l666;
assign a4668 = l662 & ~l536;
assign a4670 = a4320 & l586;
assign a4672 = ~a4670 & ~a4668;
assign a4674 = a4672 & ~a4666;
assign a4676 = a4674 & ~a4660;
assign a4678 = a992 & a990;
assign a4680 = a3596 & l542;
assign a4682 = ~a4680 & ~a4678;
assign a4684 = a4682 & a4676;
assign a4686 = ~a4684 & l86;
assign a4688 = l668 & ~l86;
assign a4690 = ~a4688 & ~a4686;
assign a4692 = ~a4690 & a832;
assign a4694 = ~a832 & l662;
assign a4696 = ~a4694 & ~a4692;
assign a4698 = ~a4664 & l666;
assign a4700 = ~a4698 & a3984;
assign a4702 = ~a4700 & l86;
assign a4704 = l670 & ~l86;
assign a4706 = ~a4704 & ~a4702;
assign a4708 = ~a4706 & a832;
assign a4710 = ~a832 & l666;
assign a4712 = ~a4710 & ~a4708;
assign a4714 = ~l666 & ~l662;
assign a4716 = ~a4714 & a4070;
assign a4718 = l676 & l86;
assign a4720 = a4718 & a4716;
assign a4722 = l678 & ~l86;
assign a4724 = ~a4722 & ~a4720;
assign a4726 = ~a4724 & a832;
assign a4728 = ~a832 & l672;
assign a4730 = ~a4728 & ~a4726;
assign a4732 = ~a4716 & l676;
assign a4734 = a3986 & l656;
assign a4736 = ~a4008 & l496;
assign a4738 = ~a4736 & ~a4734;
assign a4740 = a4738 & ~a4732;
assign a4742 = ~a4740 & l86;
assign a4744 = l680 & ~l86;
assign a4746 = ~a4744 & ~a4742;
assign a4748 = ~a4746 & a832;
assign a4750 = ~a832 & l676;
assign a4752 = ~a4750 & ~a4748;
assign a4754 = ~a3788 & ~l518;
assign a4756 = a4754 & l698;
assign a4758 = l698 & ~l522;
assign a4760 = l710 & ~l522;
assign a4762 = l712 & ~l522;
assign a4764 = ~a4762 & ~a4760;
assign a4766 = a4764 & ~a4758;
assign a4768 = ~a4764 & a4758;
assign a4770 = ~a4768 & ~a4766;
assign a4772 = ~a4770 & ~a4754;
assign a4774 = ~a4772 & ~a4756;
assign a4776 = ~a4774 & l86;
assign a4778 = l734 & ~l86;
assign a4780 = ~a4778 & ~a4776;
assign a4782 = ~a4780 & a832;
assign a4784 = ~a832 & l698;
assign a4786 = ~a4784 & ~a4782;
assign a4788 = a4754 & l700;
assign a4790 = l714 & ~l522;
assign a4792 = ~a4790 & a4766;
assign a4794 = l700 & ~l522;
assign a4796 = ~a4794 & a4792;
assign a4798 = a4794 & ~a4792;
assign a4800 = ~a4798 & ~a4796;
assign a4802 = ~a4800 & ~a4754;
assign a4804 = ~a4802 & ~a4788;
assign a4806 = ~a4804 & l86;
assign a4808 = l732 & ~l86;
assign a4810 = ~a4808 & ~a4806;
assign a4812 = ~a4810 & a832;
assign a4814 = ~a832 & l700;
assign a4816 = ~a4814 & ~a4812;
assign a4818 = a4754 & l702;
assign a4820 = l702 & ~l522;
assign a4822 = ~a4820 & a4796;
assign a4824 = a4820 & ~a4796;
assign a4826 = ~a4824 & ~a4822;
assign a4828 = ~a4826 & ~a4754;
assign a4830 = ~a4828 & ~a4818;
assign a4832 = ~a4830 & l86;
assign a4834 = l730 & ~l86;
assign a4836 = ~a4834 & ~a4832;
assign a4838 = ~a4836 & a832;
assign a4840 = ~a832 & l702;
assign a4842 = ~a4840 & ~a4838;
assign a4844 = a4754 & l704;
assign a4846 = l704 & ~l522;
assign a4848 = ~a4846 & a4822;
assign a4850 = a4846 & ~a4822;
assign a4852 = ~a4850 & ~a4848;
assign a4854 = ~a4852 & ~a4754;
assign a4856 = ~a4854 & ~a4844;
assign a4858 = ~a4856 & l86;
assign a4860 = l728 & ~l86;
assign a4862 = ~a4860 & ~a4858;
assign a4864 = ~a4862 & a832;
assign a4866 = ~a832 & l704;
assign a4868 = ~a4866 & ~a4864;
assign a4870 = a4754 & l706;
assign a4872 = l708 & ~l522;
assign a4874 = ~a4872 & a4848;
assign a4876 = l706 & ~l522;
assign a4878 = a4876 & ~a4874;
assign a4880 = ~a4876 & a4874;
assign a4882 = ~a4880 & ~a4878;
assign a4884 = ~a4882 & ~a4754;
assign a4886 = ~a4884 & ~a4870;
assign a4888 = ~a4886 & l86;
assign a4890 = l726 & ~l86;
assign a4892 = ~a4890 & ~a4888;
assign a4894 = ~a4892 & a832;
assign a4896 = ~a832 & l706;
assign a4898 = ~a4896 & ~a4894;
assign a4900 = a4754 & l708;
assign a4902 = a4872 & ~a4848;
assign a4904 = ~a4902 & ~a4874;
assign a4906 = ~a4904 & ~a4754;
assign a4908 = ~a4906 & ~a4900;
assign a4910 = ~a4908 & l86;
assign a4912 = l724 & ~l86;
assign a4914 = ~a4912 & ~a4910;
assign a4916 = ~a4914 & a832;
assign a4918 = ~a832 & l708;
assign a4920 = ~a4918 & ~a4916;
assign a4922 = a4754 & l710;
assign a4924 = a4760 & l712;
assign a4926 = ~a4924 & ~a4764;
assign a4928 = ~a4926 & ~a4754;
assign a4930 = ~a4928 & ~a4922;
assign a4932 = ~a4930 & l86;
assign a4934 = l722 & ~l86;
assign a4936 = ~a4934 & ~a4932;
assign a4938 = ~a4936 & a832;
assign a4940 = ~a832 & l710;
assign a4942 = ~a4940 & ~a4938;
assign a4944 = a4754 & l712;
assign a4946 = ~a4762 & ~a4754;
assign a4948 = ~a4946 & ~a4944;
assign a4950 = ~a4948 & l86;
assign a4952 = l720 & ~l86;
assign a4954 = ~a4952 & ~a4950;
assign a4956 = ~a4954 & a832;
assign a4958 = ~a832 & l712;
assign a4960 = ~a4958 & ~a4956;
assign a4962 = a4754 & l714;
assign a4964 = a4790 & ~a4766;
assign a4966 = ~a4964 & ~a4792;
assign a4968 = ~a4966 & ~a4754;
assign a4970 = ~a4968 & ~a4962;
assign a4972 = ~a4970 & l86;
assign a4974 = l718 & ~l86;
assign a4976 = ~a4974 & ~a4972;
assign a4978 = ~a4976 & a832;
assign a4980 = ~a832 & l714;
assign a4982 = ~a4980 & ~a4978;
assign a4984 = l748 & l86;
assign a4986 = l750 & ~l86;
assign a4988 = ~a4986 & ~a4984;
assign a4990 = ~a4988 & a832;
assign a4992 = ~a832 & l744;
assign a4994 = ~a4992 & ~a4990;
assign a4996 = l752 & l86;
assign a4998 = l754 & ~l86;
assign a5000 = ~a4998 & ~a4996;
assign a5002 = ~a5000 & a832;
assign a5004 = ~a832 & l748;
assign a5006 = ~a5004 & ~a5002;
assign a5008 = l756 & l86;
assign a5010 = l758 & ~l86;
assign a5012 = ~a5010 & ~a5008;
assign a5014 = ~a5012 & a832;
assign a5016 = ~a832 & l752;
assign a5018 = ~a5016 & ~a5014;
assign a5020 = l760 & l86;
assign a5022 = l762 & ~l86;
assign a5024 = ~a5022 & ~a5020;
assign a5026 = ~a5024 & a832;
assign a5028 = ~a832 & l756;
assign a5030 = ~a5028 & ~a5026;
assign a5032 = l764 & l86;
assign a5034 = l766 & ~l86;
assign a5036 = ~a5034 & ~a5032;
assign a5038 = ~a5036 & a832;
assign a5040 = ~a832 & l760;
assign a5042 = ~a5040 & ~a5038;
assign a5044 = l768 & l86;
assign a5046 = l770 & ~l86;
assign a5048 = ~a5046 & ~a5044;
assign a5050 = ~a5048 & a832;
assign a5052 = ~a832 & l764;
assign a5054 = ~a5052 & ~a5050;
assign a5056 = l772 & l86;
assign a5058 = l774 & ~l86;
assign a5060 = ~a5058 & ~a5056;
assign a5062 = ~a5060 & a832;
assign a5064 = ~a832 & l768;
assign a5066 = ~a5064 & ~a5062;
assign a5068 = l776 & l86;
assign a5070 = l778 & ~l86;
assign a5072 = ~a5070 & ~a5068;
assign a5074 = ~a5072 & a832;
assign a5076 = ~a832 & l772;
assign a5078 = ~a5076 & ~a5074;
assign a5080 = l780 & l86;
assign a5082 = l782 & ~l86;
assign a5084 = ~a5082 & ~a5080;
assign a5086 = ~a5084 & a832;
assign a5088 = ~a832 & l776;
assign a5090 = ~a5088 & ~a5086;
assign a5092 = l784 & l86;
assign a5094 = l786 & ~l86;
assign a5096 = ~a5094 & ~a5092;
assign a5098 = ~a5096 & a832;
assign a5100 = ~a832 & l780;
assign a5102 = ~a5100 & ~a5098;
assign a5104 = a3622 & l86;
assign a5106 = l788 & ~l86;
assign a5108 = ~a5106 & ~a5104;
assign a5110 = ~a5108 & a832;
assign a5112 = ~a832 & l784;
assign a5114 = ~a5112 & ~a5110;
assign a5116 = ~a3258 & a832;
assign a5118 = ~a832 & l818;
assign a5120 = ~a5118 & ~a5116;
assign p0 = ~a826;

assert property (~p0);

endmodule
