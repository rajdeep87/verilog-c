module m139442p (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338;

output p0;

wire a858,a874,a902,a946,a962,a982,a1042,a1066,a1088,a1100,a1254,a1264,a1274,a1284,a1342,
a1358,a1386,a1430,a1446,a1466,a1526,a1550,a1572,a1584,a1738,a1748,a1758,a1768,a1826,a1842,
a1870,a1914,a1930,a1950,a2010,a2034,a2056,a2068,a2222,a2232,a2242,a2252,a2310,a2326,a2354,
a2398,a2414,a2434,a2494,a2518,a2540,a2552,a2706,a2716,a2726,a2736,a2742,a2750,a2760,a2768,
a2770,a7676,c1,a802,a804,a806,a808,a810,a812,a814,a816,a818,a820,a822,a824,
a826,a828,a830,a832,a834,a836,a838,a840,a842,a844,a846,a848,a850,a852,a854,
a856,a860,a862,a864,a866,a868,a870,a872,a876,a878,a880,a882,a884,a886,a888,
a890,a892,a894,a896,a898,a900,a904,a906,a908,a910,a912,a914,a916,a918,a920,
a922,a924,a926,a928,a930,a932,a934,a936,a938,a940,a942,a944,a948,a950,a952,
a954,a956,a958,a960,a964,a966,a968,a970,a972,a974,a976,a978,a980,a984,a986,
a988,a990,a992,a994,a996,a998,a1000,a1002,a1004,a1006,a1008,a1010,a1012,a1014,a1016,
a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,a1038,a1040,a1044,a1046,a1048,
a1050,a1052,a1054,a1056,a1058,a1060,a1062,a1064,a1068,a1070,a1072,a1074,a1076,a1078,a1080,
a1082,a1084,a1086,a1090,a1092,a1094,a1096,a1098,a1102,a1104,a1106,a1108,a1110,a1112,a1114,
a1116,a1118,a1120,a1122,a1124,a1126,a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,
a1146,a1148,a1150,a1152,a1154,a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,
a1176,a1178,a1180,a1182,a1184,a1186,a1188,a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,
a1206,a1208,a1210,a1212,a1214,a1216,a1218,a1220,a1222,a1224,a1226,a1228,a1230,a1232,a1234,
a1236,a1238,a1240,a1242,a1244,a1246,a1248,a1250,a1252,a1256,a1258,a1260,a1262,a1266,a1268,
a1270,a1272,a1276,a1278,a1280,a1282,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,
a1304,a1306,a1308,a1310,a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,
a1334,a1336,a1338,a1340,a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1360,a1362,a1364,a1366,
a1368,a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1388,a1390,a1392,a1394,a1396,a1398,
a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1426,a1428,
a1432,a1434,a1436,a1438,a1440,a1442,a1444,a1448,a1450,a1452,a1454,a1456,a1458,a1460,a1462,
a1464,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1482,a1484,a1486,a1488,a1490,a1492,a1494,
a1496,a1498,a1500,a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,a1518,a1520,a1522,a1524,
a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,a1548,a1552,a1554,a1556,a1558,
a1560,a1562,a1564,a1566,a1568,a1570,a1574,a1576,a1578,a1580,a1582,a1586,a1588,a1590,a1592,
a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,a1610,a1612,a1614,a1616,a1618,a1620,a1622,
a1624,a1626,a1628,a1630,a1632,a1634,a1636,a1638,a1640,a1642,a1644,a1646,a1648,a1650,a1652,
a1654,a1656,a1658,a1660,a1662,a1664,a1666,a1668,a1670,a1672,a1674,a1676,a1678,a1680,a1682,
a1684,a1686,a1688,a1690,a1692,a1694,a1696,a1698,a1700,a1702,a1704,a1706,a1708,a1710,a1712,
a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,a1732,a1734,a1736,a1740,a1742,a1744,
a1746,a1750,a1752,a1754,a1756,a1760,a1762,a1764,a1766,a1770,a1772,a1774,a1776,a1778,a1780,
a1782,a1784,a1786,a1788,a1790,a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,
a1812,a1814,a1816,a1818,a1820,a1822,a1824,a1828,a1830,a1832,a1834,a1836,a1838,a1840,a1844,
a1846,a1848,a1850,a1852,a1854,a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1872,a1874,a1876,
a1878,a1880,a1882,a1884,a1886,a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,
a1908,a1910,a1912,a1916,a1918,a1920,a1922,a1924,a1926,a1928,a1932,a1934,a1936,a1938,a1940,
a1942,a1944,a1946,a1948,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,a1972,
a1974,a1976,a1978,a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,a1998,a2000,a2002,
a2004,a2006,a2008,a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,a2030,a2032,a2036,
a2038,a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2058,a2060,a2062,a2064,a2066,a2070,
a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,a2090,a2092,a2094,a2096,a2098,a2100,
a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,a2120,a2122,a2124,a2126,a2128,a2130,
a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,a2152,a2154,a2156,a2158,a2160,
a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,a2178,a2180,a2182,a2184,a2186,a2188,a2190,
a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,a2208,a2210,a2212,a2214,a2216,a2218,a2220,
a2224,a2226,a2228,a2230,a2234,a2236,a2238,a2240,a2244,a2246,a2248,a2250,a2254,a2256,a2258,
a2260,a2262,a2264,a2266,a2268,a2270,a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,
a2290,a2292,a2294,a2296,a2298,a2300,a2302,a2304,a2306,a2308,a2312,a2314,a2316,a2318,a2320,
a2322,a2324,a2328,a2330,a2332,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,a2350,a2352,
a2356,a2358,a2360,a2362,a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,
a2386,a2388,a2390,a2392,a2394,a2396,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2416,a2418,
a2420,a2422,a2424,a2426,a2428,a2430,a2432,a2436,a2438,a2440,a2442,a2444,a2446,a2448,a2450,
a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,a2478,a2480,
a2482,a2484,a2486,a2488,a2490,a2492,a2496,a2498,a2500,a2502,a2504,a2506,a2508,a2510,a2512,
a2514,a2516,a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,a2542,a2544,a2546,
a2548,a2550,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,a2572,a2574,a2576,a2578,
a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,a2602,a2604,a2606,a2608,
a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,a2630,a2632,a2634,a2636,a2638,
a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,a2662,a2664,a2666,a2668,
a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,a2692,a2694,a2696,a2698,
a2700,a2702,a2704,a2708,a2710,a2712,a2714,a2718,a2720,a2722,a2724,a2728,a2730,a2732,a2734,
a2738,a2740,a2744,a2746,a2748,a2752,a2754,a2756,a2758,a2762,a2764,a2766,a2772,a2774,a2776,
a2778,a2780,a2782,a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,
a2808,a2810,a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,
a2838,a2840,a2842,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,
a2868,a2870,a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,
a2898,a2900,a2902,a2904,a2906,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,
a2928,a2930,a2932,a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,
a2958,a2960,a2962,a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,
a2988,a2990,a2992,a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,
a3018,a3020,a3022,a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,
a3048,a3050,a3052,a3054,a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,
a3078,a3080,a3082,a3084,a3086,a3088,a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,
a3108,a3110,a3112,a3114,a3116,a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,
a3138,a3140,a3142,a3144,a3146,a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,
a3168,a3170,a3172,a3174,a3176,a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,
a3198,a3200,a3202,a3204,a3206,a3208,a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,
a3228,a3230,a3232,a3234,a3236,a3238,a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,
a3258,a3260,a3262,a3264,a3266,a3268,a3270,a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,
a3288,a3290,a3292,a3294,a3296,a3298,a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,
a3318,a3320,a3322,a3324,a3326,a3328,a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,
a3348,a3350,a3352,a3354,a3356,a3358,a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,
a3378,a3380,a3382,a3384,a3386,a3388,a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,
a3408,a3410,a3412,a3414,a3416,a3418,a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,
a3438,a3440,a3442,a3444,a3446,a3448,a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,
a3468,a3470,a3472,a3474,a3476,a3478,a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,
a3498,a3500,a3502,a3504,a3506,a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,
a3528,a3530,a3532,a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,
a3558,a3560,a3562,a3564,a3566,a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,
a3588,a3590,a3592,a3594,a3596,a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,
a3618,a3620,a3622,a3624,a3626,a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,
a3648,a3650,a3652,a3654,a3656,a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,
a3678,a3680,a3682,a3684,a3686,a3688,a3690,a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,
a3708,a3710,a3712,a3714,a3716,a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,
a3738,a3740,a3742,a3744,a3746,a3748,a3750,a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,
a3768,a3770,a3772,a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,
a3798,a3800,a3802,a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,
a3828,a3830,a3832,a3834,a3836,a3838,a3840,a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,
a3858,a3860,a3862,a3864,a3866,a3868,a3870,a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,
a3888,a3890,a3892,a3894,a3896,a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,
a3918,a3920,a3922,a3924,a3926,a3928,a3930,a3932,a3934,a3936,a3938,a3940,a3942,a3944,a3946,
a3948,a3950,a3952,a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,
a3978,a3980,a3982,a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,
a4008,a4010,a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,
a4038,a4040,a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,
a4068,a4070,a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,a4096,
a4098,a4100,a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4124,a4126,
a4128,a4130,a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,a4152,a4154,a4156,
a4158,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,a4184,a4186,
a4188,a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,a4214,a4216,
a4218,a4220,a4222,a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,a4244,a4246,
a4248,a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,a4274,a4276,
a4278,a4280,a4282,a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,a4306,
a4308,a4310,a4312,a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,a4334,a4336,
a4338,a4340,a4342,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,
a4368,a4370,a4372,a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,a4394,a4396,
a4398,a4400,a4402,a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,
a4428,a4430,a4432,a4434,a4436,a4438,a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,
a4458,a4460,a4462,a4464,a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4482,a4484,a4486,
a4488,a4490,a4492,a4494,a4496,a4498,a4500,a4502,a4504,a4506,a4508,a4510,a4512,a4514,a4516,
a4518,a4520,a4522,a4524,a4526,a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,
a4548,a4550,a4552,a4554,a4556,a4558,a4560,a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,
a4578,a4580,a4582,a4584,a4586,a4588,a4590,a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,
a4608,a4610,a4612,a4614,a4616,a4618,a4620,a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,
a4638,a4640,a4642,a4644,a4646,a4648,a4650,a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,
a4668,a4670,a4672,a4674,a4676,a4678,a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,a4696,
a4698,a4700,a4702,a4704,a4706,a4708,a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,a4726,
a4728,a4730,a4732,a4734,a4736,a4738,a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,a4756,
a4758,a4760,a4762,a4764,a4766,a4768,a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4784,a4786,
a4788,a4790,a4792,a4794,a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,
a4818,a4820,a4822,a4824,a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,a4844,a4846,
a4848,a4850,a4852,a4854,a4856,a4858,a4860,a4862,a4864,a4866,a4868,a4870,a4872,a4874,a4876,
a4878,a4880,a4882,a4884,a4886,a4888,a4890,a4892,a4894,a4896,a4898,a4900,a4902,a4904,a4906,
a4908,a4910,a4912,a4914,a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,
a4938,a4940,a4942,a4944,a4946,a4948,a4950,a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,
a4968,a4970,a4972,a4974,a4976,a4978,a4980,a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,
a4998,a5000,a5002,a5004,a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,
a5028,a5030,a5032,a5034,a5036,a5038,a5040,a5042,a5044,a5046,a5048,a5050,a5052,a5054,a5056,
a5058,a5060,a5062,a5064,a5066,a5068,a5070,a5072,a5074,a5076,a5078,a5080,a5082,a5084,a5086,
a5088,a5090,a5092,a5094,a5096,a5098,a5100,a5102,a5104,a5106,a5108,a5110,a5112,a5114,a5116,
a5118,a5120,a5122,a5124,a5126,a5128,a5130,a5132,a5134,a5136,a5138,a5140,a5142,a5144,a5146,
a5148,a5150,a5152,a5154,a5156,a5158,a5160,a5162,a5164,a5166,a5168,a5170,a5172,a5174,a5176,
a5178,a5180,a5182,a5184,a5186,a5188,a5190,a5192,a5194,a5196,a5198,a5200,a5202,a5204,a5206,
a5208,a5210,a5212,a5214,a5216,a5218,a5220,a5222,a5224,a5226,a5228,a5230,a5232,a5234,a5236,
a5238,a5240,a5242,a5244,a5246,a5248,a5250,a5252,a5254,a5256,a5258,a5260,a5262,a5264,a5266,
a5268,a5270,a5272,a5274,a5276,a5278,a5280,a5282,a5284,a5286,a5288,a5290,a5292,a5294,a5296,
a5298,a5300,a5302,a5304,a5306,a5308,a5310,a5312,a5314,a5316,a5318,a5320,a5322,a5324,a5326,
a5328,a5330,a5332,a5334,a5336,a5338,a5340,a5342,a5344,a5346,a5348,a5350,a5352,a5354,a5356,
a5358,a5360,a5362,a5364,a5366,a5368,a5370,a5372,a5374,a5376,a5378,a5380,a5382,a5384,a5386,
a5388,a5390,a5392,a5394,a5396,a5398,a5400,a5402,a5404,a5406,a5408,a5410,a5412,a5414,a5416,
a5418,a5420,a5422,a5424,a5426,a5428,a5430,a5432,a5434,a5436,a5438,a5440,a5442,a5444,a5446,
a5448,a5450,a5452,a5454,a5456,a5458,a5460,a5462,a5464,a5466,a5468,a5470,a5472,a5474,a5476,
a5478,a5480,a5482,a5484,a5486,a5488,a5490,a5492,a5494,a5496,a5498,a5500,a5502,a5504,a5506,
a5508,a5510,a5512,a5514,a5516,a5518,a5520,a5522,a5524,a5526,a5528,a5530,a5532,a5534,a5536,
a5538,a5540,a5542,a5544,a5546,a5548,a5550,a5552,a5554,a5556,a5558,a5560,a5562,a5564,a5566,
a5568,a5570,a5572,a5574,a5576,a5578,a5580,a5582,a5584,a5586,a5588,a5590,a5592,a5594,a5596,
a5598,a5600,a5602,a5604,a5606,a5608,a5610,a5612,a5614,a5616,a5618,a5620,a5622,a5624,a5626,
a5628,a5630,a5632,a5634,a5636,a5638,a5640,a5642,a5644,a5646,a5648,a5650,a5652,a5654,a5656,
a5658,a5660,a5662,a5664,a5666,a5668,a5670,a5672,a5674,a5676,a5678,a5680,a5682,a5684,a5686,
a5688,a5690,a5692,a5694,a5696,a5698,a5700,a5702,a5704,a5706,a5708,a5710,a5712,a5714,a5716,
a5718,a5720,a5722,a5724,a5726,a5728,a5730,a5732,a5734,a5736,a5738,a5740,a5742,a5744,a5746,
a5748,a5750,a5752,a5754,a5756,a5758,a5760,a5762,a5764,a5766,a5768,a5770,a5772,a5774,a5776,
a5778,a5780,a5782,a5784,a5786,a5788,a5790,a5792,a5794,a5796,a5798,a5800,a5802,a5804,a5806,
a5808,a5810,a5812,a5814,a5816,a5818,a5820,a5822,a5824,a5826,a5828,a5830,a5832,a5834,a5836,
a5838,a5840,a5842,a5844,a5846,a5848,a5850,a5852,a5854,a5856,a5858,a5860,a5862,a5864,a5866,
a5868,a5870,a5872,a5874,a5876,a5878,a5880,a5882,a5884,a5886,a5888,a5890,a5892,a5894,a5896,
a5898,a5900,a5902,a5904,a5906,a5908,a5910,a5912,a5914,a5916,a5918,a5920,a5922,a5924,a5926,
a5928,a5930,a5932,a5934,a5936,a5938,a5940,a5942,a5944,a5946,a5948,a5950,a5952,a5954,a5956,
a5958,a5960,a5962,a5964,a5966,a5968,a5970,a5972,a5974,a5976,a5978,a5980,a5982,a5984,a5986,
a5988,a5990,a5992,a5994,a5996,a5998,a6000,a6002,a6004,a6006,a6008,a6010,a6012,a6014,a6016,
a6018,a6020,a6022,a6024,a6026,a6028,a6030,a6032,a6034,a6036,a6038,a6040,a6042,a6044,a6046,
a6048,a6050,a6052,a6054,a6056,a6058,a6060,a6062,a6064,a6066,a6068,a6070,a6072,a6074,a6076,
a6078,a6080,a6082,a6084,a6086,a6088,a6090,a6092,a6094,a6096,a6098,a6100,a6102,a6104,a6106,
a6108,a6110,a6112,a6114,a6116,a6118,a6120,a6122,a6124,a6126,a6128,a6130,a6132,a6134,a6136,
a6138,a6140,a6142,a6144,a6146,a6148,a6150,a6152,a6154,a6156,a6158,a6160,a6162,a6164,a6166,
a6168,a6170,a6172,a6174,a6176,a6178,a6180,a6182,a6184,a6186,a6188,a6190,a6192,a6194,a6196,
a6198,a6200,a6202,a6204,a6206,a6208,a6210,a6212,a6214,a6216,a6218,a6220,a6222,a6224,a6226,
a6228,a6230,a6232,a6234,a6236,a6238,a6240,a6242,a6244,a6246,a6248,a6250,a6252,a6254,a6256,
a6258,a6260,a6262,a6264,a6266,a6268,a6270,a6272,a6274,a6276,a6278,a6280,a6282,a6284,a6286,
a6288,a6290,a6292,a6294,a6296,a6298,a6300,a6302,a6304,a6306,a6308,a6310,a6312,a6314,a6316,
a6318,a6320,a6322,a6324,a6326,a6328,a6330,a6332,a6334,a6336,a6338,a6340,a6342,a6344,a6346,
a6348,a6350,a6352,a6354,a6356,a6358,a6360,a6362,a6364,a6366,a6368,a6370,a6372,a6374,a6376,
a6378,a6380,a6382,a6384,a6386,a6388,a6390,a6392,a6394,a6396,a6398,a6400,a6402,a6404,a6406,
a6408,a6410,a6412,a6414,a6416,a6418,a6420,a6422,a6424,a6426,a6428,a6430,a6432,a6434,a6436,
a6438,a6440,a6442,a6444,a6446,a6448,a6450,a6452,a6454,a6456,a6458,a6460,a6462,a6464,a6466,
a6468,a6470,a6472,a6474,a6476,a6478,a6480,a6482,a6484,a6486,a6488,a6490,a6492,a6494,a6496,
a6498,a6500,a6502,a6504,a6506,a6508,a6510,a6512,a6514,a6516,a6518,a6520,a6522,a6524,a6526,
a6528,a6530,a6532,a6534,a6536,a6538,a6540,a6542,a6544,a6546,a6548,a6550,a6552,a6554,a6556,
a6558,a6560,a6562,a6564,a6566,a6568,a6570,a6572,a6574,a6576,a6578,a6580,a6582,a6584,a6586,
a6588,a6590,a6592,a6594,a6596,a6598,a6600,a6602,a6604,a6606,a6608,a6610,a6612,a6614,a6616,
a6618,a6620,a6622,a6624,a6626,a6628,a6630,a6632,a6634,a6636,a6638,a6640,a6642,a6644,a6646,
a6648,a6650,a6652,a6654,a6656,a6658,a6660,a6662,a6664,a6666,a6668,a6670,a6672,a6674,a6676,
a6678,a6680,a6682,a6684,a6686,a6688,a6690,a6692,a6694,a6696,a6698,a6700,a6702,a6704,a6706,
a6708,a6710,a6712,a6714,a6716,a6718,a6720,a6722,a6724,a6726,a6728,a6730,a6732,a6734,a6736,
a6738,a6740,a6742,a6744,a6746,a6748,a6750,a6752,a6754,a6756,a6758,a6760,a6762,a6764,a6766,
a6768,a6770,a6772,a6774,a6776,a6778,a6780,a6782,a6784,a6786,a6788,a6790,a6792,a6794,a6796,
a6798,a6800,a6802,a6804,a6806,a6808,a6810,a6812,a6814,a6816,a6818,a6820,a6822,a6824,a6826,
a6828,a6830,a6832,a6834,a6836,a6838,a6840,a6842,a6844,a6846,a6848,a6850,a6852,a6854,a6856,
a6858,a6860,a6862,a6864,a6866,a6868,a6870,a6872,a6874,a6876,a6878,a6880,a6882,a6884,a6886,
a6888,a6890,a6892,a6894,a6896,a6898,a6900,a6902,a6904,a6906,a6908,a6910,a6912,a6914,a6916,
a6918,a6920,a6922,a6924,a6926,a6928,a6930,a6932,a6934,a6936,a6938,a6940,a6942,a6944,a6946,
a6948,a6950,a6952,a6954,a6956,a6958,a6960,a6962,a6964,a6966,a6968,a6970,a6972,a6974,a6976,
a6978,a6980,a6982,a6984,a6986,a6988,a6990,a6992,a6994,a6996,a6998,a7000,a7002,a7004,a7006,
a7008,a7010,a7012,a7014,a7016,a7018,a7020,a7022,a7024,a7026,a7028,a7030,a7032,a7034,a7036,
a7038,a7040,a7042,a7044,a7046,a7048,a7050,a7052,a7054,a7056,a7058,a7060,a7062,a7064,a7066,
a7068,a7070,a7072,a7074,a7076,a7078,a7080,a7082,a7084,a7086,a7088,a7090,a7092,a7094,a7096,
a7098,a7100,a7102,a7104,a7106,a7108,a7110,a7112,a7114,a7116,a7118,a7120,a7122,a7124,a7126,
a7128,a7130,a7132,a7134,a7136,a7138,a7140,a7142,a7144,a7146,a7148,a7150,a7152,a7154,a7156,
a7158,a7160,a7162,a7164,a7166,a7168,a7170,a7172,a7174,a7176,a7178,a7180,a7182,a7184,a7186,
a7188,a7190,a7192,a7194,a7196,a7198,a7200,a7202,a7204,a7206,a7208,a7210,a7212,a7214,a7216,
a7218,a7220,a7222,a7224,a7226,a7228,a7230,a7232,a7234,a7236,a7238,a7240,a7242,a7244,a7246,
a7248,a7250,a7252,a7254,a7256,a7258,a7260,a7262,a7264,a7266,a7268,a7270,a7272,a7274,a7276,
a7278,a7280,a7282,a7284,a7286,a7288,a7290,a7292,a7294,a7296,a7298,a7300,a7302,a7304,a7306,
a7308,a7310,a7312,a7314,a7316,a7318,a7320,a7322,a7324,a7326,a7328,a7330,a7332,a7334,a7336,
a7338,a7340,a7342,a7344,a7346,a7348,a7350,a7352,a7354,a7356,a7358,a7360,a7362,a7364,a7366,
a7368,a7370,a7372,a7374,a7376,a7378,a7380,a7382,a7384,a7386,a7388,a7390,a7392,a7394,a7396,
a7398,a7400,a7402,a7404,a7406,a7408,a7410,a7412,a7414,a7416,a7418,a7420,a7422,a7424,a7426,
a7428,a7430,a7432,a7434,a7436,a7438,a7440,a7442,a7444,a7446,a7448,a7450,a7452,a7454,a7456,
a7458,a7460,a7462,a7464,a7466,a7468,a7470,a7472,a7474,a7476,a7478,a7480,a7482,a7484,a7486,
a7488,a7490,a7492,a7494,a7496,a7498,a7500,a7502,a7504,a7506,a7508,a7510,a7512,a7514,a7516,
a7518,a7520,a7522,a7524,a7526,a7528,a7530,a7532,a7534,a7536,a7538,a7540,a7542,a7544,a7546,
a7548,a7550,a7552,a7554,a7556,a7558,a7560,a7562,a7564,a7566,a7568,a7570,a7572,a7574,a7576,
a7578,a7580,a7582,a7584,a7586,a7588,a7590,a7592,a7594,a7596,a7598,a7600,a7602,a7604,a7606,
a7608,a7610,a7612,a7614,a7616,a7618,a7620,a7622,a7624,a7626,a7628,a7630,a7632,a7634,a7636,
a7638,a7640,a7642,a7644,a7646,a7648,a7650,a7652,a7654,a7656,a7658,a7660,a7662,a7664,a7666,
a7668,a7670,a7672,a7674,a7678,p0;

reg l340,l342,l344,l346,l348,l350,l352,l354,l356,l358,l360,l362,l364,l366,l368,
l370,l372,l374,l376,l378,l380,l382,l384,l386,l388,l390,l392,l394,l396,l398,
l400,l402,l404,l406,l408,l410,l412,l414,l416,l418,l420,l422,l424,l426,l428,
l430,l432,l434,l436,l438,l440,l442,l444,l446,l448,l450,l452,l454,l456,l458,
l460,l462,l464,l466,l468,l470,l472,l474,l476,l478,l480,l482,l484,l486,l488,
l490,l492,l494,l496,l498,l500,l502,l504,l506,l508,l510,l512,l514,l516,l518,
l520,l522,l524,l526,l528,l530,l532,l534,l536,l538,l540,l542,l544,l546,l548,
l550,l552,l554,l556,l558,l560,l562,l564,l566,l568,l570,l572,l574,l576,l578,
l580,l582,l584,l586,l588,l590,l592,l594,l596,l598,l600,l602,l604,l606,l608,
l610,l612,l614,l616,l618,l620,l622,l624,l626,l628,l630,l632,l634,l636,l638,
l640,l642,l644,l646,l648,l650,l652,l654,l656,l658,l660,l662,l664,l666,l668,
l670,l672,l674,l676,l678,l680,l682,l684,l686,l688,l690,l692,l694,l696,l698,
l700,l702,l704,l706,l708,l710,l712,l714,l716,l718,l720,l722,l724,l726,l728,
l730,l732,l734,l736,l738,l740,l742,l744,l746,l748,l750,l752,l754,l756,l758,
l760,l762,l764,l766,l768,l770,l772,l774,l776,l778,l780,l782,l784,l786,l788,
l790,l792,l794,l796,l798,l800;

initial
begin
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
   l392 = 0;
   l394 = 0;
   l396 = 0;
   l398 = 0;
   l400 = 0;
   l402 = 0;
   l404 = 0;
   l406 = 0;
   l408 = 0;
   l410 = 0;
   l412 = 0;
   l414 = 0;
   l416 = 0;
   l418 = 0;
   l420 = 0;
   l422 = 0;
   l424 = 0;
   l426 = 0;
   l428 = 0;
   l430 = 0;
   l432 = 0;
   l434 = 0;
   l436 = 0;
   l438 = 0;
   l440 = 0;
   l442 = 0;
   l444 = 0;
   l446 = 0;
   l448 = 0;
   l450 = 0;
   l452 = 0;
   l454 = 0;
   l456 = 0;
   l458 = 0;
   l460 = 0;
   l462 = 0;
   l464 = 0;
   l466 = 0;
   l468 = 0;
   l470 = 0;
   l472 = 0;
   l474 = 0;
   l476 = 0;
   l478 = 0;
   l480 = 0;
   l482 = 0;
   l484 = 0;
   l486 = 0;
   l488 = 0;
   l490 = 0;
   l492 = 0;
   l494 = 0;
   l496 = 0;
   l498 = 0;
   l500 = 0;
   l502 = 0;
   l504 = 0;
   l506 = 0;
   l508 = 0;
   l510 = 0;
   l512 = 0;
   l514 = 0;
   l516 = 0;
   l518 = 0;
   l520 = 0;
   l522 = 0;
   l524 = 0;
   l526 = 0;
   l528 = 0;
   l530 = 0;
   l532 = 0;
   l534 = 0;
   l536 = 0;
   l538 = 0;
   l540 = 0;
   l542 = 0;
   l544 = 0;
   l546 = 0;
   l548 = 0;
   l550 = 0;
   l552 = 0;
   l554 = 0;
   l556 = 0;
   l558 = 0;
   l560 = 0;
   l562 = 0;
   l564 = 0;
   l566 = 0;
   l568 = 0;
   l570 = 0;
   l572 = 0;
   l574 = 0;
   l576 = 0;
   l578 = 0;
   l580 = 0;
   l582 = 0;
   l584 = 0;
   l586 = 0;
   l588 = 0;
   l590 = 0;
   l592 = 0;
   l594 = 0;
   l596 = 0;
   l598 = 0;
   l600 = 0;
   l602 = 0;
   l604 = 0;
   l606 = 0;
   l608 = 0;
   l610 = 0;
   l612 = 0;
   l614 = 0;
   l616 = 0;
   l618 = 0;
   l620 = 0;
   l622 = 0;
   l624 = 0;
   l626 = 0;
   l628 = 0;
   l630 = 0;
   l632 = 0;
   l634 = 0;
   l636 = 0;
   l638 = 0;
   l640 = 0;
   l642 = 0;
   l644 = 0;
   l646 = 0;
   l648 = 0;
   l650 = 0;
   l652 = 0;
   l654 = 0;
   l656 = 0;
   l658 = 0;
   l660 = 0;
   l662 = 0;
   l664 = 0;
   l666 = 0;
   l668 = 0;
   l670 = 0;
   l672 = 0;
   l674 = 0;
   l676 = 0;
   l678 = 0;
   l680 = 0;
   l682 = 0;
   l684 = 0;
   l686 = 0;
   l688 = 0;
   l690 = 0;
   l692 = 0;
   l694 = 0;
   l696 = 0;
   l698 = 0;
   l700 = 0;
   l702 = 0;
   l704 = 0;
   l706 = 0;
   l708 = 0;
   l710 = 0;
   l712 = 0;
   l714 = 0;
   l716 = 0;
   l718 = 0;
   l720 = 0;
   l722 = 0;
   l724 = 0;
   l726 = 0;
   l728 = 0;
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
end

always @(posedge i2)
   l340 <= i2;

always @(posedge i4)
   l342 <= i4;

always @(posedge i6)
   l344 <= i6;

always @(posedge i8)
   l346 <= i8;

always @(posedge i10)
   l348 <= i10;

always @(posedge i12)
   l350 <= i12;

always @(posedge i14)
   l352 <= i14;

always @(posedge i16)
   l354 <= i16;

always @(posedge i18)
   l356 <= i18;

always @(posedge i20)
   l358 <= i20;

always @(posedge i22)
   l360 <= i22;

always @(posedge i24)
   l362 <= i24;

always @(posedge i26)
   l364 <= i26;

always @(posedge i28)
   l366 <= i28;

always @(posedge i30)
   l368 <= i30;

always @(posedge i32)
   l370 <= i32;

always @(posedge i34)
   l372 <= i34;

always @(posedge i36)
   l374 <= i36;

always @(posedge i38)
   l376 <= i38;

always @(posedge i40)
   l378 <= i40;

always @(posedge i42)
   l380 <= i42;

always @(posedge i44)
   l382 <= i44;

always @(posedge i46)
   l384 <= i46;

always @(posedge i48)
   l386 <= i48;

always @(posedge i50)
   l388 <= i50;

always @(posedge i52)
   l390 <= i52;

always @(posedge i54)
   l392 <= i54;

always @(posedge i56)
   l394 <= i56;

always @(posedge i58)
   l396 <= i58;

always @(posedge i60)
   l398 <= i60;

always @(posedge i62)
   l400 <= i62;

always @(posedge i64)
   l402 <= i64;

always @(posedge i66)
   l404 <= i66;

always @(posedge i68)
   l406 <= i68;

always @(posedge a858)
   l408 <= a858;

always @(posedge a874)
   l410 <= a874;

always @(posedge i70)
   l412 <= i70;

always @(posedge i72)
   l414 <= i72;

always @(posedge a902)
   l416 <= a902;

always @(posedge i74)
   l418 <= i74;

always @(posedge i76)
   l420 <= i76;

always @(posedge a946)
   l422 <= a946;

always @(posedge a962)
   l424 <= a962;

always @(posedge i78)
   l426 <= i78;

always @(posedge i80)
   l428 <= i80;

always @(posedge a982)
   l430 <= a982;

always @(posedge a1042)
   l432 <= a1042;

always @(posedge a1066)
   l434 <= a1066;

always @(posedge a1088)
   l436 <= a1088;

always @(posedge i82)
   l438 <= i82;

always @(posedge i84)
   l440 <= i84;

always @(posedge i86)
   l442 <= i86;

always @(posedge i88)
   l444 <= i88;

always @(posedge a1100)
   l446 <= a1100;

always @(posedge a1254)
   l448 <= a1254;

always @(posedge a1264)
   l450 <= a1264;

always @(posedge a1274)
   l452 <= a1274;

always @(posedge a1284)
   l454 <= a1284;

always @(posedge i90)
   l456 <= i90;

always @(posedge i92)
   l458 <= i92;

always @(posedge a1342)
   l460 <= a1342;

always @(posedge a1358)
   l462 <= a1358;

always @(posedge i94)
   l464 <= i94;

always @(posedge i96)
   l466 <= i96;

always @(posedge a1386)
   l468 <= a1386;

always @(posedge i98)
   l470 <= i98;

always @(posedge i100)
   l472 <= i100;

always @(posedge a1430)
   l474 <= a1430;

always @(posedge a1446)
   l476 <= a1446;

always @(posedge i102)
   l478 <= i102;

always @(posedge i104)
   l480 <= i104;

always @(posedge a1466)
   l482 <= a1466;

always @(posedge a1526)
   l484 <= a1526;

always @(posedge a1550)
   l486 <= a1550;

always @(posedge a1572)
   l488 <= a1572;

always @(posedge i106)
   l490 <= i106;

always @(posedge i108)
   l492 <= i108;

always @(posedge i110)
   l494 <= i110;

always @(posedge i112)
   l496 <= i112;

always @(posedge a1584)
   l498 <= a1584;

always @(posedge a1738)
   l500 <= a1738;

always @(posedge a1748)
   l502 <= a1748;

always @(posedge a1758)
   l504 <= a1758;

always @(posedge a1768)
   l506 <= a1768;

always @(posedge i114)
   l508 <= i114;

always @(posedge i116)
   l510 <= i116;

always @(posedge a1826)
   l512 <= a1826;

always @(posedge a1842)
   l514 <= a1842;

always @(posedge i118)
   l516 <= i118;

always @(posedge i120)
   l518 <= i120;

always @(posedge a1870)
   l520 <= a1870;

always @(posedge i122)
   l522 <= i122;

always @(posedge i124)
   l524 <= i124;

always @(posedge a1914)
   l526 <= a1914;

always @(posedge a1930)
   l528 <= a1930;

always @(posedge i126)
   l530 <= i126;

always @(posedge i128)
   l532 <= i128;

always @(posedge a1950)
   l534 <= a1950;

always @(posedge a2010)
   l536 <= a2010;

always @(posedge a2034)
   l538 <= a2034;

always @(posedge a2056)
   l540 <= a2056;

always @(posedge i130)
   l542 <= i130;

always @(posedge i132)
   l544 <= i132;

always @(posedge i134)
   l546 <= i134;

always @(posedge i136)
   l548 <= i136;

always @(posedge a2068)
   l550 <= a2068;

always @(posedge a2222)
   l552 <= a2222;

always @(posedge a2232)
   l554 <= a2232;

always @(posedge a2242)
   l556 <= a2242;

always @(posedge a2252)
   l558 <= a2252;

always @(posedge i138)
   l560 <= i138;

always @(posedge i140)
   l562 <= i140;

always @(posedge a2310)
   l564 <= a2310;

always @(posedge a2326)
   l566 <= a2326;

always @(posedge i142)
   l568 <= i142;

always @(posedge i144)
   l570 <= i144;

always @(posedge a2354)
   l572 <= a2354;

always @(posedge i146)
   l574 <= i146;

always @(posedge i148)
   l576 <= i148;

always @(posedge a2398)
   l578 <= a2398;

always @(posedge a2414)
   l580 <= a2414;

always @(posedge i150)
   l582 <= i150;

always @(posedge i152)
   l584 <= i152;

always @(posedge a2434)
   l586 <= a2434;

always @(posedge a2494)
   l588 <= a2494;

always @(posedge a2518)
   l590 <= a2518;

always @(posedge a2540)
   l592 <= a2540;

always @(posedge i154)
   l594 <= i154;

always @(posedge i156)
   l596 <= i156;

always @(posedge i158)
   l598 <= i158;

always @(posedge i160)
   l600 <= i160;

always @(posedge a2552)
   l602 <= a2552;

always @(posedge a2706)
   l604 <= a2706;

always @(posedge a2716)
   l606 <= a2716;

always @(posedge a2726)
   l608 <= a2726;

always @(posedge a2736)
   l610 <= a2736;

always @(posedge i162)
   l612 <= i162;

always @(posedge a2742)
   l614 <= a2742;

always @(posedge i164)
   l616 <= i164;

always @(posedge i166)
   l618 <= i166;

always @(posedge i168)
   l620 <= i168;

always @(posedge i170)
   l622 <= i170;

always @(posedge i172)
   l624 <= i172;

always @(posedge i174)
   l626 <= i174;

always @(posedge i176)
   l628 <= i176;

always @(posedge i178)
   l630 <= i178;

always @(posedge i180)
   l632 <= i180;

always @(posedge i182)
   l634 <= i182;

always @(posedge i184)
   l636 <= i184;

always @(posedge i186)
   l638 <= i186;

always @(posedge i188)
   l640 <= i188;

always @(posedge i190)
   l642 <= i190;

always @(posedge i192)
   l644 <= i192;

always @(posedge i194)
   l646 <= i194;

always @(posedge i196)
   l648 <= i196;

always @(posedge i198)
   l650 <= i198;

always @(posedge i200)
   l652 <= i200;

always @(posedge i202)
   l654 <= i202;

always @(posedge i204)
   l656 <= i204;

always @(posedge i206)
   l658 <= i206;

always @(posedge i208)
   l660 <= i208;

always @(posedge i210)
   l662 <= i210;

always @(posedge i212)
   l664 <= i212;

always @(posedge i214)
   l666 <= i214;

always @(posedge i216)
   l668 <= i216;

always @(posedge i218)
   l670 <= i218;

always @(posedge i220)
   l672 <= i220;

always @(posedge i222)
   l674 <= i222;

always @(posedge i224)
   l676 <= i224;

always @(posedge i226)
   l678 <= i226;

always @(posedge i228)
   l680 <= i228;

always @(posedge i230)
   l682 <= i230;

always @(posedge i232)
   l684 <= i232;

always @(posedge i234)
   l686 <= i234;

always @(posedge i236)
   l688 <= i236;

always @(posedge i238)
   l690 <= i238;

always @(posedge i240)
   l692 <= i240;

always @(posedge i242)
   l694 <= i242;

always @(posedge i244)
   l696 <= i244;

always @(posedge i246)
   l698 <= i246;

always @(posedge i248)
   l700 <= i248;

always @(posedge i250)
   l702 <= i250;

always @(posedge i252)
   l704 <= i252;

always @(posedge i254)
   l706 <= i254;

always @(posedge i256)
   l708 <= i256;

always @(posedge i258)
   l710 <= i258;

always @(posedge i260)
   l712 <= i260;

always @(posedge i262)
   l714 <= i262;

always @(posedge i264)
   l716 <= i264;

always @(posedge i266)
   l718 <= i266;

always @(posedge i268)
   l720 <= i268;

always @(posedge i270)
   l722 <= i270;

always @(posedge i272)
   l724 <= i272;

always @(posedge i274)
   l726 <= i274;

always @(posedge i276)
   l728 <= i276;

always @(posedge i278)
   l730 <= i278;

always @(posedge i280)
   l732 <= i280;

always @(posedge i282)
   l734 <= i282;

always @(posedge i284)
   l736 <= i284;

always @(posedge i286)
   l738 <= i286;

always @(posedge i288)
   l740 <= i288;

always @(posedge i290)
   l742 <= i290;

always @(posedge i292)
   l744 <= i292;

always @(posedge i294)
   l746 <= i294;

always @(posedge i296)
   l748 <= i296;

always @(posedge i298)
   l750 <= i298;

always @(posedge i300)
   l752 <= i300;

always @(posedge i302)
   l754 <= i302;

always @(posedge i304)
   l756 <= i304;

always @(posedge i306)
   l758 <= i306;

always @(posedge i308)
   l760 <= i308;

always @(posedge i310)
   l762 <= i310;

always @(posedge i312)
   l764 <= i312;

always @(posedge i314)
   l766 <= i314;

always @(posedge i316)
   l768 <= i316;

always @(posedge i318)
   l770 <= i318;

always @(posedge i320)
   l772 <= i320;

always @(posedge i322)
   l774 <= i322;

always @(posedge i324)
   l776 <= i324;

always @(posedge i326)
   l778 <= i326;

always @(posedge a2750)
   l780 <= a2750;

always @(posedge a2760)
   l782 <= a2760;

always @(posedge a2768)
   l784 <= a2768;

always @(posedge i328)
   l786 <= i328;

always @(posedge a2770)
   l788 <= a2770;

always @(posedge i332)
   l790 <= i332;

always @(posedge i334)
   l792 <= i334;

always @(posedge i336)
   l794 <= i336;

always @(posedge i338)
   l796 <= i338;

always @(posedge a7676)
   l798 <= a7676;

always @(posedge c1)
   l800 <= c1;


assign a858 = a856 & l800;
assign a874 = ~a872 & l800;
assign a902 = ~a900 & l800;
assign a946 = a944 & l800;
assign a962 = ~a960 & l800;
assign a982 = ~a980 & l800;
assign a1042 = a1040 & l800;
assign a1066 = ~a1064 & l800;
assign a1088 = ~a1086 & l800;
assign a1100 = ~a1098 & l800;
assign a1254 = a1252 & l800;
assign a1264 = a1262 & l800;
assign a1274 = a1272 & l800;
assign a1284 = a1282 & l800;
assign a1342 = a1340 & l800;
assign a1358 = ~a1356 & l800;
assign a1386 = ~a1384 & l800;
assign a1430 = a1428 & l800;
assign a1446 = ~a1444 & l800;
assign a1466 = ~a1464 & l800;
assign a1526 = a1524 & l800;
assign a1550 = ~a1548 & l800;
assign a1572 = ~a1570 & l800;
assign a1584 = ~a1582 & l800;
assign a1738 = a1736 & l800;
assign a1748 = a1746 & l800;
assign a1758 = a1756 & l800;
assign a1768 = a1766 & l800;
assign a1826 = a1824 & l800;
assign a1842 = ~a1840 & l800;
assign a1870 = ~a1868 & l800;
assign a1914 = a1912 & l800;
assign a1930 = ~a1928 & l800;
assign a1950 = ~a1948 & l800;
assign a2010 = a2008 & l800;
assign a2034 = ~a2032 & l800;
assign a2056 = ~a2054 & l800;
assign a2068 = ~a2066 & l800;
assign a2222 = a2220 & l800;
assign a2232 = a2230 & l800;
assign a2242 = a2240 & l800;
assign a2252 = a2250 & l800;
assign a2310 = a2308 & l800;
assign a2326 = ~a2324 & l800;
assign a2354 = ~a2352 & l800;
assign a2398 = a2396 & l800;
assign a2414 = ~a2412 & l800;
assign a2434 = ~a2432 & l800;
assign a2494 = a2492 & l800;
assign a2518 = ~a2516 & l800;
assign a2540 = ~a2538 & l800;
assign a2552 = ~a2550 & l800;
assign a2706 = a2704 & l800;
assign a2716 = a2714 & l800;
assign a2726 = a2724 & l800;
assign a2736 = a2734 & l800;
assign a2742 = ~a2740 & l800;
assign a2750 = ~a2748 & l800;
assign a2760 = ~a2758 & l800;
assign a2768 = ~a2766 & l800;
assign a2770 = ~a2744 & l800;
assign a7676 = a7674 & l800;
assign c1 = 1;
assign a802 = l416 & ~l414;
assign a804 = l436 & l434;
assign a806 = a804 & ~l432;
assign a808 = a806 & a802;
assign a810 = ~l416 & l414;
assign a812 = a810 & a806;
assign a814 = l436 & ~l434;
assign a816 = a814 & l432;
assign a818 = a816 & a810;
assign a820 = l406 & ~l404;
assign a822 = a804 & l432;
assign a824 = a822 & a810;
assign a826 = a824 & a820;
assign a828 = ~l406 & ~l404;
assign a830 = l416 & l414;
assign a832 = a814 & ~l432;
assign a834 = a832 & a830;
assign a836 = a834 & a828;
assign a838 = a832 & a802;
assign a840 = a838 & a820;
assign a842 = a832 & l438;
assign a844 = ~a842 & l408;
assign a846 = a844 & ~a840;
assign a848 = a846 & ~a836;
assign a850 = ~a848 & ~a826;
assign a852 = ~a850 & ~a818;
assign a854 = ~a852 & ~a812;
assign a856 = ~a854 & ~a808;
assign a860 = ~a842 & l410;
assign a862 = a860 & ~a840;
assign a864 = a862 & ~a836;
assign a866 = ~a864 & ~a826;
assign a868 = ~a866 & ~a818;
assign a870 = ~a868 & ~a812;
assign a872 = a870 & ~a808;
assign a876 = ~l406 & l404;
assign a878 = ~l436 & ~l434;
assign a880 = a878 & ~l432;
assign a882 = a880 & a810;
assign a884 = a882 & a876;
assign a886 = ~l436 & l434;
assign a888 = a886 & ~l432;
assign a890 = a888 & a810;
assign a892 = a890 & a828;
assign a894 = a876 & a824;
assign a896 = ~a894 & ~l416;
assign a898 = a896 & ~a892;
assign a900 = a898 & ~a884;
assign a904 = l430 & ~l428;
assign a906 = a904 & a806;
assign a908 = ~l430 & l428;
assign a910 = a908 & a806;
assign a912 = a908 & a816;
assign a914 = l420 & ~l418;
assign a916 = a908 & a822;
assign a918 = a916 & a914;
assign a920 = ~l420 & ~l418;
assign a922 = l430 & l428;
assign a924 = a922 & a832;
assign a926 = a924 & a920;
assign a928 = a904 & a832;
assign a930 = a928 & a914;
assign a932 = ~a842 & l422;
assign a934 = a932 & ~a930;
assign a936 = a934 & ~a926;
assign a938 = ~a936 & ~a918;
assign a940 = ~a938 & ~a912;
assign a942 = ~a940 & ~a910;
assign a944 = ~a942 & ~a906;
assign a948 = ~a842 & l424;
assign a950 = a948 & ~a930;
assign a952 = a950 & ~a926;
assign a954 = ~a952 & ~a918;
assign a956 = ~a954 & ~a912;
assign a958 = ~a956 & ~a910;
assign a960 = a958 & ~a906;
assign a964 = ~l420 & l418;
assign a966 = a908 & a880;
assign a968 = a966 & a964;
assign a970 = a908 & a888;
assign a972 = a970 & a920;
assign a974 = a964 & a916;
assign a976 = ~a974 & ~l430;
assign a978 = a976 & ~a972;
assign a980 = a978 & ~a968;
assign a984 = ~l448 & l442;
assign a986 = a908 & a810;
assign a988 = ~a986 & a880;
assign a990 = a988 & ~a984;
assign a992 = ~a820 & a802;
assign a994 = ~a992 & a806;
assign a996 = ~a914 & a904;
assign a998 = ~a996 & a994;
assign a1000 = ~a828 & a810;
assign a1002 = ~a1000 & a888;
assign a1004 = ~a920 & a908;
assign a1006 = ~a1004 & a1002;
assign a1008 = ~a964 & a908;
assign a1010 = ~a876 & a810;
assign a1012 = ~a1010 & a888;
assign a1014 = a1012 & ~a1008;
assign a1016 = ~a820 & a810;
assign a1018 = ~a914 & a908;
assign a1020 = ~a1018 & ~a1016;
assign a1022 = ~a1010 & ~a1008;
assign a1024 = ~a1022 & ~a1020;
assign a1026 = ~a1024 & ~a814;
assign a1028 = a1026 & a822;
assign a1030 = a1028 & ~a878;
assign a1032 = ~a1030 & l432;
assign a1034 = ~a1032 & ~a1014;
assign a1036 = ~a1034 & ~a1006;
assign a1038 = a1036 & ~a998;
assign a1040 = a1038 & ~a990;
assign a1044 = a816 & ~l444;
assign a1046 = a878 & l432;
assign a1048 = l436 & l432;
assign a1050 = a1048 & l444;
assign a1052 = ~a1050 & a1046;
assign a1054 = ~a1052 & ~l434;
assign a1056 = a1054 & ~a1044;
assign a1058 = ~a1056 & ~a1014;
assign a1060 = a1058 & ~a1006;
assign a1062 = ~a1060 & ~a998;
assign a1064 = a1062 & ~a990;
assign a1068 = a816 & l444;
assign a1070 = a1020 & a822;
assign a1072 = ~a1070 & l436;
assign a1074 = ~a1072 & ~a1046;
assign a1076 = ~a1074 & ~a1068;
assign a1078 = ~a1076 & ~a1044;
assign a1080 = a1078 & ~a1014;
assign a1082 = a1080 & ~a1006;
assign a1084 = ~a1082 & ~a998;
assign a1086 = ~a1084 & ~a990;
assign a1090 = ~l454 & ~l452;
assign a1092 = ~a1090 & l450;
assign a1094 = a1092 & l448;
assign a1096 = a1094 & a880;
assign a1098 = ~a1096 & ~l446;
assign a1102 = ~l452 & ~l450;
assign a1104 = a1102 & ~l448;
assign a1106 = l454 & ~l452;
assign a1108 = a1106 & ~l450;
assign a1110 = a1108 & ~l448;
assign a1112 = l452 & ~l450;
assign a1114 = a1112 & ~l448;
assign a1116 = l454 & l452;
assign a1118 = a1116 & ~l450;
assign a1120 = a1118 & ~l448;
assign a1122 = ~l452 & l450;
assign a1124 = a1122 & ~l448;
assign a1126 = a1106 & l450;
assign a1128 = a1126 & ~l448;
assign a1130 = l452 & l450;
assign a1132 = a1130 & ~l448;
assign a1134 = a1108 & l448;
assign a1136 = a1118 & l448;
assign a1138 = ~a1136 & a1122;
assign a1140 = ~a1138 & ~a1112;
assign a1142 = ~a1140 & ~a1134;
assign a1144 = ~a1142 & ~a1102;
assign a1146 = ~a1144 & l448;
assign a1148 = ~a1146 & ~a1132;
assign a1150 = ~a1148 & ~a1128;
assign a1152 = ~a1150 & ~a1124;
assign a1154 = ~a1152 & ~a1120;
assign a1156 = ~a1154 & ~a1114;
assign a1158 = ~a1156 & ~a1110;
assign a1160 = ~a1158 & ~a1104;
assign a1162 = ~a1160 & ~l454;
assign a1164 = a1090 & ~l450;
assign a1166 = a1164 & ~l448;
assign a1168 = l454 & ~l450;
assign a1170 = a1168 & ~l448;
assign a1172 = a1090 & l450;
assign a1174 = a1172 & ~l448;
assign a1176 = l454 & l450;
assign a1178 = a1176 & ~l448;
assign a1180 = a1164 & l448;
assign a1182 = ~l450 & l448;
assign a1184 = a1182 & ~a1106;
assign a1186 = a1184 & ~a1180;
assign a1188 = ~a1186 & ~a1178;
assign a1190 = ~l454 & l450;
assign a1192 = a1190 & ~l448;
assign a1194 = ~a1192 & a1188;
assign a1196 = ~a1194 & ~a1128;
assign a1198 = a1196 & ~a1174;
assign a1200 = ~a1198 & ~a1170;
assign a1202 = ~l454 & ~l450;
assign a1204 = a1202 & ~l448;
assign a1206 = ~a1204 & a1200;
assign a1208 = ~a1206 & l452;
assign a1210 = a1208 & ~a1110;
assign a1212 = a1210 & ~a1166;
assign a1214 = a1212 & a1162;
assign a1216 = ~l454 & l452;
assign a1218 = ~a1116 & ~l448;
assign a1220 = a1218 & ~a1216;
assign a1222 = a1106 & ~l448;
assign a1224 = ~a1222 & a1220;
assign a1226 = a1090 & ~l448;
assign a1228 = ~a1226 & a1224;
assign a1230 = ~a1228 & ~l450;
assign a1232 = ~a1230 & a1214;
assign a1234 = ~a1116 & ~l450;
assign a1236 = a1234 & ~a1216;
assign a1238 = a1236 & ~a1108;
assign a1240 = a1238 & ~a1164;
assign a1242 = ~a1240 & ~l448;
assign a1244 = ~a1242 & a1232;
assign a1246 = ~a1244 & l448;
assign a1248 = ~a1246 & a880;
assign a1250 = ~a880 & ~l448;
assign a1252 = ~a1250 & ~a1248;
assign a1256 = ~a1244 & l450;
assign a1258 = ~a1256 & a880;
assign a1260 = ~a880 & ~l450;
assign a1262 = ~a1260 & ~a1258;
assign a1266 = ~a1244 & l452;
assign a1268 = ~a1266 & a880;
assign a1270 = ~a880 & ~l452;
assign a1272 = ~a1270 & ~a1268;
assign a1276 = ~a1244 & ~l454;
assign a1278 = ~a1276 & a880;
assign a1280 = ~a880 & ~l454;
assign a1282 = ~a1280 & ~a1278;
assign a1286 = l468 & ~l466;
assign a1288 = l488 & l486;
assign a1290 = a1288 & ~l484;
assign a1292 = a1290 & a1286;
assign a1294 = ~l468 & l466;
assign a1296 = a1294 & a1290;
assign a1298 = l488 & ~l486;
assign a1300 = a1298 & l484;
assign a1302 = a1300 & a1294;
assign a1304 = l458 & ~l456;
assign a1306 = a1288 & l484;
assign a1308 = a1306 & a1294;
assign a1310 = a1308 & a1304;
assign a1312 = ~l458 & ~l456;
assign a1314 = l468 & l466;
assign a1316 = a1298 & ~l484;
assign a1318 = a1316 & a1314;
assign a1320 = a1318 & a1312;
assign a1322 = a1316 & a1286;
assign a1324 = a1322 & a1304;
assign a1326 = a1316 & l490;
assign a1328 = ~a1326 & l460;
assign a1330 = a1328 & ~a1324;
assign a1332 = a1330 & ~a1320;
assign a1334 = ~a1332 & ~a1310;
assign a1336 = ~a1334 & ~a1302;
assign a1338 = ~a1336 & ~a1296;
assign a1340 = ~a1338 & ~a1292;
assign a1344 = ~a1326 & l462;
assign a1346 = a1344 & ~a1324;
assign a1348 = a1346 & ~a1320;
assign a1350 = ~a1348 & ~a1310;
assign a1352 = ~a1350 & ~a1302;
assign a1354 = ~a1352 & ~a1296;
assign a1356 = a1354 & ~a1292;
assign a1360 = ~l458 & l456;
assign a1362 = ~l488 & ~l486;
assign a1364 = a1362 & ~l484;
assign a1366 = a1364 & a1294;
assign a1368 = a1366 & a1360;
assign a1370 = ~l488 & l486;
assign a1372 = a1370 & ~l484;
assign a1374 = a1372 & a1294;
assign a1376 = a1374 & a1312;
assign a1378 = a1360 & a1308;
assign a1380 = ~a1378 & ~l468;
assign a1382 = a1380 & ~a1376;
assign a1384 = a1382 & ~a1368;
assign a1388 = l482 & ~l480;
assign a1390 = a1388 & a1290;
assign a1392 = ~l482 & l480;
assign a1394 = a1392 & a1290;
assign a1396 = a1392 & a1300;
assign a1398 = l472 & ~l470;
assign a1400 = a1392 & a1306;
assign a1402 = a1400 & a1398;
assign a1404 = ~l472 & ~l470;
assign a1406 = l482 & l480;
assign a1408 = a1406 & a1316;
assign a1410 = a1408 & a1404;
assign a1412 = a1388 & a1316;
assign a1414 = a1412 & a1398;
assign a1416 = ~a1326 & l474;
assign a1418 = a1416 & ~a1414;
assign a1420 = a1418 & ~a1410;
assign a1422 = ~a1420 & ~a1402;
assign a1424 = ~a1422 & ~a1396;
assign a1426 = ~a1424 & ~a1394;
assign a1428 = ~a1426 & ~a1390;
assign a1432 = ~a1326 & l476;
assign a1434 = a1432 & ~a1414;
assign a1436 = a1434 & ~a1410;
assign a1438 = ~a1436 & ~a1402;
assign a1440 = ~a1438 & ~a1396;
assign a1442 = ~a1440 & ~a1394;
assign a1444 = a1442 & ~a1390;
assign a1448 = ~l472 & l470;
assign a1450 = a1392 & a1364;
assign a1452 = a1450 & a1448;
assign a1454 = a1392 & a1372;
assign a1456 = a1454 & a1404;
assign a1458 = a1448 & a1400;
assign a1460 = ~a1458 & ~l482;
assign a1462 = a1460 & ~a1456;
assign a1464 = a1462 & ~a1452;
assign a1468 = ~l500 & l494;
assign a1470 = a1392 & a1294;
assign a1472 = ~a1470 & a1364;
assign a1474 = a1472 & ~a1468;
assign a1476 = ~a1304 & a1286;
assign a1478 = ~a1476 & a1290;
assign a1480 = ~a1398 & a1388;
assign a1482 = ~a1480 & a1478;
assign a1484 = ~a1312 & a1294;
assign a1486 = ~a1484 & a1372;
assign a1488 = ~a1404 & a1392;
assign a1490 = ~a1488 & a1486;
assign a1492 = ~a1448 & a1392;
assign a1494 = ~a1360 & a1294;
assign a1496 = ~a1494 & a1372;
assign a1498 = a1496 & ~a1492;
assign a1500 = ~a1304 & a1294;
assign a1502 = ~a1398 & a1392;
assign a1504 = ~a1502 & ~a1500;
assign a1506 = ~a1494 & ~a1492;
assign a1508 = ~a1506 & ~a1504;
assign a1510 = ~a1508 & ~a1298;
assign a1512 = a1510 & a1306;
assign a1514 = a1512 & ~a1362;
assign a1516 = ~a1514 & l484;
assign a1518 = ~a1516 & ~a1498;
assign a1520 = ~a1518 & ~a1490;
assign a1522 = a1520 & ~a1482;
assign a1524 = a1522 & ~a1474;
assign a1528 = a1300 & ~l496;
assign a1530 = a1362 & l484;
assign a1532 = l488 & l484;
assign a1534 = a1532 & l496;
assign a1536 = ~a1534 & a1530;
assign a1538 = ~a1536 & ~l486;
assign a1540 = a1538 & ~a1528;
assign a1542 = ~a1540 & ~a1498;
assign a1544 = a1542 & ~a1490;
assign a1546 = ~a1544 & ~a1482;
assign a1548 = a1546 & ~a1474;
assign a1552 = a1300 & l496;
assign a1554 = a1504 & a1306;
assign a1556 = ~a1554 & l488;
assign a1558 = ~a1556 & ~a1530;
assign a1560 = ~a1558 & ~a1552;
assign a1562 = ~a1560 & ~a1528;
assign a1564 = a1562 & ~a1498;
assign a1566 = a1564 & ~a1490;
assign a1568 = ~a1566 & ~a1482;
assign a1570 = ~a1568 & ~a1474;
assign a1574 = ~l506 & ~l504;
assign a1576 = ~a1574 & l502;
assign a1578 = a1576 & l500;
assign a1580 = a1578 & a1364;
assign a1582 = ~a1580 & ~l498;
assign a1586 = ~l504 & ~l502;
assign a1588 = a1586 & ~l500;
assign a1590 = l506 & ~l504;
assign a1592 = a1590 & ~l502;
assign a1594 = a1592 & ~l500;
assign a1596 = l504 & ~l502;
assign a1598 = a1596 & ~l500;
assign a1600 = l506 & l504;
assign a1602 = a1600 & ~l502;
assign a1604 = a1602 & ~l500;
assign a1606 = ~l504 & l502;
assign a1608 = a1606 & ~l500;
assign a1610 = a1590 & l502;
assign a1612 = a1610 & ~l500;
assign a1614 = l504 & l502;
assign a1616 = a1614 & ~l500;
assign a1618 = a1592 & l500;
assign a1620 = a1602 & l500;
assign a1622 = ~a1620 & a1606;
assign a1624 = ~a1622 & ~a1596;
assign a1626 = ~a1624 & ~a1618;
assign a1628 = ~a1626 & ~a1586;
assign a1630 = ~a1628 & l500;
assign a1632 = ~a1630 & ~a1616;
assign a1634 = ~a1632 & ~a1612;
assign a1636 = ~a1634 & ~a1608;
assign a1638 = ~a1636 & ~a1604;
assign a1640 = ~a1638 & ~a1598;
assign a1642 = ~a1640 & ~a1594;
assign a1644 = ~a1642 & ~a1588;
assign a1646 = ~a1644 & ~l506;
assign a1648 = a1574 & ~l502;
assign a1650 = a1648 & ~l500;
assign a1652 = l506 & ~l502;
assign a1654 = a1652 & ~l500;
assign a1656 = a1574 & l502;
assign a1658 = a1656 & ~l500;
assign a1660 = l506 & l502;
assign a1662 = a1660 & ~l500;
assign a1664 = a1648 & l500;
assign a1666 = ~l502 & l500;
assign a1668 = a1666 & ~a1590;
assign a1670 = a1668 & ~a1664;
assign a1672 = ~a1670 & ~a1662;
assign a1674 = ~l506 & l502;
assign a1676 = a1674 & ~l500;
assign a1678 = ~a1676 & a1672;
assign a1680 = ~a1678 & ~a1612;
assign a1682 = a1680 & ~a1658;
assign a1684 = ~a1682 & ~a1654;
assign a1686 = ~l506 & ~l502;
assign a1688 = a1686 & ~l500;
assign a1690 = ~a1688 & a1684;
assign a1692 = ~a1690 & l504;
assign a1694 = a1692 & ~a1594;
assign a1696 = a1694 & ~a1650;
assign a1698 = a1696 & a1646;
assign a1700 = ~l506 & l504;
assign a1702 = ~a1600 & ~l500;
assign a1704 = a1702 & ~a1700;
assign a1706 = a1590 & ~l500;
assign a1708 = ~a1706 & a1704;
assign a1710 = a1574 & ~l500;
assign a1712 = ~a1710 & a1708;
assign a1714 = ~a1712 & ~l502;
assign a1716 = ~a1714 & a1698;
assign a1718 = ~a1600 & ~l502;
assign a1720 = a1718 & ~a1700;
assign a1722 = a1720 & ~a1592;
assign a1724 = a1722 & ~a1648;
assign a1726 = ~a1724 & ~l500;
assign a1728 = ~a1726 & a1716;
assign a1730 = ~a1728 & l500;
assign a1732 = ~a1730 & a1364;
assign a1734 = ~a1364 & ~l500;
assign a1736 = ~a1734 & ~a1732;
assign a1740 = ~a1728 & l502;
assign a1742 = ~a1740 & a1364;
assign a1744 = ~a1364 & ~l502;
assign a1746 = ~a1744 & ~a1742;
assign a1750 = ~a1728 & l504;
assign a1752 = ~a1750 & a1364;
assign a1754 = ~a1364 & ~l504;
assign a1756 = ~a1754 & ~a1752;
assign a1760 = ~a1728 & ~l506;
assign a1762 = ~a1760 & a1364;
assign a1764 = ~a1364 & ~l506;
assign a1766 = ~a1764 & ~a1762;
assign a1770 = l520 & ~l518;
assign a1772 = l540 & l538;
assign a1774 = a1772 & ~l536;
assign a1776 = a1774 & a1770;
assign a1778 = ~l520 & l518;
assign a1780 = a1778 & a1774;
assign a1782 = l540 & ~l538;
assign a1784 = a1782 & l536;
assign a1786 = a1784 & a1778;
assign a1788 = l510 & ~l508;
assign a1790 = a1772 & l536;
assign a1792 = a1790 & a1778;
assign a1794 = a1792 & a1788;
assign a1796 = ~l510 & ~l508;
assign a1798 = l520 & l518;
assign a1800 = a1782 & ~l536;
assign a1802 = a1800 & a1798;
assign a1804 = a1802 & a1796;
assign a1806 = a1800 & a1770;
assign a1808 = a1806 & a1788;
assign a1810 = a1800 & l542;
assign a1812 = ~a1810 & l512;
assign a1814 = a1812 & ~a1808;
assign a1816 = a1814 & ~a1804;
assign a1818 = ~a1816 & ~a1794;
assign a1820 = ~a1818 & ~a1786;
assign a1822 = ~a1820 & ~a1780;
assign a1824 = ~a1822 & ~a1776;
assign a1828 = ~a1810 & l514;
assign a1830 = a1828 & ~a1808;
assign a1832 = a1830 & ~a1804;
assign a1834 = ~a1832 & ~a1794;
assign a1836 = ~a1834 & ~a1786;
assign a1838 = ~a1836 & ~a1780;
assign a1840 = a1838 & ~a1776;
assign a1844 = ~l510 & l508;
assign a1846 = ~l540 & ~l538;
assign a1848 = a1846 & ~l536;
assign a1850 = a1848 & a1778;
assign a1852 = a1850 & a1844;
assign a1854 = ~l540 & l538;
assign a1856 = a1854 & ~l536;
assign a1858 = a1856 & a1778;
assign a1860 = a1858 & a1796;
assign a1862 = a1844 & a1792;
assign a1864 = ~a1862 & ~l520;
assign a1866 = a1864 & ~a1860;
assign a1868 = a1866 & ~a1852;
assign a1872 = l534 & ~l532;
assign a1874 = a1872 & a1774;
assign a1876 = ~l534 & l532;
assign a1878 = a1876 & a1774;
assign a1880 = a1876 & a1784;
assign a1882 = l524 & ~l522;
assign a1884 = a1876 & a1790;
assign a1886 = a1884 & a1882;
assign a1888 = ~l524 & ~l522;
assign a1890 = l534 & l532;
assign a1892 = a1890 & a1800;
assign a1894 = a1892 & a1888;
assign a1896 = a1872 & a1800;
assign a1898 = a1896 & a1882;
assign a1900 = ~a1810 & l526;
assign a1902 = a1900 & ~a1898;
assign a1904 = a1902 & ~a1894;
assign a1906 = ~a1904 & ~a1886;
assign a1908 = ~a1906 & ~a1880;
assign a1910 = ~a1908 & ~a1878;
assign a1912 = ~a1910 & ~a1874;
assign a1916 = ~a1810 & l528;
assign a1918 = a1916 & ~a1898;
assign a1920 = a1918 & ~a1894;
assign a1922 = ~a1920 & ~a1886;
assign a1924 = ~a1922 & ~a1880;
assign a1926 = ~a1924 & ~a1878;
assign a1928 = a1926 & ~a1874;
assign a1932 = ~l524 & l522;
assign a1934 = a1876 & a1848;
assign a1936 = a1934 & a1932;
assign a1938 = a1876 & a1856;
assign a1940 = a1938 & a1888;
assign a1942 = a1932 & a1884;
assign a1944 = ~a1942 & ~l534;
assign a1946 = a1944 & ~a1940;
assign a1948 = a1946 & ~a1936;
assign a1952 = ~l552 & l546;
assign a1954 = a1876 & a1778;
assign a1956 = ~a1954 & a1848;
assign a1958 = a1956 & ~a1952;
assign a1960 = ~a1788 & a1770;
assign a1962 = ~a1960 & a1774;
assign a1964 = ~a1882 & a1872;
assign a1966 = ~a1964 & a1962;
assign a1968 = ~a1796 & a1778;
assign a1970 = ~a1968 & a1856;
assign a1972 = ~a1888 & a1876;
assign a1974 = ~a1972 & a1970;
assign a1976 = ~a1932 & a1876;
assign a1978 = ~a1844 & a1778;
assign a1980 = ~a1978 & a1856;
assign a1982 = a1980 & ~a1976;
assign a1984 = ~a1788 & a1778;
assign a1986 = ~a1882 & a1876;
assign a1988 = ~a1986 & ~a1984;
assign a1990 = ~a1978 & ~a1976;
assign a1992 = ~a1990 & ~a1988;
assign a1994 = ~a1992 & ~a1782;
assign a1996 = a1994 & a1790;
assign a1998 = a1996 & ~a1846;
assign a2000 = ~a1998 & l536;
assign a2002 = ~a2000 & ~a1982;
assign a2004 = ~a2002 & ~a1974;
assign a2006 = a2004 & ~a1966;
assign a2008 = a2006 & ~a1958;
assign a2012 = a1784 & ~l548;
assign a2014 = a1846 & l536;
assign a2016 = l540 & l536;
assign a2018 = a2016 & l548;
assign a2020 = ~a2018 & a2014;
assign a2022 = ~a2020 & ~l538;
assign a2024 = a2022 & ~a2012;
assign a2026 = ~a2024 & ~a1982;
assign a2028 = a2026 & ~a1974;
assign a2030 = ~a2028 & ~a1966;
assign a2032 = a2030 & ~a1958;
assign a2036 = a1784 & l548;
assign a2038 = a1988 & a1790;
assign a2040 = ~a2038 & l540;
assign a2042 = ~a2040 & ~a2014;
assign a2044 = ~a2042 & ~a2036;
assign a2046 = ~a2044 & ~a2012;
assign a2048 = a2046 & ~a1982;
assign a2050 = a2048 & ~a1974;
assign a2052 = ~a2050 & ~a1966;
assign a2054 = ~a2052 & ~a1958;
assign a2058 = ~l558 & ~l556;
assign a2060 = ~a2058 & l554;
assign a2062 = a2060 & l552;
assign a2064 = a2062 & a1848;
assign a2066 = ~a2064 & ~l550;
assign a2070 = ~l556 & ~l554;
assign a2072 = a2070 & ~l552;
assign a2074 = l558 & ~l556;
assign a2076 = a2074 & ~l554;
assign a2078 = a2076 & ~l552;
assign a2080 = l556 & ~l554;
assign a2082 = a2080 & ~l552;
assign a2084 = l558 & l556;
assign a2086 = a2084 & ~l554;
assign a2088 = a2086 & ~l552;
assign a2090 = ~l556 & l554;
assign a2092 = a2090 & ~l552;
assign a2094 = a2074 & l554;
assign a2096 = a2094 & ~l552;
assign a2098 = l556 & l554;
assign a2100 = a2098 & ~l552;
assign a2102 = a2076 & l552;
assign a2104 = a2086 & l552;
assign a2106 = ~a2104 & a2090;
assign a2108 = ~a2106 & ~a2080;
assign a2110 = ~a2108 & ~a2102;
assign a2112 = ~a2110 & ~a2070;
assign a2114 = ~a2112 & l552;
assign a2116 = ~a2114 & ~a2100;
assign a2118 = ~a2116 & ~a2096;
assign a2120 = ~a2118 & ~a2092;
assign a2122 = ~a2120 & ~a2088;
assign a2124 = ~a2122 & ~a2082;
assign a2126 = ~a2124 & ~a2078;
assign a2128 = ~a2126 & ~a2072;
assign a2130 = ~a2128 & ~l558;
assign a2132 = a2058 & ~l554;
assign a2134 = a2132 & ~l552;
assign a2136 = l558 & ~l554;
assign a2138 = a2136 & ~l552;
assign a2140 = a2058 & l554;
assign a2142 = a2140 & ~l552;
assign a2144 = l558 & l554;
assign a2146 = a2144 & ~l552;
assign a2148 = a2132 & l552;
assign a2150 = ~l554 & l552;
assign a2152 = a2150 & ~a2074;
assign a2154 = a2152 & ~a2148;
assign a2156 = ~a2154 & ~a2146;
assign a2158 = ~l558 & l554;
assign a2160 = a2158 & ~l552;
assign a2162 = ~a2160 & a2156;
assign a2164 = ~a2162 & ~a2096;
assign a2166 = a2164 & ~a2142;
assign a2168 = ~a2166 & ~a2138;
assign a2170 = ~l558 & ~l554;
assign a2172 = a2170 & ~l552;
assign a2174 = ~a2172 & a2168;
assign a2176 = ~a2174 & l556;
assign a2178 = a2176 & ~a2078;
assign a2180 = a2178 & ~a2134;
assign a2182 = a2180 & a2130;
assign a2184 = ~l558 & l556;
assign a2186 = ~a2084 & ~l552;
assign a2188 = a2186 & ~a2184;
assign a2190 = a2074 & ~l552;
assign a2192 = ~a2190 & a2188;
assign a2194 = a2058 & ~l552;
assign a2196 = ~a2194 & a2192;
assign a2198 = ~a2196 & ~l554;
assign a2200 = ~a2198 & a2182;
assign a2202 = ~a2084 & ~l554;
assign a2204 = a2202 & ~a2184;
assign a2206 = a2204 & ~a2076;
assign a2208 = a2206 & ~a2132;
assign a2210 = ~a2208 & ~l552;
assign a2212 = ~a2210 & a2200;
assign a2214 = ~a2212 & l552;
assign a2216 = ~a2214 & a1848;
assign a2218 = ~a1848 & ~l552;
assign a2220 = ~a2218 & ~a2216;
assign a2224 = ~a2212 & l554;
assign a2226 = ~a2224 & a1848;
assign a2228 = ~a1848 & ~l554;
assign a2230 = ~a2228 & ~a2226;
assign a2234 = ~a2212 & l556;
assign a2236 = ~a2234 & a1848;
assign a2238 = ~a1848 & ~l556;
assign a2240 = ~a2238 & ~a2236;
assign a2244 = ~a2212 & ~l558;
assign a2246 = ~a2244 & a1848;
assign a2248 = ~a1848 & ~l558;
assign a2250 = ~a2248 & ~a2246;
assign a2254 = l572 & ~l570;
assign a2256 = l592 & l590;
assign a2258 = a2256 & ~l588;
assign a2260 = a2258 & a2254;
assign a2262 = ~l572 & l570;
assign a2264 = a2262 & a2258;
assign a2266 = l592 & ~l590;
assign a2268 = a2266 & l588;
assign a2270 = a2268 & a2262;
assign a2272 = l562 & ~l560;
assign a2274 = a2256 & l588;
assign a2276 = a2274 & a2262;
assign a2278 = a2276 & a2272;
assign a2280 = ~l562 & ~l560;
assign a2282 = l572 & l570;
assign a2284 = a2266 & ~l588;
assign a2286 = a2284 & a2282;
assign a2288 = a2286 & a2280;
assign a2290 = a2284 & a2254;
assign a2292 = a2290 & a2272;
assign a2294 = a2284 & l594;
assign a2296 = ~a2294 & l564;
assign a2298 = a2296 & ~a2292;
assign a2300 = a2298 & ~a2288;
assign a2302 = ~a2300 & ~a2278;
assign a2304 = ~a2302 & ~a2270;
assign a2306 = ~a2304 & ~a2264;
assign a2308 = ~a2306 & ~a2260;
assign a2312 = ~a2294 & l566;
assign a2314 = a2312 & ~a2292;
assign a2316 = a2314 & ~a2288;
assign a2318 = ~a2316 & ~a2278;
assign a2320 = ~a2318 & ~a2270;
assign a2322 = ~a2320 & ~a2264;
assign a2324 = a2322 & ~a2260;
assign a2328 = ~l562 & l560;
assign a2330 = ~l592 & ~l590;
assign a2332 = a2330 & ~l588;
assign a2334 = a2332 & a2262;
assign a2336 = a2334 & a2328;
assign a2338 = ~l592 & l590;
assign a2340 = a2338 & ~l588;
assign a2342 = a2340 & a2262;
assign a2344 = a2342 & a2280;
assign a2346 = a2328 & a2276;
assign a2348 = ~a2346 & ~l572;
assign a2350 = a2348 & ~a2344;
assign a2352 = a2350 & ~a2336;
assign a2356 = l586 & ~l584;
assign a2358 = a2356 & a2258;
assign a2360 = ~l586 & l584;
assign a2362 = a2360 & a2258;
assign a2364 = a2360 & a2268;
assign a2366 = l576 & ~l574;
assign a2368 = a2360 & a2274;
assign a2370 = a2368 & a2366;
assign a2372 = ~l576 & ~l574;
assign a2374 = l586 & l584;
assign a2376 = a2374 & a2284;
assign a2378 = a2376 & a2372;
assign a2380 = a2356 & a2284;
assign a2382 = a2380 & a2366;
assign a2384 = ~a2294 & l578;
assign a2386 = a2384 & ~a2382;
assign a2388 = a2386 & ~a2378;
assign a2390 = ~a2388 & ~a2370;
assign a2392 = ~a2390 & ~a2364;
assign a2394 = ~a2392 & ~a2362;
assign a2396 = ~a2394 & ~a2358;
assign a2400 = ~a2294 & l580;
assign a2402 = a2400 & ~a2382;
assign a2404 = a2402 & ~a2378;
assign a2406 = ~a2404 & ~a2370;
assign a2408 = ~a2406 & ~a2364;
assign a2410 = ~a2408 & ~a2362;
assign a2412 = a2410 & ~a2358;
assign a2416 = ~l576 & l574;
assign a2418 = a2360 & a2332;
assign a2420 = a2418 & a2416;
assign a2422 = a2360 & a2340;
assign a2424 = a2422 & a2372;
assign a2426 = a2416 & a2368;
assign a2428 = ~a2426 & ~l586;
assign a2430 = a2428 & ~a2424;
assign a2432 = a2430 & ~a2420;
assign a2436 = ~l604 & l598;
assign a2438 = a2360 & a2262;
assign a2440 = ~a2438 & a2332;
assign a2442 = a2440 & ~a2436;
assign a2444 = ~a2272 & a2254;
assign a2446 = ~a2444 & a2258;
assign a2448 = ~a2366 & a2356;
assign a2450 = ~a2448 & a2446;
assign a2452 = ~a2280 & a2262;
assign a2454 = ~a2452 & a2340;
assign a2456 = ~a2372 & a2360;
assign a2458 = ~a2456 & a2454;
assign a2460 = ~a2416 & a2360;
assign a2462 = ~a2328 & a2262;
assign a2464 = ~a2462 & a2340;
assign a2466 = a2464 & ~a2460;
assign a2468 = ~a2272 & a2262;
assign a2470 = ~a2366 & a2360;
assign a2472 = ~a2470 & ~a2468;
assign a2474 = ~a2462 & ~a2460;
assign a2476 = ~a2474 & ~a2472;
assign a2478 = ~a2476 & ~a2266;
assign a2480 = a2478 & a2274;
assign a2482 = a2480 & ~a2330;
assign a2484 = ~a2482 & l588;
assign a2486 = ~a2484 & ~a2466;
assign a2488 = ~a2486 & ~a2458;
assign a2490 = a2488 & ~a2450;
assign a2492 = a2490 & ~a2442;
assign a2496 = a2268 & ~l600;
assign a2498 = a2330 & l588;
assign a2500 = l592 & l588;
assign a2502 = a2500 & l600;
assign a2504 = ~a2502 & a2498;
assign a2506 = ~a2504 & ~l590;
assign a2508 = a2506 & ~a2496;
assign a2510 = ~a2508 & ~a2466;
assign a2512 = a2510 & ~a2458;
assign a2514 = ~a2512 & ~a2450;
assign a2516 = a2514 & ~a2442;
assign a2520 = a2268 & l600;
assign a2522 = a2472 & a2274;
assign a2524 = ~a2522 & l592;
assign a2526 = ~a2524 & ~a2498;
assign a2528 = ~a2526 & ~a2520;
assign a2530 = ~a2528 & ~a2496;
assign a2532 = a2530 & ~a2466;
assign a2534 = a2532 & ~a2458;
assign a2536 = ~a2534 & ~a2450;
assign a2538 = ~a2536 & ~a2442;
assign a2542 = ~l610 & ~l608;
assign a2544 = ~a2542 & l606;
assign a2546 = a2544 & l604;
assign a2548 = a2546 & a2332;
assign a2550 = ~a2548 & ~l602;
assign a2554 = ~l608 & ~l606;
assign a2556 = a2554 & ~l604;
assign a2558 = l610 & ~l608;
assign a2560 = a2558 & ~l606;
assign a2562 = a2560 & ~l604;
assign a2564 = l608 & ~l606;
assign a2566 = a2564 & ~l604;
assign a2568 = l610 & l608;
assign a2570 = a2568 & ~l606;
assign a2572 = a2570 & ~l604;
assign a2574 = ~l608 & l606;
assign a2576 = a2574 & ~l604;
assign a2578 = a2558 & l606;
assign a2580 = a2578 & ~l604;
assign a2582 = l608 & l606;
assign a2584 = a2582 & ~l604;
assign a2586 = a2560 & l604;
assign a2588 = a2570 & l604;
assign a2590 = ~a2588 & a2574;
assign a2592 = ~a2590 & ~a2564;
assign a2594 = ~a2592 & ~a2586;
assign a2596 = ~a2594 & ~a2554;
assign a2598 = ~a2596 & l604;
assign a2600 = ~a2598 & ~a2584;
assign a2602 = ~a2600 & ~a2580;
assign a2604 = ~a2602 & ~a2576;
assign a2606 = ~a2604 & ~a2572;
assign a2608 = ~a2606 & ~a2566;
assign a2610 = ~a2608 & ~a2562;
assign a2612 = ~a2610 & ~a2556;
assign a2614 = ~a2612 & ~l610;
assign a2616 = a2542 & ~l606;
assign a2618 = a2616 & ~l604;
assign a2620 = l610 & ~l606;
assign a2622 = a2620 & ~l604;
assign a2624 = a2542 & l606;
assign a2626 = a2624 & ~l604;
assign a2628 = l610 & l606;
assign a2630 = a2628 & ~l604;
assign a2632 = a2616 & l604;
assign a2634 = ~l606 & l604;
assign a2636 = a2634 & ~a2558;
assign a2638 = a2636 & ~a2632;
assign a2640 = ~a2638 & ~a2630;
assign a2642 = ~l610 & l606;
assign a2644 = a2642 & ~l604;
assign a2646 = ~a2644 & a2640;
assign a2648 = ~a2646 & ~a2580;
assign a2650 = a2648 & ~a2626;
assign a2652 = ~a2650 & ~a2622;
assign a2654 = ~l610 & ~l606;
assign a2656 = a2654 & ~l604;
assign a2658 = ~a2656 & a2652;
assign a2660 = ~a2658 & l608;
assign a2662 = a2660 & ~a2562;
assign a2664 = a2662 & ~a2618;
assign a2666 = a2664 & a2614;
assign a2668 = ~l610 & l608;
assign a2670 = ~a2568 & ~l604;
assign a2672 = a2670 & ~a2668;
assign a2674 = a2558 & ~l604;
assign a2676 = ~a2674 & a2672;
assign a2678 = a2542 & ~l604;
assign a2680 = ~a2678 & a2676;
assign a2682 = ~a2680 & ~l606;
assign a2684 = ~a2682 & a2666;
assign a2686 = ~a2568 & ~l606;
assign a2688 = a2686 & ~a2668;
assign a2690 = a2688 & ~a2560;
assign a2692 = a2690 & ~a2616;
assign a2694 = ~a2692 & ~l604;
assign a2696 = ~a2694 & a2684;
assign a2698 = ~a2696 & l604;
assign a2700 = ~a2698 & a2332;
assign a2702 = ~a2332 & ~l604;
assign a2704 = ~a2702 & ~a2700;
assign a2708 = ~a2696 & l606;
assign a2710 = ~a2708 & a2332;
assign a2712 = ~a2332 & ~l606;
assign a2714 = ~a2712 & ~a2710;
assign a2718 = ~a2696 & l608;
assign a2720 = ~a2718 & a2332;
assign a2722 = ~a2332 & ~l608;
assign a2724 = ~a2722 & ~a2720;
assign a2728 = ~a2696 & ~l610;
assign a2730 = ~a2728 & a2332;
assign a2732 = ~a2332 & ~l610;
assign a2734 = ~a2732 & ~a2730;
assign a2738 = ~a1530 & l614;
assign a2740 = ~a2738 & ~a1046;
assign a2744 = ~l788 & ~l786;
assign a2746 = ~a2744 & l612;
assign a2748 = ~a2746 & ~l780;
assign a2752 = ~l616 & l490;
assign a2754 = ~a2752 & l618;
assign a2756 = ~a2754 & ~a2744;
assign a2758 = ~a2756 & ~l782;
assign a2762 = l616 & l490;
assign a2764 = ~a2762 & ~a2744;
assign a2766 = ~a2764 & ~l784;
assign a2772 = ~l616 & ~l490;
assign a2774 = l612 & ~i162;
assign a2776 = a2752 & ~l618;
assign a2778 = ~a2776 & ~a2774;
assign a2780 = a2778 & ~a2772;
assign a2782 = l340 & ~i2;
assign a2784 = ~l340 & i2;
assign a2786 = ~a2784 & ~a2782;
assign a2788 = a2786 & a2780;
assign a2790 = l342 & ~i4;
assign a2792 = ~l342 & i4;
assign a2794 = ~a2792 & ~a2790;
assign a2796 = a2794 & a2788;
assign a2798 = l344 & ~i6;
assign a2800 = ~l344 & i6;
assign a2802 = ~a2800 & ~a2798;
assign a2804 = a2802 & a2796;
assign a2806 = l346 & ~i8;
assign a2808 = ~l346 & i8;
assign a2810 = ~a2808 & ~a2806;
assign a2812 = a2810 & a2804;
assign a2814 = l348 & ~i10;
assign a2816 = ~l348 & i10;
assign a2818 = ~a2816 & ~a2814;
assign a2820 = a2818 & a2812;
assign a2822 = l350 & ~i12;
assign a2824 = ~l350 & i12;
assign a2826 = ~a2824 & ~a2822;
assign a2828 = a2826 & a2820;
assign a2830 = l352 & ~i14;
assign a2832 = ~l352 & i14;
assign a2834 = ~a2832 & ~a2830;
assign a2836 = a2834 & a2828;
assign a2838 = l354 & ~i16;
assign a2840 = ~l354 & i16;
assign a2842 = ~a2840 & ~a2838;
assign a2844 = a2842 & a2836;
assign a2846 = l356 & ~i18;
assign a2848 = ~l356 & i18;
assign a2850 = ~a2848 & ~a2846;
assign a2852 = a2850 & a2844;
assign a2854 = l358 & ~i20;
assign a2856 = ~l358 & i20;
assign a2858 = ~a2856 & ~a2854;
assign a2860 = a2858 & a2852;
assign a2862 = l360 & ~i22;
assign a2864 = ~l360 & i22;
assign a2866 = ~a2864 & ~a2862;
assign a2868 = a2866 & a2860;
assign a2870 = l362 & ~i24;
assign a2872 = ~l362 & i24;
assign a2874 = ~a2872 & ~a2870;
assign a2876 = a2874 & a2868;
assign a2878 = l364 & ~i26;
assign a2880 = ~l364 & i26;
assign a2882 = ~a2880 & ~a2878;
assign a2884 = a2882 & a2876;
assign a2886 = l366 & ~i28;
assign a2888 = ~l366 & i28;
assign a2890 = ~a2888 & ~a2886;
assign a2892 = a2890 & a2884;
assign a2894 = l368 & ~i30;
assign a2896 = ~l368 & i30;
assign a2898 = ~a2896 & ~a2894;
assign a2900 = a2898 & a2892;
assign a2902 = l370 & ~i32;
assign a2904 = ~l370 & i32;
assign a2906 = ~a2904 & ~a2902;
assign a2908 = a2906 & a2900;
assign a2910 = l372 & ~i34;
assign a2912 = ~l372 & i34;
assign a2914 = ~a2912 & ~a2910;
assign a2916 = a2914 & a2908;
assign a2918 = l374 & ~i36;
assign a2920 = ~l374 & i36;
assign a2922 = ~a2920 & ~a2918;
assign a2924 = a2922 & a2916;
assign a2926 = l376 & ~i38;
assign a2928 = ~l376 & i38;
assign a2930 = ~a2928 & ~a2926;
assign a2932 = a2930 & a2924;
assign a2934 = l378 & ~i40;
assign a2936 = ~l378 & i40;
assign a2938 = ~a2936 & ~a2934;
assign a2940 = a2938 & a2932;
assign a2942 = l380 & ~i42;
assign a2944 = ~l380 & i42;
assign a2946 = ~a2944 & ~a2942;
assign a2948 = a2946 & a2940;
assign a2950 = l382 & ~i44;
assign a2952 = ~l382 & i44;
assign a2954 = ~a2952 & ~a2950;
assign a2956 = a2954 & a2948;
assign a2958 = l384 & ~i46;
assign a2960 = ~l384 & i46;
assign a2962 = ~a2960 & ~a2958;
assign a2964 = a2962 & a2956;
assign a2966 = l386 & ~i48;
assign a2968 = ~l386 & i48;
assign a2970 = ~a2968 & ~a2966;
assign a2972 = a2970 & a2964;
assign a2974 = l388 & ~i50;
assign a2976 = ~l388 & i50;
assign a2978 = ~a2976 & ~a2974;
assign a2980 = a2978 & a2972;
assign a2982 = l390 & ~i52;
assign a2984 = ~l390 & i52;
assign a2986 = ~a2984 & ~a2982;
assign a2988 = a2986 & a2980;
assign a2990 = l392 & ~i54;
assign a2992 = ~l392 & i54;
assign a2994 = ~a2992 & ~a2990;
assign a2996 = a2994 & a2988;
assign a2998 = l394 & ~i56;
assign a3000 = ~l394 & i56;
assign a3002 = ~a3000 & ~a2998;
assign a3004 = a3002 & a2996;
assign a3006 = l396 & ~i58;
assign a3008 = ~l396 & i58;
assign a3010 = ~a3008 & ~a3006;
assign a3012 = a3010 & a3004;
assign a3014 = l398 & ~i60;
assign a3016 = ~l398 & i60;
assign a3018 = ~a3016 & ~a3014;
assign a3020 = a3018 & a3012;
assign a3022 = l400 & ~i62;
assign a3024 = ~l400 & i62;
assign a3026 = ~a3024 & ~a3022;
assign a3028 = a3026 & a3020;
assign a3030 = l402 & ~i64;
assign a3032 = ~l402 & i64;
assign a3034 = ~a3032 & ~a3030;
assign a3036 = a3034 & a3028;
assign a3038 = l412 & ~i70;
assign a3040 = ~l412 & i70;
assign a3042 = ~a3040 & ~a3038;
assign a3044 = a3042 & a3036;
assign a3046 = a888 & ~l416;
assign a3048 = a3046 & a828;
assign a3050 = ~a3048 & a894;
assign a3052 = ~a3050 & l414;
assign a3054 = a3052 & ~a884;
assign a3056 = a3054 & ~i72;
assign a3058 = ~a3054 & i72;
assign a3060 = ~a3058 & ~a3056;
assign a3062 = a3060 & a3044;
assign a3064 = l426 & ~i78;
assign a3066 = ~l426 & i78;
assign a3068 = ~a3066 & ~a3064;
assign a3070 = a3068 & a3062;
assign a3072 = a888 & ~l430;
assign a3074 = a3072 & a920;
assign a3076 = ~a3074 & a974;
assign a3078 = ~a3076 & l428;
assign a3080 = a3078 & ~a968;
assign a3082 = a3080 & ~i80;
assign a3084 = ~a3080 & i80;
assign a3086 = ~a3084 & ~a3082;
assign a3088 = a3086 & a3070;
assign a3090 = ~a908 & ~a810;
assign a3092 = ~a3090 & a806;
assign a3094 = ~a806 & ~l438;
assign a3096 = ~a3094 & ~a3092;
assign a3098 = a3096 & ~i82;
assign a3100 = ~a3096 & i82;
assign a3102 = ~a3100 & ~a3098;
assign a3104 = a3102 & a3088;
assign a3106 = ~a910 & ~l440;
assign a3108 = ~a3106 & ~a812;
assign a3110 = a3108 & ~i84;
assign a3112 = ~a3108 & i84;
assign a3114 = ~a3112 & ~a3110;
assign a3116 = a3114 & a3104;
assign a3118 = l442 & ~i86;
assign a3120 = ~l442 & i86;
assign a3122 = ~a3120 & ~a3118;
assign a3124 = a3122 & a3116;
assign a3126 = a888 & l790;
assign a3128 = ~a888 & ~l444;
assign a3130 = ~a3128 & ~a3126;
assign a3132 = a3130 & ~i88;
assign a3134 = ~a3130 & i88;
assign a3136 = ~a3134 & ~a3132;
assign a3138 = a3136 & a3124;
assign a3140 = l464 & ~i94;
assign a3142 = ~l464 & i94;
assign a3144 = ~a3142 & ~a3140;
assign a3146 = a3144 & a3138;
assign a3148 = a1372 & ~l468;
assign a3150 = a3148 & a1312;
assign a3152 = ~a3150 & a1378;
assign a3154 = ~a3152 & l466;
assign a3156 = a3154 & ~a1368;
assign a3158 = a3156 & ~i96;
assign a3160 = ~a3156 & i96;
assign a3162 = ~a3160 & ~a3158;
assign a3164 = a3162 & a3146;
assign a3166 = l478 & ~i102;
assign a3168 = ~l478 & i102;
assign a3170 = ~a3168 & ~a3166;
assign a3172 = a3170 & a3164;
assign a3174 = a1372 & ~l482;
assign a3176 = a3174 & a1404;
assign a3178 = ~a3176 & a1458;
assign a3180 = ~a3178 & l480;
assign a3182 = a3180 & ~a1452;
assign a3184 = a3182 & ~i104;
assign a3186 = ~a3182 & i104;
assign a3188 = ~a3186 & ~a3184;
assign a3190 = a3188 & a3172;
assign a3192 = ~a1392 & ~a1294;
assign a3194 = ~a3192 & a1290;
assign a3196 = ~a1290 & ~l490;
assign a3198 = ~a3196 & ~a3194;
assign a3200 = a3198 & ~i106;
assign a3202 = ~a3198 & i106;
assign a3204 = ~a3202 & ~a3200;
assign a3206 = a3204 & a3190;
assign a3208 = ~a1394 & ~l492;
assign a3210 = ~a3208 & ~a1296;
assign a3212 = a3210 & ~i108;
assign a3214 = ~a3210 & i108;
assign a3216 = ~a3214 & ~a3212;
assign a3218 = a3216 & a3206;
assign a3220 = l494 & ~i110;
assign a3222 = ~l494 & i110;
assign a3224 = ~a3222 & ~a3220;
assign a3226 = a3224 & a3218;
assign a3228 = a1372 & l792;
assign a3230 = ~a1372 & ~l496;
assign a3232 = ~a3230 & ~a3228;
assign a3234 = a3232 & ~i112;
assign a3236 = ~a3232 & i112;
assign a3238 = ~a3236 & ~a3234;
assign a3240 = a3238 & a3226;
assign a3242 = l516 & ~i118;
assign a3244 = ~l516 & i118;
assign a3246 = ~a3244 & ~a3242;
assign a3248 = a3246 & a3240;
assign a3250 = a1856 & ~l520;
assign a3252 = a3250 & a1796;
assign a3254 = ~a3252 & a1862;
assign a3256 = ~a3254 & l518;
assign a3258 = a3256 & ~a1852;
assign a3260 = a3258 & ~i120;
assign a3262 = ~a3258 & i120;
assign a3264 = ~a3262 & ~a3260;
assign a3266 = a3264 & a3248;
assign a3268 = l530 & ~i126;
assign a3270 = ~l530 & i126;
assign a3272 = ~a3270 & ~a3268;
assign a3274 = a3272 & a3266;
assign a3276 = a1856 & ~l534;
assign a3278 = a3276 & a1888;
assign a3280 = ~a3278 & a1942;
assign a3282 = ~a3280 & l532;
assign a3284 = a3282 & ~a1936;
assign a3286 = a3284 & ~i128;
assign a3288 = ~a3284 & i128;
assign a3290 = ~a3288 & ~a3286;
assign a3292 = a3290 & a3274;
assign a3294 = ~a1876 & ~a1778;
assign a3296 = ~a3294 & a1774;
assign a3298 = ~a1774 & ~l542;
assign a3300 = ~a3298 & ~a3296;
assign a3302 = a3300 & ~i130;
assign a3304 = ~a3300 & i130;
assign a3306 = ~a3304 & ~a3302;
assign a3308 = a3306 & a3292;
assign a3310 = ~a1878 & ~l544;
assign a3312 = ~a3310 & ~a1780;
assign a3314 = a3312 & ~i132;
assign a3316 = ~a3312 & i132;
assign a3318 = ~a3316 & ~a3314;
assign a3320 = a3318 & a3308;
assign a3322 = l546 & ~i134;
assign a3324 = ~l546 & i134;
assign a3326 = ~a3324 & ~a3322;
assign a3328 = a3326 & a3320;
assign a3330 = a1856 & l794;
assign a3332 = ~a1856 & ~l548;
assign a3334 = ~a3332 & ~a3330;
assign a3336 = a3334 & ~i136;
assign a3338 = ~a3334 & i136;
assign a3340 = ~a3338 & ~a3336;
assign a3342 = a3340 & a3328;
assign a3344 = l568 & ~i142;
assign a3346 = ~l568 & i142;
assign a3348 = ~a3346 & ~a3344;
assign a3350 = a3348 & a3342;
assign a3352 = a2340 & ~l572;
assign a3354 = a3352 & a2280;
assign a3356 = ~a3354 & a2346;
assign a3358 = ~a3356 & l570;
assign a3360 = a3358 & ~a2336;
assign a3362 = a3360 & ~i144;
assign a3364 = ~a3360 & i144;
assign a3366 = ~a3364 & ~a3362;
assign a3368 = a3366 & a3350;
assign a3370 = l582 & ~i150;
assign a3372 = ~l582 & i150;
assign a3374 = ~a3372 & ~a3370;
assign a3376 = a3374 & a3368;
assign a3378 = a2340 & ~l586;
assign a3380 = a3378 & a2372;
assign a3382 = ~a3380 & a2426;
assign a3384 = ~a3382 & l584;
assign a3386 = a3384 & ~a2420;
assign a3388 = a3386 & ~i152;
assign a3390 = ~a3386 & i152;
assign a3392 = ~a3390 & ~a3388;
assign a3394 = a3392 & a3376;
assign a3396 = ~a2360 & ~a2262;
assign a3398 = ~a3396 & a2258;
assign a3400 = ~a2258 & ~l594;
assign a3402 = ~a3400 & ~a3398;
assign a3404 = a3402 & ~i154;
assign a3406 = ~a3402 & i154;
assign a3408 = ~a3406 & ~a3404;
assign a3410 = a3408 & a3394;
assign a3412 = ~a2362 & ~l596;
assign a3414 = ~a3412 & ~a2264;
assign a3416 = a3414 & ~i156;
assign a3418 = ~a3414 & i156;
assign a3420 = ~a3418 & ~a3416;
assign a3422 = a3420 & a3410;
assign a3424 = l598 & ~i158;
assign a3426 = ~l598 & i158;
assign a3428 = ~a3426 & ~a3424;
assign a3430 = a3428 & a3422;
assign a3432 = a2340 & l796;
assign a3434 = ~a2340 & ~l600;
assign a3436 = ~a3434 & ~a3432;
assign a3438 = a3436 & ~i160;
assign a3440 = ~a3436 & i160;
assign a3442 = ~a3440 & ~a3438;
assign a3444 = a3442 & a3430;
assign a3446 = ~l788 & l786;
assign a3448 = a3446 & ~l408;
assign a3450 = ~a3446 & ~l620;
assign a3452 = ~a3450 & ~a3448;
assign a3454 = a3452 & ~i168;
assign a3456 = ~a3452 & i168;
assign a3458 = ~a3456 & ~a3454;
assign a3460 = a3458 & a3444;
assign a3462 = ~a3446 & ~l622;
assign a3464 = a3446 & l410;
assign a3466 = ~a3464 & ~a3462;
assign a3468 = a3466 & ~i170;
assign a3470 = ~a3466 & i170;
assign a3472 = ~a3470 & ~a3468;
assign a3474 = a3472 & a3460;
assign a3476 = a3446 & ~l414;
assign a3478 = ~a3446 & ~l624;
assign a3480 = ~a3478 & ~a3476;
assign a3482 = a3480 & ~i172;
assign a3484 = ~a3480 & i172;
assign a3486 = ~a3484 & ~a3482;
assign a3488 = a3486 & a3474;
assign a3490 = ~a3446 & ~l626;
assign a3492 = a3446 & l416;
assign a3494 = ~a3492 & ~a3490;
assign a3496 = a3494 & ~i174;
assign a3498 = ~a3494 & i174;
assign a3500 = ~a3498 & ~a3496;
assign a3502 = a3500 & a3488;
assign a3504 = a3446 & ~l422;
assign a3506 = ~a3446 & ~l628;
assign a3508 = ~a3506 & ~a3504;
assign a3510 = a3508 & ~i176;
assign a3512 = ~a3508 & i176;
assign a3514 = ~a3512 & ~a3510;
assign a3516 = a3514 & a3502;
assign a3518 = ~a3446 & ~l630;
assign a3520 = a3446 & l424;
assign a3522 = ~a3520 & ~a3518;
assign a3524 = a3522 & ~i178;
assign a3526 = ~a3522 & i178;
assign a3528 = ~a3526 & ~a3524;
assign a3530 = a3528 & a3516;
assign a3532 = a3446 & ~l428;
assign a3534 = ~a3446 & ~l632;
assign a3536 = ~a3534 & ~a3532;
assign a3538 = a3536 & ~i180;
assign a3540 = ~a3536 & i180;
assign a3542 = ~a3540 & ~a3538;
assign a3544 = a3542 & a3530;
assign a3546 = ~a3446 & ~l634;
assign a3548 = a3446 & l430;
assign a3550 = ~a3548 & ~a3546;
assign a3552 = a3550 & ~i182;
assign a3554 = ~a3550 & i182;
assign a3556 = ~a3554 & ~a3552;
assign a3558 = a3556 & a3544;
assign a3560 = a3446 & ~l432;
assign a3562 = ~a3446 & ~l636;
assign a3564 = ~a3562 & ~a3560;
assign a3566 = a3564 & ~i184;
assign a3568 = ~a3564 & i184;
assign a3570 = ~a3568 & ~a3566;
assign a3572 = a3570 & a3558;
assign a3574 = a3446 & ~l434;
assign a3576 = ~a3446 & ~l638;
assign a3578 = ~a3576 & ~a3574;
assign a3580 = a3578 & ~i186;
assign a3582 = ~a3578 & i186;
assign a3584 = ~a3582 & ~a3580;
assign a3586 = a3584 & a3572;
assign a3588 = ~a3446 & ~l640;
assign a3590 = a3446 & l436;
assign a3592 = ~a3590 & ~a3588;
assign a3594 = a3592 & ~i188;
assign a3596 = ~a3592 & i188;
assign a3598 = ~a3596 & ~a3594;
assign a3600 = a3598 & a3586;
assign a3602 = a3446 & ~l438;
assign a3604 = ~a3446 & ~l642;
assign a3606 = ~a3604 & ~a3602;
assign a3608 = a3606 & ~i190;
assign a3610 = ~a3606 & i190;
assign a3612 = ~a3610 & ~a3608;
assign a3614 = a3612 & a3600;
assign a3616 = a3446 & ~l440;
assign a3618 = ~a3446 & ~l644;
assign a3620 = ~a3618 & ~a3616;
assign a3622 = a3620 & ~i192;
assign a3624 = ~a3620 & i192;
assign a3626 = ~a3624 & ~a3622;
assign a3628 = a3626 & a3614;
assign a3630 = a3446 & ~l444;
assign a3632 = ~a3446 & ~l646;
assign a3634 = ~a3632 & ~a3630;
assign a3636 = a3634 & ~i194;
assign a3638 = ~a3634 & i194;
assign a3640 = ~a3638 & ~a3636;
assign a3642 = a3640 & a3628;
assign a3644 = a3446 & ~l446;
assign a3646 = ~a3446 & ~l648;
assign a3648 = ~a3646 & ~a3644;
assign a3650 = a3648 & ~i196;
assign a3652 = ~a3648 & i196;
assign a3654 = ~a3652 & ~a3650;
assign a3656 = a3654 & a3642;
assign a3658 = a3446 & ~l448;
assign a3660 = ~a3446 & ~l650;
assign a3662 = ~a3660 & ~a3658;
assign a3664 = a3662 & ~i198;
assign a3666 = ~a3662 & i198;
assign a3668 = ~a3666 & ~a3664;
assign a3670 = a3668 & a3656;
assign a3672 = a3446 & ~l450;
assign a3674 = ~a3446 & ~l652;
assign a3676 = ~a3674 & ~a3672;
assign a3678 = a3676 & ~i200;
assign a3680 = ~a3676 & i200;
assign a3682 = ~a3680 & ~a3678;
assign a3684 = a3682 & a3670;
assign a3686 = a3446 & ~l452;
assign a3688 = ~a3446 & ~l654;
assign a3690 = ~a3688 & ~a3686;
assign a3692 = a3690 & ~i202;
assign a3694 = ~a3690 & i202;
assign a3696 = ~a3694 & ~a3692;
assign a3698 = a3696 & a3684;
assign a3700 = a3446 & ~l454;
assign a3702 = ~a3446 & ~l656;
assign a3704 = ~a3702 & ~a3700;
assign a3706 = a3704 & ~i204;
assign a3708 = ~a3704 & i204;
assign a3710 = ~a3708 & ~a3706;
assign a3712 = a3710 & a3698;
assign a3714 = a3446 & ~l460;
assign a3716 = ~a3446 & ~l658;
assign a3718 = ~a3716 & ~a3714;
assign a3720 = a3718 & ~i206;
assign a3722 = ~a3718 & i206;
assign a3724 = ~a3722 & ~a3720;
assign a3726 = a3724 & a3712;
assign a3728 = ~a3446 & ~l660;
assign a3730 = a3446 & l462;
assign a3732 = ~a3730 & ~a3728;
assign a3734 = a3732 & ~i208;
assign a3736 = ~a3732 & i208;
assign a3738 = ~a3736 & ~a3734;
assign a3740 = a3738 & a3726;
assign a3742 = a3446 & ~l466;
assign a3744 = ~a3446 & ~l662;
assign a3746 = ~a3744 & ~a3742;
assign a3748 = a3746 & ~i210;
assign a3750 = ~a3746 & i210;
assign a3752 = ~a3750 & ~a3748;
assign a3754 = a3752 & a3740;
assign a3756 = ~a3446 & ~l664;
assign a3758 = a3446 & l468;
assign a3760 = ~a3758 & ~a3756;
assign a3762 = a3760 & ~i212;
assign a3764 = ~a3760 & i212;
assign a3766 = ~a3764 & ~a3762;
assign a3768 = a3766 & a3754;
assign a3770 = a3446 & ~l474;
assign a3772 = ~a3446 & ~l666;
assign a3774 = ~a3772 & ~a3770;
assign a3776 = a3774 & ~i214;
assign a3778 = ~a3774 & i214;
assign a3780 = ~a3778 & ~a3776;
assign a3782 = a3780 & a3768;
assign a3784 = ~a3446 & ~l668;
assign a3786 = a3446 & l476;
assign a3788 = ~a3786 & ~a3784;
assign a3790 = a3788 & ~i216;
assign a3792 = ~a3788 & i216;
assign a3794 = ~a3792 & ~a3790;
assign a3796 = a3794 & a3782;
assign a3798 = a3446 & ~l480;
assign a3800 = ~a3446 & ~l670;
assign a3802 = ~a3800 & ~a3798;
assign a3804 = a3802 & ~i218;
assign a3806 = ~a3802 & i218;
assign a3808 = ~a3806 & ~a3804;
assign a3810 = a3808 & a3796;
assign a3812 = ~a3446 & ~l672;
assign a3814 = a3446 & l482;
assign a3816 = ~a3814 & ~a3812;
assign a3818 = a3816 & ~i220;
assign a3820 = ~a3816 & i220;
assign a3822 = ~a3820 & ~a3818;
assign a3824 = a3822 & a3810;
assign a3826 = a3446 & ~l484;
assign a3828 = ~a3446 & ~l674;
assign a3830 = ~a3828 & ~a3826;
assign a3832 = a3830 & ~i222;
assign a3834 = ~a3830 & i222;
assign a3836 = ~a3834 & ~a3832;
assign a3838 = a3836 & a3824;
assign a3840 = a3446 & ~l486;
assign a3842 = ~a3446 & ~l676;
assign a3844 = ~a3842 & ~a3840;
assign a3846 = a3844 & ~i224;
assign a3848 = ~a3844 & i224;
assign a3850 = ~a3848 & ~a3846;
assign a3852 = a3850 & a3838;
assign a3854 = ~a3446 & ~l678;
assign a3856 = a3446 & l488;
assign a3858 = ~a3856 & ~a3854;
assign a3860 = a3858 & ~i226;
assign a3862 = ~a3858 & i226;
assign a3864 = ~a3862 & ~a3860;
assign a3866 = a3864 & a3852;
assign a3868 = a3446 & ~l490;
assign a3870 = ~a3446 & ~l680;
assign a3872 = ~a3870 & ~a3868;
assign a3874 = a3872 & ~i228;
assign a3876 = ~a3872 & i228;
assign a3878 = ~a3876 & ~a3874;
assign a3880 = a3878 & a3866;
assign a3882 = a3446 & ~l492;
assign a3884 = ~a3446 & ~l682;
assign a3886 = ~a3884 & ~a3882;
assign a3888 = a3886 & ~i230;
assign a3890 = ~a3886 & i230;
assign a3892 = ~a3890 & ~a3888;
assign a3894 = a3892 & a3880;
assign a3896 = a3446 & ~l496;
assign a3898 = ~a3446 & ~l684;
assign a3900 = ~a3898 & ~a3896;
assign a3902 = a3900 & ~i232;
assign a3904 = ~a3900 & i232;
assign a3906 = ~a3904 & ~a3902;
assign a3908 = a3906 & a3894;
assign a3910 = a3446 & ~l498;
assign a3912 = ~a3446 & ~l686;
assign a3914 = ~a3912 & ~a3910;
assign a3916 = a3914 & ~i234;
assign a3918 = ~a3914 & i234;
assign a3920 = ~a3918 & ~a3916;
assign a3922 = a3920 & a3908;
assign a3924 = a3446 & ~l500;
assign a3926 = ~a3446 & ~l688;
assign a3928 = ~a3926 & ~a3924;
assign a3930 = a3928 & ~i236;
assign a3932 = ~a3928 & i236;
assign a3934 = ~a3932 & ~a3930;
assign a3936 = a3934 & a3922;
assign a3938 = a3446 & ~l502;
assign a3940 = ~a3446 & ~l690;
assign a3942 = ~a3940 & ~a3938;
assign a3944 = a3942 & ~i238;
assign a3946 = ~a3942 & i238;
assign a3948 = ~a3946 & ~a3944;
assign a3950 = a3948 & a3936;
assign a3952 = a3446 & ~l504;
assign a3954 = ~a3446 & ~l692;
assign a3956 = ~a3954 & ~a3952;
assign a3958 = a3956 & ~i240;
assign a3960 = ~a3956 & i240;
assign a3962 = ~a3960 & ~a3958;
assign a3964 = a3962 & a3950;
assign a3966 = a3446 & ~l506;
assign a3968 = ~a3446 & ~l694;
assign a3970 = ~a3968 & ~a3966;
assign a3972 = a3970 & ~i242;
assign a3974 = ~a3970 & i242;
assign a3976 = ~a3974 & ~a3972;
assign a3978 = a3976 & a3964;
assign a3980 = a3446 & ~l512;
assign a3982 = ~a3446 & ~l696;
assign a3984 = ~a3982 & ~a3980;
assign a3986 = a3984 & ~i244;
assign a3988 = ~a3984 & i244;
assign a3990 = ~a3988 & ~a3986;
assign a3992 = a3990 & a3978;
assign a3994 = ~a3446 & ~l698;
assign a3996 = a3446 & l514;
assign a3998 = ~a3996 & ~a3994;
assign a4000 = a3998 & ~i246;
assign a4002 = ~a3998 & i246;
assign a4004 = ~a4002 & ~a4000;
assign a4006 = a4004 & a3992;
assign a4008 = a3446 & ~l518;
assign a4010 = ~a3446 & ~l700;
assign a4012 = ~a4010 & ~a4008;
assign a4014 = a4012 & ~i248;
assign a4016 = ~a4012 & i248;
assign a4018 = ~a4016 & ~a4014;
assign a4020 = a4018 & a4006;
assign a4022 = ~a3446 & ~l702;
assign a4024 = a3446 & l520;
assign a4026 = ~a4024 & ~a4022;
assign a4028 = a4026 & ~i250;
assign a4030 = ~a4026 & i250;
assign a4032 = ~a4030 & ~a4028;
assign a4034 = a4032 & a4020;
assign a4036 = a3446 & ~l526;
assign a4038 = ~a3446 & ~l704;
assign a4040 = ~a4038 & ~a4036;
assign a4042 = a4040 & ~i252;
assign a4044 = ~a4040 & i252;
assign a4046 = ~a4044 & ~a4042;
assign a4048 = a4046 & a4034;
assign a4050 = ~a3446 & ~l706;
assign a4052 = a3446 & l528;
assign a4054 = ~a4052 & ~a4050;
assign a4056 = a4054 & ~i254;
assign a4058 = ~a4054 & i254;
assign a4060 = ~a4058 & ~a4056;
assign a4062 = a4060 & a4048;
assign a4064 = a3446 & ~l532;
assign a4066 = ~a3446 & ~l708;
assign a4068 = ~a4066 & ~a4064;
assign a4070 = a4068 & ~i256;
assign a4072 = ~a4068 & i256;
assign a4074 = ~a4072 & ~a4070;
assign a4076 = a4074 & a4062;
assign a4078 = ~a3446 & ~l710;
assign a4080 = a3446 & l534;
assign a4082 = ~a4080 & ~a4078;
assign a4084 = a4082 & ~i258;
assign a4086 = ~a4082 & i258;
assign a4088 = ~a4086 & ~a4084;
assign a4090 = a4088 & a4076;
assign a4092 = a3446 & ~l536;
assign a4094 = ~a3446 & ~l712;
assign a4096 = ~a4094 & ~a4092;
assign a4098 = a4096 & ~i260;
assign a4100 = ~a4096 & i260;
assign a4102 = ~a4100 & ~a4098;
assign a4104 = a4102 & a4090;
assign a4106 = a3446 & ~l538;
assign a4108 = ~a3446 & ~l714;
assign a4110 = ~a4108 & ~a4106;
assign a4112 = a4110 & ~i262;
assign a4114 = ~a4110 & i262;
assign a4116 = ~a4114 & ~a4112;
assign a4118 = a4116 & a4104;
assign a4120 = ~a3446 & ~l716;
assign a4122 = a3446 & l540;
assign a4124 = ~a4122 & ~a4120;
assign a4126 = a4124 & ~i264;
assign a4128 = ~a4124 & i264;
assign a4130 = ~a4128 & ~a4126;
assign a4132 = a4130 & a4118;
assign a4134 = a3446 & ~l542;
assign a4136 = ~a3446 & ~l718;
assign a4138 = ~a4136 & ~a4134;
assign a4140 = a4138 & ~i266;
assign a4142 = ~a4138 & i266;
assign a4144 = ~a4142 & ~a4140;
assign a4146 = a4144 & a4132;
assign a4148 = a3446 & ~l544;
assign a4150 = ~a3446 & ~l720;
assign a4152 = ~a4150 & ~a4148;
assign a4154 = a4152 & ~i268;
assign a4156 = ~a4152 & i268;
assign a4158 = ~a4156 & ~a4154;
assign a4160 = a4158 & a4146;
assign a4162 = a3446 & ~l548;
assign a4164 = ~a3446 & ~l722;
assign a4166 = ~a4164 & ~a4162;
assign a4168 = a4166 & ~i270;
assign a4170 = ~a4166 & i270;
assign a4172 = ~a4170 & ~a4168;
assign a4174 = a4172 & a4160;
assign a4176 = a3446 & ~l550;
assign a4178 = ~a3446 & ~l724;
assign a4180 = ~a4178 & ~a4176;
assign a4182 = a4180 & ~i272;
assign a4184 = ~a4180 & i272;
assign a4186 = ~a4184 & ~a4182;
assign a4188 = a4186 & a4174;
assign a4190 = a3446 & ~l552;
assign a4192 = ~a3446 & ~l726;
assign a4194 = ~a4192 & ~a4190;
assign a4196 = a4194 & ~i274;
assign a4198 = ~a4194 & i274;
assign a4200 = ~a4198 & ~a4196;
assign a4202 = a4200 & a4188;
assign a4204 = a3446 & ~l554;
assign a4206 = ~a3446 & ~l728;
assign a4208 = ~a4206 & ~a4204;
assign a4210 = a4208 & ~i276;
assign a4212 = ~a4208 & i276;
assign a4214 = ~a4212 & ~a4210;
assign a4216 = a4214 & a4202;
assign a4218 = a3446 & ~l556;
assign a4220 = ~a3446 & ~l730;
assign a4222 = ~a4220 & ~a4218;
assign a4224 = a4222 & ~i278;
assign a4226 = ~a4222 & i278;
assign a4228 = ~a4226 & ~a4224;
assign a4230 = a4228 & a4216;
assign a4232 = a3446 & ~l558;
assign a4234 = ~a3446 & ~l732;
assign a4236 = ~a4234 & ~a4232;
assign a4238 = a4236 & ~i280;
assign a4240 = ~a4236 & i280;
assign a4242 = ~a4240 & ~a4238;
assign a4244 = a4242 & a4230;
assign a4246 = a3446 & ~l564;
assign a4248 = ~a3446 & ~l734;
assign a4250 = ~a4248 & ~a4246;
assign a4252 = a4250 & ~i282;
assign a4254 = ~a4250 & i282;
assign a4256 = ~a4254 & ~a4252;
assign a4258 = a4256 & a4244;
assign a4260 = ~a3446 & ~l736;
assign a4262 = a3446 & l566;
assign a4264 = ~a4262 & ~a4260;
assign a4266 = a4264 & ~i284;
assign a4268 = ~a4264 & i284;
assign a4270 = ~a4268 & ~a4266;
assign a4272 = a4270 & a4258;
assign a4274 = a3446 & ~l570;
assign a4276 = ~a3446 & ~l738;
assign a4278 = ~a4276 & ~a4274;
assign a4280 = a4278 & ~i286;
assign a4282 = ~a4278 & i286;
assign a4284 = ~a4282 & ~a4280;
assign a4286 = a4284 & a4272;
assign a4288 = ~a3446 & ~l740;
assign a4290 = a3446 & l572;
assign a4292 = ~a4290 & ~a4288;
assign a4294 = a4292 & ~i288;
assign a4296 = ~a4292 & i288;
assign a4298 = ~a4296 & ~a4294;
assign a4300 = a4298 & a4286;
assign a4302 = a3446 & ~l578;
assign a4304 = ~a3446 & ~l742;
assign a4306 = ~a4304 & ~a4302;
assign a4308 = a4306 & ~i290;
assign a4310 = ~a4306 & i290;
assign a4312 = ~a4310 & ~a4308;
assign a4314 = a4312 & a4300;
assign a4316 = ~a3446 & ~l744;
assign a4318 = a3446 & l580;
assign a4320 = ~a4318 & ~a4316;
assign a4322 = a4320 & ~i292;
assign a4324 = ~a4320 & i292;
assign a4326 = ~a4324 & ~a4322;
assign a4328 = a4326 & a4314;
assign a4330 = a3446 & ~l584;
assign a4332 = ~a3446 & ~l746;
assign a4334 = ~a4332 & ~a4330;
assign a4336 = a4334 & ~i294;
assign a4338 = ~a4334 & i294;
assign a4340 = ~a4338 & ~a4336;
assign a4342 = a4340 & a4328;
assign a4344 = ~a3446 & ~l748;
assign a4346 = a3446 & l586;
assign a4348 = ~a4346 & ~a4344;
assign a4350 = a4348 & ~i296;
assign a4352 = ~a4348 & i296;
assign a4354 = ~a4352 & ~a4350;
assign a4356 = a4354 & a4342;
assign a4358 = a3446 & ~l588;
assign a4360 = ~a3446 & ~l750;
assign a4362 = ~a4360 & ~a4358;
assign a4364 = a4362 & ~i298;
assign a4366 = ~a4362 & i298;
assign a4368 = ~a4366 & ~a4364;
assign a4370 = a4368 & a4356;
assign a4372 = a3446 & ~l590;
assign a4374 = ~a3446 & ~l752;
assign a4376 = ~a4374 & ~a4372;
assign a4378 = a4376 & ~i300;
assign a4380 = ~a4376 & i300;
assign a4382 = ~a4380 & ~a4378;
assign a4384 = a4382 & a4370;
assign a4386 = ~a3446 & ~l754;
assign a4388 = a3446 & l592;
assign a4390 = ~a4388 & ~a4386;
assign a4392 = a4390 & ~i302;
assign a4394 = ~a4390 & i302;
assign a4396 = ~a4394 & ~a4392;
assign a4398 = a4396 & a4384;
assign a4400 = a3446 & ~l594;
assign a4402 = ~a3446 & ~l756;
assign a4404 = ~a4402 & ~a4400;
assign a4406 = a4404 & ~i304;
assign a4408 = ~a4404 & i304;
assign a4410 = ~a4408 & ~a4406;
assign a4412 = a4410 & a4398;
assign a4414 = a3446 & ~l596;
assign a4416 = ~a3446 & ~l758;
assign a4418 = ~a4416 & ~a4414;
assign a4420 = a4418 & ~i306;
assign a4422 = ~a4418 & i306;
assign a4424 = ~a4422 & ~a4420;
assign a4426 = a4424 & a4412;
assign a4428 = a3446 & ~l600;
assign a4430 = ~a3446 & ~l760;
assign a4432 = ~a4430 & ~a4428;
assign a4434 = a4432 & ~i308;
assign a4436 = ~a4432 & i308;
assign a4438 = ~a4436 & ~a4434;
assign a4440 = a4438 & a4426;
assign a4442 = a3446 & ~l602;
assign a4444 = ~a3446 & ~l762;
assign a4446 = ~a4444 & ~a4442;
assign a4448 = a4446 & ~i310;
assign a4450 = ~a4446 & i310;
assign a4452 = ~a4450 & ~a4448;
assign a4454 = a4452 & a4440;
assign a4456 = a3446 & ~l604;
assign a4458 = ~a3446 & ~l764;
assign a4460 = ~a4458 & ~a4456;
assign a4462 = a4460 & ~i312;
assign a4464 = ~a4460 & i312;
assign a4466 = ~a4464 & ~a4462;
assign a4468 = a4466 & a4454;
assign a4470 = a3446 & ~l606;
assign a4472 = ~a3446 & ~l766;
assign a4474 = ~a4472 & ~a4470;
assign a4476 = a4474 & ~i314;
assign a4478 = ~a4474 & i314;
assign a4480 = ~a4478 & ~a4476;
assign a4482 = a4480 & a4468;
assign a4484 = a3446 & ~l608;
assign a4486 = ~a3446 & ~l768;
assign a4488 = ~a4486 & ~a4484;
assign a4490 = a4488 & ~i316;
assign a4492 = ~a4488 & i316;
assign a4494 = ~a4492 & ~a4490;
assign a4496 = a4494 & a4482;
assign a4498 = a3446 & ~l610;
assign a4500 = ~a3446 & ~l770;
assign a4502 = ~a4500 & ~a4498;
assign a4504 = a4502 & ~i318;
assign a4506 = ~a4502 & i318;
assign a4508 = ~a4506 & ~a4504;
assign a4510 = a4508 & a4496;
assign a4512 = a3446 & ~l612;
assign a4514 = ~a3446 & ~l772;
assign a4516 = ~a4514 & ~a4512;
assign a4518 = a4516 & ~i320;
assign a4520 = ~a4516 & i320;
assign a4522 = ~a4520 & ~a4518;
assign a4524 = a4522 & a4510;
assign a4526 = a3446 & ~l614;
assign a4528 = ~a3446 & ~l774;
assign a4530 = ~a4528 & ~a4526;
assign a4532 = a4530 & ~i322;
assign a4534 = ~a4530 & i322;
assign a4536 = ~a4534 & ~a4532;
assign a4538 = a4536 & a4524;
assign a4540 = a3446 & ~l616;
assign a4542 = ~a3446 & ~l776;
assign a4544 = ~a4542 & ~a4540;
assign a4546 = a4544 & ~i324;
assign a4548 = ~a4544 & i324;
assign a4550 = ~a4548 & ~a4546;
assign a4552 = a4550 & a4538;
assign a4554 = a3446 & ~l618;
assign a4556 = ~a3446 & ~l778;
assign a4558 = ~a4556 & ~a4554;
assign a4560 = a4558 & ~i326;
assign a4562 = ~a4558 & i326;
assign a4564 = ~a4562 & ~a4560;
assign a4566 = a4564 & a4552;
assign a4568 = ~l344 & ~l342;
assign a4570 = ~a4568 & l340;
assign a4572 = ~l352 & ~l350;
assign a4574 = ~a4572 & l348;
assign a4576 = ~l360 & ~l358;
assign a4578 = ~a4576 & l356;
assign a4580 = ~l368 & ~l366;
assign a4582 = ~a4580 & l364;
assign a4584 = ~l376 & ~l374;
assign a4586 = ~a4584 & l372;
assign a4588 = ~l384 & ~l382;
assign a4590 = ~a4588 & l380;
assign a4592 = ~l392 & ~l390;
assign a4594 = ~a4592 & l388;
assign a4596 = ~l400 & ~l398;
assign a4598 = ~a4596 & l396;
assign a4600 = l406 & l404;
assign a4602 = ~l410 & l408;
assign a4604 = l420 & l418;
assign a4606 = ~l424 & l422;
assign a4608 = a886 & l432;
assign a4610 = a1130 & l448;
assign a4612 = l458 & l456;
assign a4614 = ~l462 & l460;
assign a4616 = l472 & l470;
assign a4618 = ~l476 & l474;
assign a4620 = a1370 & l484;
assign a4622 = a1614 & l500;
assign a4624 = l510 & l508;
assign a4626 = ~l514 & l512;
assign a4628 = l524 & l522;
assign a4630 = ~l528 & l526;
assign a4632 = a1854 & l536;
assign a4634 = a2098 & l552;
assign a4636 = l562 & l560;
assign a4638 = ~l566 & l564;
assign a4640 = l576 & l574;
assign a4642 = ~l580 & l578;
assign a4644 = a2338 & l588;
assign a4646 = a2582 & l604;
assign a4648 = l622 & l620;
assign a4650 = l630 & l628;
assign a4652 = l640 & l638;
assign a4654 = a4652 & l636;
assign a4656 = l654 & l652;
assign a4658 = a4656 & l650;
assign a4660 = l660 & l658;
assign a4662 = l668 & l666;
assign a4664 = l678 & l676;
assign a4666 = a4664 & l674;
assign a4668 = l692 & l690;
assign a4670 = a4668 & l688;
assign a4672 = l698 & l696;
assign a4674 = l706 & l704;
assign a4676 = l716 & l714;
assign a4678 = a4676 & l712;
assign a4680 = l730 & l728;
assign a4682 = a4680 & l726;
assign a4684 = l736 & l734;
assign a4686 = l744 & l742;
assign a4688 = l754 & l752;
assign a4690 = a4688 & l750;
assign a4692 = l768 & l766;
assign a4694 = a4692 & l764;
assign a4696 = ~l548 & ~l496;
assign a4698 = l548 & l496;
assign a4700 = ~a4698 & ~a4696;
assign a4702 = a1784 & a1300;
assign a4704 = a4702 & ~a4700;
assign a4706 = ~l496 & ~l444;
assign a4708 = l496 & l444;
assign a4710 = ~a4708 & ~a4706;
assign a4712 = ~a4710 & a1300;
assign a4714 = ~l548 & ~l444;
assign a4716 = l548 & l444;
assign a4718 = ~a4716 & ~a4714;
assign a4720 = ~a4718 & a1784;
assign a4722 = ~l600 & ~l444;
assign a4724 = l600 & l444;
assign a4726 = ~a4724 & ~a4722;
assign a4728 = ~a4726 & a2268;
assign a4730 = ~a4728 & ~a4720;
assign a4732 = a4730 & ~a4712;
assign a4734 = ~a4732 & a816;
assign a4736 = ~l600 & ~l496;
assign a4738 = l600 & l496;
assign a4740 = ~a4738 & ~a4736;
assign a4742 = a2268 & a1300;
assign a4744 = a4742 & ~a4740;
assign a4746 = ~l600 & ~l548;
assign a4748 = l600 & l548;
assign a4750 = ~a4748 & ~a4746;
assign a4752 = a2268 & a1784;
assign a4754 = a4752 & ~a4750;
assign a4756 = ~a4754 & ~a4744;
assign a4758 = a4756 & ~a4734;
assign a4760 = a4758 & ~a4704;
assign a4762 = ~a4760 & l612;
assign a4764 = a4568 & ~l340;
assign a4766 = l344 & ~l342;
assign a4768 = a4766 & ~l340;
assign a4770 = ~l344 & l342;
assign a4772 = a4770 & ~l340;
assign a4774 = l344 & l342;
assign a4776 = a4774 & ~l340;
assign a4778 = ~l564 & ~l346;
assign a4780 = ~l578 & l346;
assign a4782 = ~a4780 & ~a4778;
assign a4784 = a4568 & l340;
assign a4786 = a4784 & ~a4782;
assign a4788 = a4786 & ~a4776;
assign a4790 = ~l512 & ~l346;
assign a4792 = ~l526 & l346;
assign a4794 = ~a4792 & ~a4790;
assign a4796 = ~a4794 & a4776;
assign a4798 = ~a4796 & ~a4788;
assign a4800 = ~a4798 & ~a4772;
assign a4802 = ~l460 & ~l346;
assign a4804 = ~l474 & l346;
assign a4806 = ~a4804 & ~a4802;
assign a4808 = ~a4806 & a4772;
assign a4810 = ~a4808 & ~a4800;
assign a4812 = ~a4810 & ~a4768;
assign a4814 = ~l408 & ~l346;
assign a4816 = ~l422 & l346;
assign a4818 = ~a4816 & ~a4814;
assign a4820 = ~a4818 & a4768;
assign a4822 = ~a4820 & ~a4812;
assign a4824 = a4822 & ~l404;
assign a4826 = ~a4822 & l404;
assign a4828 = ~a4826 & ~a4824;
assign a4830 = l566 & ~l346;
assign a4832 = l580 & l346;
assign a4834 = ~a4832 & ~a4830;
assign a4836 = ~a4834 & a4784;
assign a4838 = a4836 & ~a4776;
assign a4840 = l514 & ~l346;
assign a4842 = l528 & l346;
assign a4844 = ~a4842 & ~a4840;
assign a4846 = ~a4844 & a4776;
assign a4848 = ~a4846 & ~a4838;
assign a4850 = ~a4848 & ~a4772;
assign a4852 = l462 & ~l346;
assign a4854 = l476 & l346;
assign a4856 = ~a4854 & ~a4852;
assign a4858 = ~a4856 & a4772;
assign a4860 = ~a4858 & ~a4850;
assign a4862 = ~a4860 & ~a4768;
assign a4864 = l410 & ~l346;
assign a4866 = l424 & l346;
assign a4868 = ~a4866 & ~a4864;
assign a4870 = ~a4868 & a4768;
assign a4872 = ~a4870 & ~a4862;
assign a4874 = a4872 & ~l406;
assign a4876 = ~a4872 & l406;
assign a4878 = ~a4876 & ~a4874;
assign a4880 = a4878 & a4828;
assign a4882 = ~a4880 & ~a4764;
assign a4884 = a4572 & ~l348;
assign a4886 = l352 & ~l350;
assign a4888 = a4886 & ~l348;
assign a4890 = ~l352 & l350;
assign a4892 = a4890 & ~l348;
assign a4894 = l352 & l350;
assign a4896 = a4894 & ~l348;
assign a4898 = ~l564 & ~l354;
assign a4900 = ~l578 & l354;
assign a4902 = ~a4900 & ~a4898;
assign a4904 = a4572 & l348;
assign a4906 = a4904 & ~a4902;
assign a4908 = a4906 & ~a4896;
assign a4910 = ~l512 & ~l354;
assign a4912 = ~l526 & l354;
assign a4914 = ~a4912 & ~a4910;
assign a4916 = ~a4914 & a4896;
assign a4918 = ~a4916 & ~a4908;
assign a4920 = ~a4918 & ~a4892;
assign a4922 = ~l460 & ~l354;
assign a4924 = ~l474 & l354;
assign a4926 = ~a4924 & ~a4922;
assign a4928 = ~a4926 & a4892;
assign a4930 = ~a4928 & ~a4920;
assign a4932 = ~a4930 & ~a4888;
assign a4934 = ~l408 & ~l354;
assign a4936 = ~l422 & l354;
assign a4938 = ~a4936 & ~a4934;
assign a4940 = ~a4938 & a4888;
assign a4942 = ~a4940 & ~a4932;
assign a4944 = a4942 & ~l418;
assign a4946 = ~a4942 & l418;
assign a4948 = ~a4946 & ~a4944;
assign a4950 = l566 & ~l354;
assign a4952 = l580 & l354;
assign a4954 = ~a4952 & ~a4950;
assign a4956 = ~a4954 & a4904;
assign a4958 = a4956 & ~a4896;
assign a4960 = l514 & ~l354;
assign a4962 = l528 & l354;
assign a4964 = ~a4962 & ~a4960;
assign a4966 = ~a4964 & a4896;
assign a4968 = ~a4966 & ~a4958;
assign a4970 = ~a4968 & ~a4892;
assign a4972 = l462 & ~l354;
assign a4974 = l476 & l354;
assign a4976 = ~a4974 & ~a4972;
assign a4978 = ~a4976 & a4892;
assign a4980 = ~a4978 & ~a4970;
assign a4982 = ~a4980 & ~a4888;
assign a4984 = l410 & ~l354;
assign a4986 = l424 & l354;
assign a4988 = ~a4986 & ~a4984;
assign a4990 = ~a4988 & a4888;
assign a4992 = ~a4990 & ~a4982;
assign a4994 = a4992 & ~l420;
assign a4996 = ~a4992 & l420;
assign a4998 = ~a4996 & ~a4994;
assign a5000 = a4998 & a4948;
assign a5002 = ~a5000 & ~a4884;
assign a5004 = a4576 & ~l356;
assign a5006 = l360 & ~l358;
assign a5008 = a5006 & ~l356;
assign a5010 = ~l360 & l358;
assign a5012 = a5010 & ~l356;
assign a5014 = l360 & l358;
assign a5016 = a5014 & ~l356;
assign a5018 = ~l564 & ~l362;
assign a5020 = ~l578 & l362;
assign a5022 = ~a5020 & ~a5018;
assign a5024 = a4576 & l356;
assign a5026 = a5024 & ~a5022;
assign a5028 = a5026 & ~a5016;
assign a5030 = ~l512 & ~l362;
assign a5032 = ~l526 & l362;
assign a5034 = ~a5032 & ~a5030;
assign a5036 = ~a5034 & a5016;
assign a5038 = ~a5036 & ~a5028;
assign a5040 = ~a5038 & ~a5012;
assign a5042 = ~l460 & ~l362;
assign a5044 = ~l474 & l362;
assign a5046 = ~a5044 & ~a5042;
assign a5048 = ~a5046 & a5012;
assign a5050 = ~a5048 & ~a5040;
assign a5052 = ~a5050 & ~a5008;
assign a5054 = ~l408 & ~l362;
assign a5056 = ~l422 & l362;
assign a5058 = ~a5056 & ~a5054;
assign a5060 = ~a5058 & a5008;
assign a5062 = ~a5060 & ~a5052;
assign a5064 = a5062 & ~l456;
assign a5066 = ~a5062 & l456;
assign a5068 = ~a5066 & ~a5064;
assign a5070 = l566 & ~l362;
assign a5072 = l580 & l362;
assign a5074 = ~a5072 & ~a5070;
assign a5076 = ~a5074 & a5024;
assign a5078 = a5076 & ~a5016;
assign a5080 = l514 & ~l362;
assign a5082 = l528 & l362;
assign a5084 = ~a5082 & ~a5080;
assign a5086 = ~a5084 & a5016;
assign a5088 = ~a5086 & ~a5078;
assign a5090 = ~a5088 & ~a5012;
assign a5092 = l462 & ~l362;
assign a5094 = l476 & l362;
assign a5096 = ~a5094 & ~a5092;
assign a5098 = ~a5096 & a5012;
assign a5100 = ~a5098 & ~a5090;
assign a5102 = ~a5100 & ~a5008;
assign a5104 = l410 & ~l362;
assign a5106 = l424 & l362;
assign a5108 = ~a5106 & ~a5104;
assign a5110 = ~a5108 & a5008;
assign a5112 = ~a5110 & ~a5102;
assign a5114 = a5112 & ~l458;
assign a5116 = ~a5112 & l458;
assign a5118 = ~a5116 & ~a5114;
assign a5120 = a5118 & a5068;
assign a5122 = ~a5120 & ~a5004;
assign a5124 = a4580 & ~l364;
assign a5126 = l368 & ~l366;
assign a5128 = a5126 & ~l364;
assign a5130 = ~l368 & l366;
assign a5132 = a5130 & ~l364;
assign a5134 = l368 & l366;
assign a5136 = a5134 & ~l364;
assign a5138 = ~l564 & ~l370;
assign a5140 = ~l578 & l370;
assign a5142 = ~a5140 & ~a5138;
assign a5144 = a4580 & l364;
assign a5146 = a5144 & ~a5142;
assign a5148 = a5146 & ~a5136;
assign a5150 = ~l512 & ~l370;
assign a5152 = ~l526 & l370;
assign a5154 = ~a5152 & ~a5150;
assign a5156 = ~a5154 & a5136;
assign a5158 = ~a5156 & ~a5148;
assign a5160 = ~a5158 & ~a5132;
assign a5162 = ~l460 & ~l370;
assign a5164 = ~l474 & l370;
assign a5166 = ~a5164 & ~a5162;
assign a5168 = ~a5166 & a5132;
assign a5170 = ~a5168 & ~a5160;
assign a5172 = ~a5170 & ~a5128;
assign a5174 = ~l408 & ~l370;
assign a5176 = ~l422 & l370;
assign a5178 = ~a5176 & ~a5174;
assign a5180 = ~a5178 & a5128;
assign a5182 = ~a5180 & ~a5172;
assign a5184 = a5182 & ~l470;
assign a5186 = ~a5182 & l470;
assign a5188 = ~a5186 & ~a5184;
assign a5190 = l566 & ~l370;
assign a5192 = l580 & l370;
assign a5194 = ~a5192 & ~a5190;
assign a5196 = ~a5194 & a5144;
assign a5198 = a5196 & ~a5136;
assign a5200 = l514 & ~l370;
assign a5202 = l528 & l370;
assign a5204 = ~a5202 & ~a5200;
assign a5206 = ~a5204 & a5136;
assign a5208 = ~a5206 & ~a5198;
assign a5210 = ~a5208 & ~a5132;
assign a5212 = l462 & ~l370;
assign a5214 = l476 & l370;
assign a5216 = ~a5214 & ~a5212;
assign a5218 = ~a5216 & a5132;
assign a5220 = ~a5218 & ~a5210;
assign a5222 = ~a5220 & ~a5128;
assign a5224 = l410 & ~l370;
assign a5226 = l424 & l370;
assign a5228 = ~a5226 & ~a5224;
assign a5230 = ~a5228 & a5128;
assign a5232 = ~a5230 & ~a5222;
assign a5234 = a5232 & ~l472;
assign a5236 = ~a5232 & l472;
assign a5238 = ~a5236 & ~a5234;
assign a5240 = a5238 & a5188;
assign a5242 = ~a5240 & ~a5124;
assign a5244 = a4584 & ~l372;
assign a5246 = l376 & ~l374;
assign a5248 = a5246 & ~l372;
assign a5250 = ~l376 & l374;
assign a5252 = a5250 & ~l372;
assign a5254 = l376 & l374;
assign a5256 = a5254 & ~l372;
assign a5258 = ~l564 & ~l378;
assign a5260 = ~l578 & l378;
assign a5262 = ~a5260 & ~a5258;
assign a5264 = a4584 & l372;
assign a5266 = a5264 & ~a5262;
assign a5268 = a5266 & ~a5256;
assign a5270 = ~l512 & ~l378;
assign a5272 = ~l526 & l378;
assign a5274 = ~a5272 & ~a5270;
assign a5276 = ~a5274 & a5256;
assign a5278 = ~a5276 & ~a5268;
assign a5280 = ~a5278 & ~a5252;
assign a5282 = ~l460 & ~l378;
assign a5284 = ~l474 & l378;
assign a5286 = ~a5284 & ~a5282;
assign a5288 = ~a5286 & a5252;
assign a5290 = ~a5288 & ~a5280;
assign a5292 = ~a5290 & ~a5248;
assign a5294 = ~l408 & ~l378;
assign a5296 = ~l422 & l378;
assign a5298 = ~a5296 & ~a5294;
assign a5300 = ~a5298 & a5248;
assign a5302 = ~a5300 & ~a5292;
assign a5304 = a5302 & ~l508;
assign a5306 = ~a5302 & l508;
assign a5308 = ~a5306 & ~a5304;
assign a5310 = l566 & ~l378;
assign a5312 = l580 & l378;
assign a5314 = ~a5312 & ~a5310;
assign a5316 = ~a5314 & a5264;
assign a5318 = a5316 & ~a5256;
assign a5320 = l514 & ~l378;
assign a5322 = l528 & l378;
assign a5324 = ~a5322 & ~a5320;
assign a5326 = ~a5324 & a5256;
assign a5328 = ~a5326 & ~a5318;
assign a5330 = ~a5328 & ~a5252;
assign a5332 = l462 & ~l378;
assign a5334 = l476 & l378;
assign a5336 = ~a5334 & ~a5332;
assign a5338 = ~a5336 & a5252;
assign a5340 = ~a5338 & ~a5330;
assign a5342 = ~a5340 & ~a5248;
assign a5344 = l410 & ~l378;
assign a5346 = l424 & l378;
assign a5348 = ~a5346 & ~a5344;
assign a5350 = ~a5348 & a5248;
assign a5352 = ~a5350 & ~a5342;
assign a5354 = a5352 & ~l510;
assign a5356 = ~a5352 & l510;
assign a5358 = ~a5356 & ~a5354;
assign a5360 = a5358 & a5308;
assign a5362 = ~a5360 & ~a5244;
assign a5364 = a4588 & ~l380;
assign a5366 = l384 & ~l382;
assign a5368 = a5366 & ~l380;
assign a5370 = ~l384 & l382;
assign a5372 = a5370 & ~l380;
assign a5374 = l384 & l382;
assign a5376 = a5374 & ~l380;
assign a5378 = ~l564 & ~l386;
assign a5380 = ~l578 & l386;
assign a5382 = ~a5380 & ~a5378;
assign a5384 = a4588 & l380;
assign a5386 = a5384 & ~a5382;
assign a5388 = a5386 & ~a5376;
assign a5390 = ~l512 & ~l386;
assign a5392 = ~l526 & l386;
assign a5394 = ~a5392 & ~a5390;
assign a5396 = ~a5394 & a5376;
assign a5398 = ~a5396 & ~a5388;
assign a5400 = ~a5398 & ~a5372;
assign a5402 = ~l460 & ~l386;
assign a5404 = ~l474 & l386;
assign a5406 = ~a5404 & ~a5402;
assign a5408 = ~a5406 & a5372;
assign a5410 = ~a5408 & ~a5400;
assign a5412 = ~a5410 & ~a5368;
assign a5414 = ~l408 & ~l386;
assign a5416 = ~l422 & l386;
assign a5418 = ~a5416 & ~a5414;
assign a5420 = ~a5418 & a5368;
assign a5422 = ~a5420 & ~a5412;
assign a5424 = a5422 & ~l522;
assign a5426 = ~a5422 & l522;
assign a5428 = ~a5426 & ~a5424;
assign a5430 = l566 & ~l386;
assign a5432 = l580 & l386;
assign a5434 = ~a5432 & ~a5430;
assign a5436 = ~a5434 & a5384;
assign a5438 = a5436 & ~a5376;
assign a5440 = l514 & ~l386;
assign a5442 = l528 & l386;
assign a5444 = ~a5442 & ~a5440;
assign a5446 = ~a5444 & a5376;
assign a5448 = ~a5446 & ~a5438;
assign a5450 = ~a5448 & ~a5372;
assign a5452 = l462 & ~l386;
assign a5454 = l476 & l386;
assign a5456 = ~a5454 & ~a5452;
assign a5458 = ~a5456 & a5372;
assign a5460 = ~a5458 & ~a5450;
assign a5462 = ~a5460 & ~a5368;
assign a5464 = l410 & ~l386;
assign a5466 = l424 & l386;
assign a5468 = ~a5466 & ~a5464;
assign a5470 = ~a5468 & a5368;
assign a5472 = ~a5470 & ~a5462;
assign a5474 = a5472 & ~l524;
assign a5476 = ~a5472 & l524;
assign a5478 = ~a5476 & ~a5474;
assign a5480 = a5478 & a5428;
assign a5482 = ~a5480 & ~a5364;
assign a5484 = a4592 & ~l388;
assign a5486 = l392 & ~l390;
assign a5488 = a5486 & ~l388;
assign a5490 = ~l392 & l390;
assign a5492 = a5490 & ~l388;
assign a5494 = l392 & l390;
assign a5496 = a5494 & ~l388;
assign a5498 = ~l564 & ~l394;
assign a5500 = ~l578 & l394;
assign a5502 = ~a5500 & ~a5498;
assign a5504 = a4592 & l388;
assign a5506 = a5504 & ~a5502;
assign a5508 = a5506 & ~a5496;
assign a5510 = ~l512 & ~l394;
assign a5512 = ~l526 & l394;
assign a5514 = ~a5512 & ~a5510;
assign a5516 = ~a5514 & a5496;
assign a5518 = ~a5516 & ~a5508;
assign a5520 = ~a5518 & ~a5492;
assign a5522 = ~l460 & ~l394;
assign a5524 = ~l474 & l394;
assign a5526 = ~a5524 & ~a5522;
assign a5528 = ~a5526 & a5492;
assign a5530 = ~a5528 & ~a5520;
assign a5532 = ~a5530 & ~a5488;
assign a5534 = ~l408 & ~l394;
assign a5536 = ~l422 & l394;
assign a5538 = ~a5536 & ~a5534;
assign a5540 = ~a5538 & a5488;
assign a5542 = ~a5540 & ~a5532;
assign a5544 = a5542 & ~l560;
assign a5546 = ~a5542 & l560;
assign a5548 = ~a5546 & ~a5544;
assign a5550 = l566 & ~l394;
assign a5552 = l580 & l394;
assign a5554 = ~a5552 & ~a5550;
assign a5556 = ~a5554 & a5504;
assign a5558 = a5556 & ~a5496;
assign a5560 = l514 & ~l394;
assign a5562 = l528 & l394;
assign a5564 = ~a5562 & ~a5560;
assign a5566 = ~a5564 & a5496;
assign a5568 = ~a5566 & ~a5558;
assign a5570 = ~a5568 & ~a5492;
assign a5572 = l462 & ~l394;
assign a5574 = l476 & l394;
assign a5576 = ~a5574 & ~a5572;
assign a5578 = ~a5576 & a5492;
assign a5580 = ~a5578 & ~a5570;
assign a5582 = ~a5580 & ~a5488;
assign a5584 = l410 & ~l394;
assign a5586 = l424 & l394;
assign a5588 = ~a5586 & ~a5584;
assign a5590 = ~a5588 & a5488;
assign a5592 = ~a5590 & ~a5582;
assign a5594 = a5592 & ~l562;
assign a5596 = ~a5592 & l562;
assign a5598 = ~a5596 & ~a5594;
assign a5600 = a5598 & a5548;
assign a5602 = ~a5600 & ~a5484;
assign a5604 = a4596 & ~l396;
assign a5606 = l400 & ~l398;
assign a5608 = a5606 & ~l396;
assign a5610 = ~l400 & l398;
assign a5612 = a5610 & ~l396;
assign a5614 = l400 & l398;
assign a5616 = a5614 & ~l396;
assign a5618 = ~l564 & ~l402;
assign a5620 = ~l578 & l402;
assign a5622 = ~a5620 & ~a5618;
assign a5624 = a4596 & l396;
assign a5626 = a5624 & ~a5622;
assign a5628 = a5626 & ~a5616;
assign a5630 = ~l512 & ~l402;
assign a5632 = ~l526 & l402;
assign a5634 = ~a5632 & ~a5630;
assign a5636 = ~a5634 & a5616;
assign a5638 = ~a5636 & ~a5628;
assign a5640 = ~a5638 & ~a5612;
assign a5642 = ~l460 & ~l402;
assign a5644 = ~l474 & l402;
assign a5646 = ~a5644 & ~a5642;
assign a5648 = ~a5646 & a5612;
assign a5650 = ~a5648 & ~a5640;
assign a5652 = ~a5650 & ~a5608;
assign a5654 = ~l408 & ~l402;
assign a5656 = ~l422 & l402;
assign a5658 = ~a5656 & ~a5654;
assign a5660 = ~a5658 & a5608;
assign a5662 = ~a5660 & ~a5652;
assign a5664 = a5662 & ~l574;
assign a5666 = ~a5662 & l574;
assign a5668 = ~a5666 & ~a5664;
assign a5670 = l566 & ~l402;
assign a5672 = l580 & l402;
assign a5674 = ~a5672 & ~a5670;
assign a5676 = ~a5674 & a5624;
assign a5678 = a5676 & ~a5616;
assign a5680 = l514 & ~l402;
assign a5682 = l528 & l402;
assign a5684 = ~a5682 & ~a5680;
assign a5686 = ~a5684 & a5616;
assign a5688 = ~a5686 & ~a5678;
assign a5690 = ~a5688 & ~a5612;
assign a5692 = l462 & ~l402;
assign a5694 = l476 & l402;
assign a5696 = ~a5694 & ~a5692;
assign a5698 = ~a5696 & a5612;
assign a5700 = ~a5698 & ~a5690;
assign a5702 = ~a5700 & ~a5608;
assign a5704 = l410 & ~l402;
assign a5706 = l424 & l402;
assign a5708 = ~a5706 & ~a5704;
assign a5710 = ~a5708 & a5608;
assign a5712 = ~a5710 & ~a5702;
assign a5714 = a5712 & ~l576;
assign a5716 = ~a5712 & l576;
assign a5718 = ~a5716 & ~a5714;
assign a5720 = a5718 & a5668;
assign a5722 = ~a5720 & ~a5604;
assign a5724 = a5488 & ~l394;
assign a5726 = ~a5724 & ~l346;
assign a5728 = a5608 & ~l402;
assign a5730 = ~a5728 & l346;
assign a5732 = ~a5730 & ~a5726;
assign a5734 = ~a5732 & a4784;
assign a5736 = a5734 & ~a4776;
assign a5738 = a5248 & ~l378;
assign a5740 = ~a5738 & ~l346;
assign a5742 = a5368 & ~l386;
assign a5744 = ~a5742 & l346;
assign a5746 = ~a5744 & ~a5740;
assign a5748 = ~a5746 & a4776;
assign a5750 = ~a5748 & ~a5736;
assign a5752 = ~a5750 & ~a4772;
assign a5754 = a5008 & ~l362;
assign a5756 = ~a5754 & ~l346;
assign a5758 = a5128 & ~l370;
assign a5760 = ~a5758 & l346;
assign a5762 = ~a5760 & ~a5756;
assign a5764 = ~a5762 & a4772;
assign a5766 = ~a5764 & ~a5752;
assign a5768 = ~a5766 & ~a4768;
assign a5770 = ~a4768 & ~l346;
assign a5772 = a4888 & ~l354;
assign a5774 = ~a5772 & l346;
assign a5776 = ~a5774 & ~a5770;
assign a5778 = ~a5776 & a4768;
assign a5780 = ~a5778 & ~a5768;
assign a5782 = a5488 & l394;
assign a5784 = ~a5782 & ~l354;
assign a5786 = a5608 & l402;
assign a5788 = ~a5786 & l354;
assign a5790 = ~a5788 & ~a5784;
assign a5792 = ~a5790 & a4904;
assign a5794 = a5792 & ~a4896;
assign a5796 = a5248 & l378;
assign a5798 = ~a5796 & ~l354;
assign a5800 = a5368 & l386;
assign a5802 = ~a5800 & l354;
assign a5804 = ~a5802 & ~a5798;
assign a5806 = ~a5804 & a4896;
assign a5808 = ~a5806 & ~a5794;
assign a5810 = ~a5808 & ~a4892;
assign a5812 = a5008 & l362;
assign a5814 = ~a5812 & ~l354;
assign a5816 = a5128 & l370;
assign a5818 = ~a5816 & l354;
assign a5820 = ~a5818 & ~a5814;
assign a5822 = ~a5820 & a4892;
assign a5824 = ~a5822 & ~a5810;
assign a5826 = ~a5824 & ~a4888;
assign a5828 = a4768 & l346;
assign a5830 = ~a5828 & ~l354;
assign a5832 = ~a4888 & l354;
assign a5834 = ~a5832 & ~a5830;
assign a5836 = ~a5834 & a4888;
assign a5838 = ~a5836 & ~a5826;
assign a5840 = a5492 & ~l394;
assign a5842 = ~a5840 & ~l362;
assign a5844 = a5612 & ~l402;
assign a5846 = ~a5844 & l362;
assign a5848 = ~a5846 & ~a5842;
assign a5850 = ~a5848 & a5024;
assign a5852 = a5850 & ~a5016;
assign a5854 = a5252 & ~l378;
assign a5856 = ~a5854 & ~l362;
assign a5858 = a5372 & ~l386;
assign a5860 = ~a5858 & l362;
assign a5862 = ~a5860 & ~a5856;
assign a5864 = ~a5862 & a5016;
assign a5866 = ~a5864 & ~a5852;
assign a5868 = ~a5866 & ~a5012;
assign a5870 = ~a5012 & ~l362;
assign a5872 = a5132 & ~l370;
assign a5874 = ~a5872 & l362;
assign a5876 = ~a5874 & ~a5870;
assign a5878 = ~a5876 & a5012;
assign a5880 = ~a5878 & ~a5868;
assign a5882 = ~a5880 & ~a5008;
assign a5884 = a4772 & ~l346;
assign a5886 = ~a5884 & ~l362;
assign a5888 = a4892 & ~l354;
assign a5890 = ~a5888 & l362;
assign a5892 = ~a5890 & ~a5886;
assign a5894 = ~a5892 & a5008;
assign a5896 = ~a5894 & ~a5882;
assign a5898 = a5492 & l394;
assign a5900 = ~a5898 & ~l370;
assign a5902 = a5612 & l402;
assign a5904 = ~a5902 & l370;
assign a5906 = ~a5904 & ~a5900;
assign a5908 = ~a5906 & a5144;
assign a5910 = a5908 & ~a5136;
assign a5912 = a5252 & l378;
assign a5914 = ~a5912 & ~l370;
assign a5916 = a5372 & l386;
assign a5918 = ~a5916 & l370;
assign a5920 = ~a5918 & ~a5914;
assign a5922 = ~a5920 & a5136;
assign a5924 = ~a5922 & ~a5910;
assign a5926 = ~a5924 & ~a5132;
assign a5928 = a5012 & l362;
assign a5930 = ~a5928 & ~l370;
assign a5932 = ~a5132 & l370;
assign a5934 = ~a5932 & ~a5930;
assign a5936 = ~a5934 & a5132;
assign a5938 = ~a5936 & ~a5926;
assign a5940 = ~a5938 & ~a5128;
assign a5942 = a4772 & l346;
assign a5944 = ~a5942 & ~l370;
assign a5946 = a4892 & l354;
assign a5948 = ~a5946 & l370;
assign a5950 = ~a5948 & ~a5944;
assign a5952 = ~a5950 & a5128;
assign a5954 = ~a5952 & ~a5940;
assign a5956 = a5496 & ~l394;
assign a5958 = ~a5956 & ~l378;
assign a5960 = a5616 & ~l402;
assign a5962 = ~a5960 & l378;
assign a5964 = ~a5962 & ~a5958;
assign a5966 = ~a5964 & a5264;
assign a5968 = a5966 & ~a5256;
assign a5970 = ~a5256 & ~l378;
assign a5972 = a5376 & ~l386;
assign a5974 = ~a5972 & l378;
assign a5976 = ~a5974 & ~a5970;
assign a5978 = ~a5976 & a5256;
assign a5980 = ~a5978 & ~a5968;
assign a5982 = ~a5980 & ~a5252;
assign a5984 = a5016 & ~l362;
assign a5986 = ~a5984 & ~l378;
assign a5988 = a5136 & ~l370;
assign a5990 = ~a5988 & l378;
assign a5992 = ~a5990 & ~a5986;
assign a5994 = ~a5992 & a5252;
assign a5996 = ~a5994 & ~a5982;
assign a5998 = ~a5996 & ~a5248;
assign a6000 = a4776 & ~l346;
assign a6002 = ~a6000 & ~l378;
assign a6004 = a4896 & ~l354;
assign a6006 = ~a6004 & l378;
assign a6008 = ~a6006 & ~a6002;
assign a6010 = ~a6008 & a5248;
assign a6012 = ~a6010 & ~a5998;
assign a6014 = a5496 & l394;
assign a6016 = ~a6014 & ~l386;
assign a6018 = a5616 & l402;
assign a6020 = ~a6018 & l386;
assign a6022 = ~a6020 & ~a6016;
assign a6024 = ~a6022 & a5384;
assign a6026 = a6024 & ~a5376;
assign a6028 = a5256 & l378;
assign a6030 = ~a6028 & ~l386;
assign a6032 = ~a5376 & l386;
assign a6034 = ~a6032 & ~a6030;
assign a6036 = ~a6034 & a5376;
assign a6038 = ~a6036 & ~a6026;
assign a6040 = ~a6038 & ~a5372;
assign a6042 = a5016 & l362;
assign a6044 = ~a6042 & ~l386;
assign a6046 = a5136 & l370;
assign a6048 = ~a6046 & l386;
assign a6050 = ~a6048 & ~a6044;
assign a6052 = ~a6050 & a5372;
assign a6054 = ~a6052 & ~a6040;
assign a6056 = ~a6054 & ~a5368;
assign a6058 = a4776 & l346;
assign a6060 = ~a6058 & ~l386;
assign a6062 = a4896 & l354;
assign a6064 = ~a6062 & l386;
assign a6066 = ~a6064 & ~a6060;
assign a6068 = ~a6066 & a5368;
assign a6070 = ~a6068 & ~a6056;
assign a6072 = ~a5504 & ~l394;
assign a6074 = a5624 & ~l402;
assign a6076 = ~a6074 & l394;
assign a6078 = ~a6076 & ~a6072;
assign a6080 = ~a6078 & a5504;
assign a6082 = a6080 & ~a5496;
assign a6084 = a5264 & ~l378;
assign a6086 = ~a6084 & ~l394;
assign a6088 = a5384 & ~l386;
assign a6090 = ~a6088 & l394;
assign a6092 = ~a6090 & ~a6086;
assign a6094 = ~a6092 & a5496;
assign a6096 = ~a6094 & ~a6082;
assign a6098 = ~a6096 & ~a5492;
assign a6100 = a5024 & ~l362;
assign a6102 = ~a6100 & ~l394;
assign a6104 = a5144 & ~l370;
assign a6106 = ~a6104 & l394;
assign a6108 = ~a6106 & ~a6102;
assign a6110 = ~a6108 & a5492;
assign a6112 = ~a6110 & ~a6098;
assign a6114 = ~a6112 & ~a5488;
assign a6116 = a4784 & ~l346;
assign a6118 = ~a6116 & ~l394;
assign a6120 = a4904 & ~l354;
assign a6122 = ~a6120 & l394;
assign a6124 = ~a6122 & ~a6118;
assign a6126 = ~a6124 & a5488;
assign a6128 = ~a6126 & ~a6114;
assign a6130 = a5504 & l394;
assign a6132 = ~a6130 & ~l402;
assign a6134 = ~a5624 & l402;
assign a6136 = ~a6134 & ~a6132;
assign a6138 = ~a6136 & a5624;
assign a6140 = a6138 & ~a5616;
assign a6142 = a5264 & l378;
assign a6144 = ~a6142 & ~l402;
assign a6146 = a5384 & l386;
assign a6148 = ~a6146 & l402;
assign a6150 = ~a6148 & ~a6144;
assign a6152 = ~a6150 & a5616;
assign a6154 = ~a6152 & ~a6140;
assign a6156 = ~a6154 & ~a5612;
assign a6158 = a5024 & l362;
assign a6160 = ~a6158 & ~l402;
assign a6162 = a5144 & l370;
assign a6164 = ~a6162 & l402;
assign a6166 = ~a6164 & ~a6160;
assign a6168 = ~a6166 & a5612;
assign a6170 = ~a6168 & ~a6156;
assign a6172 = ~a6170 & ~a5608;
assign a6174 = a4784 & l346;
assign a6176 = ~a6174 & ~l402;
assign a6178 = a4904 & l354;
assign a6180 = ~a6178 & l402;
assign a6182 = ~a6180 & ~a6176;
assign a6184 = ~a6182 & a5608;
assign a6186 = ~a6184 & ~a6172;
assign a6188 = ~a5816 & ~a5812;
assign a6190 = ~a5136 & ~a5016;
assign a6192 = ~a5144 & ~a5024;
assign a6194 = ~a5616 & ~a5496;
assign a6196 = ~a6194 & ~a6192;
assign a6198 = ~a6196 & a6190;
assign a6200 = ~a6198 & a5796;
assign a6202 = ~a6198 & a5800;
assign a6204 = ~a5384 & ~a5264;
assign a6206 = ~a6204 & ~a6190;
assign a6208 = ~a6206 & a6192;
assign a6210 = ~a6208 & a5782;
assign a6212 = ~a6208 & a5786;
assign a6214 = ~a6212 & ~a6210;
assign a6216 = a6214 & ~a6202;
assign a6218 = a6216 & ~a6200;
assign a6220 = a6218 & a6188;
assign a6222 = ~a6220 & a4772;
assign a6224 = ~a5758 & ~a5754;
assign a6226 = ~a6198 & a5738;
assign a6228 = ~a6198 & a5742;
assign a6230 = ~a6208 & a5724;
assign a6232 = ~a6208 & a5728;
assign a6234 = ~a6232 & ~a6230;
assign a6236 = a6234 & ~a6228;
assign a6238 = a6236 & ~a6226;
assign a6240 = a6238 & a6224;
assign a6242 = ~a6240 & a4892;
assign a6244 = ~a5372 & ~a5252;
assign a6246 = ~a5612 & ~a5492;
assign a6248 = ~a6246 & ~a6204;
assign a6250 = ~a6248 & a6244;
assign a6252 = ~a6250 & ~a6188;
assign a6254 = ~a6244 & ~a6192;
assign a6256 = ~a6254 & a6204;
assign a6258 = ~a6256 & a5782;
assign a6260 = ~a6256 & a5786;
assign a6262 = ~a6260 & ~a6258;
assign a6264 = a6262 & ~a6252;
assign a6266 = a6264 & ~a5796;
assign a6268 = a6266 & ~a5800;
assign a6270 = ~a6268 & a4776;
assign a6272 = ~a6250 & ~a6224;
assign a6274 = ~a6256 & a5724;
assign a6276 = ~a6256 & a5728;
assign a6278 = ~a6276 & ~a6274;
assign a6280 = a6278 & ~a6272;
assign a6282 = a6280 & ~a5738;
assign a6284 = a6282 & ~a5742;
assign a6286 = ~a6284 & a4896;
assign a6288 = ~a6244 & ~a6194;
assign a6290 = ~a6288 & a6246;
assign a6292 = ~a6290 & ~a6188;
assign a6294 = ~a6246 & ~a6190;
assign a6296 = ~a6294 & a6194;
assign a6298 = ~a6296 & a5796;
assign a6300 = ~a6296 & a5800;
assign a6302 = ~a6300 & ~a6298;
assign a6304 = a6302 & ~a6292;
assign a6306 = a6304 & ~a5782;
assign a6308 = a6306 & ~a5786;
assign a6310 = ~a6308 & a4784;
assign a6312 = ~a6290 & ~a6224;
assign a6314 = ~a6296 & a5738;
assign a6316 = ~a6296 & a5742;
assign a6318 = ~a6316 & ~a6314;
assign a6320 = a6318 & ~a6312;
assign a6322 = a6320 & ~a5724;
assign a6324 = a6322 & ~a5728;
assign a6326 = ~a6324 & a4904;
assign a6328 = ~a5946 & ~a5942;
assign a6330 = ~a4896 & ~a4776;
assign a6332 = ~a4904 & ~a4784;
assign a6334 = ~a6332 & ~a6194;
assign a6336 = ~a6334 & a6330;
assign a6338 = ~a6336 & a5912;
assign a6340 = ~a6336 & a5916;
assign a6342 = ~a6330 & ~a6204;
assign a6344 = ~a6342 & a6332;
assign a6346 = ~a6344 & a5898;
assign a6348 = ~a6344 & a5902;
assign a6350 = ~a6348 & ~a6346;
assign a6352 = a6350 & ~a6340;
assign a6354 = a6352 & ~a6338;
assign a6356 = a6354 & a6328;
assign a6358 = ~a6356 & a5008;
assign a6360 = ~a5888 & ~a5884;
assign a6362 = ~a6336 & a5854;
assign a6364 = ~a6336 & a5858;
assign a6366 = ~a6344 & a5840;
assign a6368 = ~a6344 & a5844;
assign a6370 = ~a6368 & ~a6366;
assign a6372 = a6370 & ~a6364;
assign a6374 = a6372 & ~a6362;
assign a6376 = a6374 & a6360;
assign a6378 = ~a6376 & a5128;
assign a6380 = ~a5368 & ~a5248;
assign a6382 = ~a5608 & ~a5488;
assign a6384 = ~a6382 & ~a6204;
assign a6386 = ~a6384 & a6380;
assign a6388 = ~a6386 & ~a6328;
assign a6390 = ~a6380 & ~a6332;
assign a6392 = ~a6390 & a6204;
assign a6394 = ~a6392 & a5898;
assign a6396 = ~a6392 & a5902;
assign a6398 = ~a6396 & ~a6394;
assign a6400 = a6398 & ~a6388;
assign a6402 = a6400 & ~a5912;
assign a6404 = a6402 & ~a5916;
assign a6406 = ~a6404 & a5016;
assign a6408 = ~a6386 & ~a6360;
assign a6410 = ~a6392 & a5840;
assign a6412 = ~a6392 & a5844;
assign a6414 = ~a6412 & ~a6410;
assign a6416 = a6414 & ~a6408;
assign a6418 = a6416 & ~a5854;
assign a6420 = a6418 & ~a5858;
assign a6422 = ~a6420 & a5136;
assign a6424 = ~a6380 & ~a6194;
assign a6426 = ~a6424 & a6382;
assign a6428 = ~a6426 & ~a6328;
assign a6430 = ~a6382 & ~a6330;
assign a6432 = ~a6430 & a6194;
assign a6434 = ~a6432 & a5912;
assign a6436 = ~a6432 & a5916;
assign a6438 = ~a6436 & ~a6434;
assign a6440 = a6438 & ~a6428;
assign a6442 = a6440 & ~a5898;
assign a6444 = a6442 & ~a5902;
assign a6446 = ~a6444 & a5024;
assign a6448 = ~a6426 & ~a6360;
assign a6450 = ~a6432 & a5854;
assign a6452 = ~a6432 & a5858;
assign a6454 = ~a6452 & ~a6450;
assign a6456 = a6454 & ~a6448;
assign a6458 = a6456 & ~a5840;
assign a6460 = a6458 & ~a5844;
assign a6462 = ~a6460 & a5144;
assign a6464 = ~a6062 & ~a6058;
assign a6466 = ~a4892 & ~a4772;
assign a6468 = ~a6332 & ~a6246;
assign a6470 = ~a6468 & a6466;
assign a6472 = ~a6470 & a6042;
assign a6474 = ~a6470 & a6046;
assign a6476 = ~a6466 & ~a6192;
assign a6478 = ~a6476 & a6332;
assign a6480 = ~a6478 & a6014;
assign a6482 = ~a6478 & a6018;
assign a6484 = ~a6482 & ~a6480;
assign a6486 = a6484 & ~a6474;
assign a6488 = a6486 & ~a6472;
assign a6490 = a6488 & a6464;
assign a6492 = ~a6490 & a5248;
assign a6494 = ~a6004 & ~a6000;
assign a6496 = ~a6470 & a5984;
assign a6498 = ~a6470 & a5988;
assign a6500 = ~a6478 & a5956;
assign a6502 = ~a6478 & a5960;
assign a6504 = ~a6502 & ~a6500;
assign a6506 = a6504 & ~a6498;
assign a6508 = a6506 & ~a6496;
assign a6510 = a6508 & a6494;
assign a6512 = ~a6510 & a5368;
assign a6514 = ~a5128 & ~a5008;
assign a6516 = ~a6382 & ~a6192;
assign a6518 = ~a6516 & a6514;
assign a6520 = ~a6518 & ~a6464;
assign a6522 = ~a6514 & ~a6332;
assign a6524 = ~a6522 & a6192;
assign a6526 = ~a6524 & a6014;
assign a6528 = ~a6524 & a6018;
assign a6530 = ~a6528 & ~a6526;
assign a6532 = a6530 & ~a6520;
assign a6534 = a6532 & ~a6042;
assign a6536 = a6534 & ~a6046;
assign a6538 = ~a6536 & a5252;
assign a6540 = ~a6518 & ~a6494;
assign a6542 = ~a6524 & a5956;
assign a6544 = ~a6524 & a5960;
assign a6546 = ~a6544 & ~a6542;
assign a6548 = a6546 & ~a6540;
assign a6550 = a6548 & ~a5984;
assign a6552 = a6550 & ~a5988;
assign a6554 = ~a6552 & a5372;
assign a6556 = ~a6514 & ~a6246;
assign a6558 = ~a6556 & a6382;
assign a6560 = ~a6558 & ~a6464;
assign a6562 = ~a6466 & ~a6382;
assign a6564 = ~a6562 & a6246;
assign a6566 = ~a6564 & a6042;
assign a6568 = ~a6564 & a6046;
assign a6570 = ~a6568 & ~a6566;
assign a6572 = a6570 & ~a6560;
assign a6574 = a6572 & ~a6014;
assign a6576 = a6574 & ~a6018;
assign a6578 = ~a6576 & a5264;
assign a6580 = ~a6558 & ~a6494;
assign a6582 = ~a6564 & a5984;
assign a6584 = ~a6564 & a5988;
assign a6586 = ~a6584 & ~a6582;
assign a6588 = a6586 & ~a6580;
assign a6590 = a6588 & ~a5956;
assign a6592 = a6590 & ~a5960;
assign a6594 = ~a6592 & a5384;
assign a6596 = ~a6178 & ~a6174;
assign a6598 = ~a6330 & ~a6244;
assign a6600 = ~a6598 & a6466;
assign a6602 = ~a6600 & a6158;
assign a6604 = ~a6600 & a6162;
assign a6606 = ~a6466 & ~a6190;
assign a6608 = ~a6606 & a6330;
assign a6610 = ~a6608 & a6142;
assign a6612 = ~a6608 & a6146;
assign a6614 = ~a6612 & ~a6610;
assign a6616 = a6614 & ~a6604;
assign a6618 = a6616 & ~a6602;
assign a6620 = a6618 & a6596;
assign a6622 = ~a6620 & a5488;
assign a6624 = ~a6120 & ~a6116;
assign a6626 = ~a6600 & a6100;
assign a6628 = ~a6600 & a6104;
assign a6630 = ~a6608 & a6084;
assign a6632 = ~a6608 & a6088;
assign a6634 = ~a6632 & ~a6630;
assign a6636 = a6634 & ~a6628;
assign a6638 = a6636 & ~a6626;
assign a6640 = a6638 & a6624;
assign a6642 = ~a6640 & a5608;
assign a6644 = ~a6380 & ~a6190;
assign a6646 = ~a6644 & a6514;
assign a6648 = ~a6646 & ~a6596;
assign a6650 = ~a6514 & ~a6330;
assign a6652 = ~a6650 & a6190;
assign a6654 = ~a6652 & a6142;
assign a6656 = ~a6652 & a6146;
assign a6658 = ~a6656 & ~a6654;
assign a6660 = a6658 & ~a6648;
assign a6662 = a6660 & ~a6158;
assign a6664 = a6662 & ~a6162;
assign a6666 = ~a6664 & a5492;
assign a6668 = ~a6646 & ~a6624;
assign a6670 = ~a6652 & a6084;
assign a6672 = ~a6652 & a6088;
assign a6674 = ~a6672 & ~a6670;
assign a6676 = a6674 & ~a6668;
assign a6678 = a6676 & ~a6100;
assign a6680 = a6678 & ~a6104;
assign a6682 = ~a6680 & a5612;
assign a6684 = ~a6514 & ~a6244;
assign a6686 = ~a6684 & a6380;
assign a6688 = ~a6686 & ~a6596;
assign a6690 = ~a6466 & ~a6380;
assign a6692 = ~a6690 & a6244;
assign a6694 = ~a6692 & a6158;
assign a6696 = ~a6692 & a6162;
assign a6698 = ~a6696 & ~a6694;
assign a6700 = a6698 & ~a6688;
assign a6702 = a6700 & ~a6142;
assign a6704 = a6702 & ~a6146;
assign a6706 = ~a6704 & a5496;
assign a6708 = ~a6686 & ~a6624;
assign a6710 = ~a6692 & a6100;
assign a6712 = ~a6692 & a6104;
assign a6714 = ~a6712 & ~a6710;
assign a6716 = a6714 & ~a6708;
assign a6718 = a6716 & ~a6084;
assign a6720 = a6718 & ~a6088;
assign a6722 = ~a6720 & a5616;
assign a6724 = ~a6330 & a6248;
assign a6726 = ~a6332 & a6288;
assign a6728 = ~a6726 & ~a6724;
assign a6730 = a6728 & ~a6598;
assign a6732 = a6730 & ~a6468;
assign a6734 = a6732 & a6466;
assign a6736 = ~a6514 & a6334;
assign a6738 = a6430 & ~a6192;
assign a6740 = ~a6738 & ~a6736;
assign a6742 = a6740 & ~a6650;
assign a6744 = a6742 & ~a6196;
assign a6746 = a6744 & a6190;
assign a6748 = a6476 & ~a6380;
assign a6750 = a6522 & ~a6244;
assign a6752 = ~a6750 & ~a6748;
assign a6754 = a6752 & ~a6390;
assign a6756 = a6754 & ~a6254;
assign a6758 = a6756 & a6204;
assign a6760 = a4764 & l412;
assign a6762 = ~a4764 & ~l412;
assign a6764 = ~a6762 & ~a6760;
assign a6766 = a4884 & l426;
assign a6768 = ~a4884 & ~l426;
assign a6770 = ~a6768 & ~a6766;
assign a6772 = a5004 & l464;
assign a6774 = ~a5004 & ~l464;
assign a6776 = ~a6774 & ~a6772;
assign a6778 = a5124 & l478;
assign a6780 = ~a5124 & ~l478;
assign a6782 = ~a6780 & ~a6778;
assign a6784 = a5244 & l516;
assign a6786 = ~a5244 & ~l516;
assign a6788 = ~a6786 & ~a6784;
assign a6790 = a5364 & l530;
assign a6792 = ~a5364 & ~l530;
assign a6794 = ~a6792 & ~a6790;
assign a6796 = a5484 & l568;
assign a6798 = ~a5484 & ~l568;
assign a6800 = ~a6798 & ~a6796;
assign a6802 = a5604 & l582;
assign a6804 = ~a5604 & ~l582;
assign a6806 = ~a6804 & ~a6802;
assign a6808 = ~l622 & ~l410;
assign a6810 = l622 & l410;
assign a6812 = ~a6810 & ~a6808;
assign a6814 = ~l620 & l408;
assign a6816 = l620 & ~l408;
assign a6818 = ~a6816 & ~a6814;
assign a6820 = ~l626 & ~l416;
assign a6822 = l626 & l416;
assign a6824 = ~a6822 & ~a6820;
assign a6826 = ~l624 & l414;
assign a6828 = l624 & ~l414;
assign a6830 = ~a6828 & ~a6826;
assign a6832 = ~l630 & ~l424;
assign a6834 = l630 & l424;
assign a6836 = ~a6834 & ~a6832;
assign a6838 = ~l628 & l422;
assign a6840 = l628 & ~l422;
assign a6842 = ~a6840 & ~a6838;
assign a6844 = ~l634 & ~l430;
assign a6846 = l634 & l430;
assign a6848 = ~a6846 & ~a6844;
assign a6850 = ~l632 & l428;
assign a6852 = l632 & ~l428;
assign a6854 = ~a6852 & ~a6850;
assign a6856 = ~l640 & ~l436;
assign a6858 = l640 & l436;
assign a6860 = ~a6858 & ~a6856;
assign a6862 = ~l638 & l434;
assign a6864 = l638 & ~l434;
assign a6866 = ~a6864 & ~a6862;
assign a6868 = ~l636 & l432;
assign a6870 = l636 & ~l432;
assign a6872 = ~a6870 & ~a6868;
assign a6874 = ~l642 & l438;
assign a6876 = l642 & ~l438;
assign a6878 = ~a6876 & ~a6874;
assign a6880 = ~l644 & l440;
assign a6882 = l644 & ~l440;
assign a6884 = ~a6882 & ~a6880;
assign a6886 = ~l646 & l444;
assign a6888 = l646 & ~l444;
assign a6890 = ~a6888 & ~a6886;
assign a6892 = ~l648 & l446;
assign a6894 = l648 & ~l446;
assign a6896 = ~a6894 & ~a6892;
assign a6898 = ~l656 & l454;
assign a6900 = l656 & ~l454;
assign a6902 = ~a6900 & ~a6898;
assign a6904 = ~l654 & l452;
assign a6906 = l654 & ~l452;
assign a6908 = ~a6906 & ~a6904;
assign a6910 = ~l652 & l450;
assign a6912 = l652 & ~l450;
assign a6914 = ~a6912 & ~a6910;
assign a6916 = ~l650 & l448;
assign a6918 = l650 & ~l448;
assign a6920 = ~a6918 & ~a6916;
assign a6922 = ~l660 & ~l462;
assign a6924 = l660 & l462;
assign a6926 = ~a6924 & ~a6922;
assign a6928 = ~l658 & l460;
assign a6930 = l658 & ~l460;
assign a6932 = ~a6930 & ~a6928;
assign a6934 = ~l664 & ~l468;
assign a6936 = l664 & l468;
assign a6938 = ~a6936 & ~a6934;
assign a6940 = ~l662 & l466;
assign a6942 = l662 & ~l466;
assign a6944 = ~a6942 & ~a6940;
assign a6946 = ~l668 & ~l476;
assign a6948 = l668 & l476;
assign a6950 = ~a6948 & ~a6946;
assign a6952 = ~l666 & l474;
assign a6954 = l666 & ~l474;
assign a6956 = ~a6954 & ~a6952;
assign a6958 = ~l672 & ~l482;
assign a6960 = l672 & l482;
assign a6962 = ~a6960 & ~a6958;
assign a6964 = ~l670 & l480;
assign a6966 = l670 & ~l480;
assign a6968 = ~a6966 & ~a6964;
assign a6970 = ~l678 & ~l488;
assign a6972 = l678 & l488;
assign a6974 = ~a6972 & ~a6970;
assign a6976 = ~l676 & l486;
assign a6978 = l676 & ~l486;
assign a6980 = ~a6978 & ~a6976;
assign a6982 = ~l674 & l484;
assign a6984 = l674 & ~l484;
assign a6986 = ~a6984 & ~a6982;
assign a6988 = ~l680 & l490;
assign a6990 = l680 & ~l490;
assign a6992 = ~a6990 & ~a6988;
assign a6994 = ~l682 & l492;
assign a6996 = l682 & ~l492;
assign a6998 = ~a6996 & ~a6994;
assign a7000 = ~l684 & l496;
assign a7002 = l684 & ~l496;
assign a7004 = ~a7002 & ~a7000;
assign a7006 = ~l686 & l498;
assign a7008 = l686 & ~l498;
assign a7010 = ~a7008 & ~a7006;
assign a7012 = ~l694 & l506;
assign a7014 = l694 & ~l506;
assign a7016 = ~a7014 & ~a7012;
assign a7018 = ~l692 & l504;
assign a7020 = l692 & ~l504;
assign a7022 = ~a7020 & ~a7018;
assign a7024 = ~l690 & l502;
assign a7026 = l690 & ~l502;
assign a7028 = ~a7026 & ~a7024;
assign a7030 = ~l688 & l500;
assign a7032 = l688 & ~l500;
assign a7034 = ~a7032 & ~a7030;
assign a7036 = ~l698 & ~l514;
assign a7038 = l698 & l514;
assign a7040 = ~a7038 & ~a7036;
assign a7042 = ~l696 & l512;
assign a7044 = l696 & ~l512;
assign a7046 = ~a7044 & ~a7042;
assign a7048 = ~l702 & ~l520;
assign a7050 = l702 & l520;
assign a7052 = ~a7050 & ~a7048;
assign a7054 = ~l700 & l518;
assign a7056 = l700 & ~l518;
assign a7058 = ~a7056 & ~a7054;
assign a7060 = ~l706 & ~l528;
assign a7062 = l706 & l528;
assign a7064 = ~a7062 & ~a7060;
assign a7066 = ~l704 & l526;
assign a7068 = l704 & ~l526;
assign a7070 = ~a7068 & ~a7066;
assign a7072 = ~l710 & ~l534;
assign a7074 = l710 & l534;
assign a7076 = ~a7074 & ~a7072;
assign a7078 = ~l708 & l532;
assign a7080 = l708 & ~l532;
assign a7082 = ~a7080 & ~a7078;
assign a7084 = ~l716 & ~l540;
assign a7086 = l716 & l540;
assign a7088 = ~a7086 & ~a7084;
assign a7090 = ~l714 & l538;
assign a7092 = l714 & ~l538;
assign a7094 = ~a7092 & ~a7090;
assign a7096 = ~l712 & l536;
assign a7098 = l712 & ~l536;
assign a7100 = ~a7098 & ~a7096;
assign a7102 = ~l718 & l542;
assign a7104 = l718 & ~l542;
assign a7106 = ~a7104 & ~a7102;
assign a7108 = ~l720 & l544;
assign a7110 = l720 & ~l544;
assign a7112 = ~a7110 & ~a7108;
assign a7114 = ~l722 & l548;
assign a7116 = l722 & ~l548;
assign a7118 = ~a7116 & ~a7114;
assign a7120 = ~l724 & l550;
assign a7122 = l724 & ~l550;
assign a7124 = ~a7122 & ~a7120;
assign a7126 = ~l732 & l558;
assign a7128 = l732 & ~l558;
assign a7130 = ~a7128 & ~a7126;
assign a7132 = ~l730 & l556;
assign a7134 = l730 & ~l556;
assign a7136 = ~a7134 & ~a7132;
assign a7138 = ~l728 & l554;
assign a7140 = l728 & ~l554;
assign a7142 = ~a7140 & ~a7138;
assign a7144 = ~l726 & l552;
assign a7146 = l726 & ~l552;
assign a7148 = ~a7146 & ~a7144;
assign a7150 = ~l736 & ~l566;
assign a7152 = l736 & l566;
assign a7154 = ~a7152 & ~a7150;
assign a7156 = ~l734 & l564;
assign a7158 = l734 & ~l564;
assign a7160 = ~a7158 & ~a7156;
assign a7162 = ~l740 & ~l572;
assign a7164 = l740 & l572;
assign a7166 = ~a7164 & ~a7162;
assign a7168 = ~l738 & l570;
assign a7170 = l738 & ~l570;
assign a7172 = ~a7170 & ~a7168;
assign a7174 = ~l744 & ~l580;
assign a7176 = l744 & l580;
assign a7178 = ~a7176 & ~a7174;
assign a7180 = ~l742 & l578;
assign a7182 = l742 & ~l578;
assign a7184 = ~a7182 & ~a7180;
assign a7186 = ~l748 & ~l586;
assign a7188 = l748 & l586;
assign a7190 = ~a7188 & ~a7186;
assign a7192 = ~l746 & l584;
assign a7194 = l746 & ~l584;
assign a7196 = ~a7194 & ~a7192;
assign a7198 = ~l752 & l590;
assign a7200 = l752 & ~l590;
assign a7202 = ~a7200 & ~a7198;
assign a7204 = ~l750 & l588;
assign a7206 = l750 & ~l588;
assign a7208 = ~a7206 & ~a7204;
assign a7210 = ~l756 & l594;
assign a7212 = l756 & ~l594;
assign a7214 = ~a7212 & ~a7210;
assign a7216 = ~l758 & l596;
assign a7218 = l758 & ~l596;
assign a7220 = ~a7218 & ~a7216;
assign a7222 = ~l760 & l600;
assign a7224 = l760 & ~l600;
assign a7226 = ~a7224 & ~a7222;
assign a7228 = ~l762 & l602;
assign a7230 = l762 & ~l602;
assign a7232 = ~a7230 & ~a7228;
assign a7234 = ~l770 & l610;
assign a7236 = l770 & ~l610;
assign a7238 = ~a7236 & ~a7234;
assign a7240 = ~l768 & l608;
assign a7242 = l768 & ~l608;
assign a7244 = ~a7242 & ~a7240;
assign a7246 = ~l766 & l606;
assign a7248 = l766 & ~l606;
assign a7250 = ~a7248 & ~a7246;
assign a7252 = ~l764 & l604;
assign a7254 = l764 & ~l604;
assign a7256 = ~a7254 & ~a7252;
assign a7258 = ~l772 & l612;
assign a7260 = l772 & ~l612;
assign a7262 = ~a7260 & ~a7258;
assign a7264 = l774 & ~l614;
assign a7266 = ~l774 & l614;
assign a7268 = ~a7266 & ~a7264;
assign a7270 = l776 & ~l616;
assign a7272 = ~l776 & l616;
assign a7274 = ~a7272 & ~a7270;
assign a7276 = l778 & ~l618;
assign a7278 = ~l778 & l618;
assign a7280 = ~a7278 & ~a7276;
assign a7282 = a7280 & a7274;
assign a7284 = a7282 & a7268;
assign a7286 = a7284 & a7262;
assign a7288 = a7286 & a7256;
assign a7290 = a7288 & a7250;
assign a7292 = a7290 & a7244;
assign a7294 = a7292 & a7238;
assign a7296 = a7294 & a7232;
assign a7298 = a7296 & a7226;
assign a7300 = a7298 & a7220;
assign a7302 = a7300 & a7214;
assign a7304 = a7302 & a7208;
assign a7306 = a7304 & a7202;
assign a7308 = ~l754 & ~l592;
assign a7310 = l754 & l592;
assign a7312 = ~a7310 & ~a7308;
assign a7314 = a7312 & a7306;
assign a7316 = a7314 & a7196;
assign a7318 = a7316 & a7190;
assign a7320 = a7318 & a7184;
assign a7322 = a7320 & a7178;
assign a7324 = a7322 & a7172;
assign a7326 = a7324 & a7166;
assign a7328 = a7326 & a7160;
assign a7330 = a7328 & a7154;
assign a7332 = a7330 & a7148;
assign a7334 = a7332 & a7142;
assign a7336 = a7334 & a7136;
assign a7338 = a7336 & a7130;
assign a7340 = a7338 & a7124;
assign a7342 = a7340 & a7118;
assign a7344 = a7342 & a7112;
assign a7346 = a7344 & a7106;
assign a7348 = a7346 & a7100;
assign a7350 = a7348 & a7094;
assign a7352 = a7350 & a7088;
assign a7354 = a7352 & a7082;
assign a7356 = a7354 & a7076;
assign a7358 = a7356 & a7070;
assign a7360 = a7358 & a7064;
assign a7362 = a7360 & a7058;
assign a7364 = a7362 & a7052;
assign a7366 = a7364 & a7046;
assign a7368 = a7366 & a7040;
assign a7370 = a7368 & a7034;
assign a7372 = a7370 & a7028;
assign a7374 = a7372 & a7022;
assign a7376 = a7374 & a7016;
assign a7378 = a7376 & a7010;
assign a7380 = a7378 & a7004;
assign a7382 = a7380 & a6998;
assign a7384 = a7382 & a6992;
assign a7386 = a7384 & a6986;
assign a7388 = a7386 & a6980;
assign a7390 = a7388 & a6974;
assign a7392 = a7390 & a6968;
assign a7394 = a7392 & a6962;
assign a7396 = a7394 & a6956;
assign a7398 = a7396 & a6950;
assign a7400 = a7398 & a6944;
assign a7402 = a7400 & a6938;
assign a7404 = a7402 & a6932;
assign a7406 = a7404 & a6926;
assign a7408 = a7406 & a6920;
assign a7410 = a7408 & a6914;
assign a7412 = a7410 & a6908;
assign a7414 = a7412 & a6902;
assign a7416 = a7414 & a6896;
assign a7418 = a7416 & a6890;
assign a7420 = a7418 & a6884;
assign a7422 = a7420 & a6878;
assign a7424 = a7422 & a6872;
assign a7426 = a7424 & a6866;
assign a7428 = a7426 & a6860;
assign a7430 = a7428 & a6854;
assign a7432 = a7430 & a6848;
assign a7434 = a7432 & a6842;
assign a7436 = a7434 & a6836;
assign a7438 = a7436 & a6830;
assign a7440 = a7438 & a6824;
assign a7442 = a7440 & a6818;
assign a7444 = a7442 & a6812;
assign a7446 = a7444 & l788;
assign a7448 = a7446 & l780;
assign a7450 = a7448 & l782;
assign a7452 = a7450 & l784;
assign a7454 = ~a7452 & i330;
assign a7456 = ~a7454 & a6806;
assign a7458 = a7456 & a6800;
assign a7460 = a7458 & a6794;
assign a7462 = a7460 & a6788;
assign a7464 = a7462 & a6782;
assign a7466 = a7464 & a6776;
assign a7468 = a7466 & a6770;
assign a7470 = a7468 & a6764;
assign a7472 = a7470 & ~a6758;
assign a7474 = a7472 & ~a6746;
assign a7476 = a7474 & ~a6734;
assign a7478 = a7476 & ~a6722;
assign a7480 = a7478 & ~a6706;
assign a7482 = a7480 & ~a6682;
assign a7484 = a7482 & ~a6666;
assign a7486 = a7484 & ~a6642;
assign a7488 = a7486 & ~a6622;
assign a7490 = a7488 & ~a6594;
assign a7492 = a7490 & ~a6578;
assign a7494 = a7492 & ~a6554;
assign a7496 = a7494 & ~a6538;
assign a7498 = a7496 & ~a6512;
assign a7500 = a7498 & ~a6492;
assign a7502 = a7500 & ~a6462;
assign a7504 = a7502 & ~a6446;
assign a7506 = a7504 & ~a6422;
assign a7508 = a7506 & ~a6406;
assign a7510 = a7508 & ~a6378;
assign a7512 = a7510 & ~a6358;
assign a7514 = a7512 & ~a6326;
assign a7516 = a7514 & ~a6310;
assign a7518 = a7516 & ~a6286;
assign a7520 = a7518 & ~a6270;
assign a7522 = a7520 & ~a6242;
assign a7524 = a7522 & ~a6222;
assign a7526 = a7524 & a6186;
assign a7528 = a7526 & ~a5624;
assign a7530 = a7528 & a6128;
assign a7532 = a7530 & ~a5504;
assign a7534 = a7532 & a6070;
assign a7536 = a7534 & ~a5376;
assign a7538 = a7536 & a6012;
assign a7540 = a7538 & ~a5256;
assign a7542 = a7540 & a5954;
assign a7544 = a7542 & ~a5132;
assign a7546 = a7544 & a5896;
assign a7548 = a7546 & ~a5012;
assign a7550 = a7548 & a5838;
assign a7552 = a7550 & ~a4888;
assign a7554 = a7552 & a5780;
assign a7556 = a7554 & ~a4768;
assign a7558 = a7556 & ~a5722;
assign a7560 = a7558 & ~a5602;
assign a7562 = a7560 & ~a5482;
assign a7564 = a7562 & ~a5362;
assign a7566 = a7564 & ~a5242;
assign a7568 = a7566 & ~a5122;
assign a7570 = a7568 & ~a5002;
assign a7572 = a7570 & ~a4882;
assign a7574 = a7572 & ~a4762;
assign a7576 = a7574 & ~a4694;
assign a7578 = a7576 & ~a4690;
assign a7580 = a7578 & ~a4686;
assign a7582 = a7580 & ~a4684;
assign a7584 = a7582 & ~a4682;
assign a7586 = a7584 & ~a4678;
assign a7588 = a7586 & ~a4674;
assign a7590 = a7588 & ~a4672;
assign a7592 = a7590 & ~a4670;
assign a7594 = a7592 & ~a4666;
assign a7596 = a7594 & ~a4662;
assign a7598 = a7596 & ~a4660;
assign a7600 = a7598 & ~a4658;
assign a7602 = a7600 & ~a4654;
assign a7604 = a7602 & ~a4650;
assign a7606 = a7604 & ~a4648;
assign a7608 = a7606 & ~a4646;
assign a7610 = a7608 & ~a4644;
assign a7612 = a7610 & ~a4642;
assign a7614 = a7612 & ~a4640;
assign a7616 = a7614 & ~a4638;
assign a7618 = a7616 & ~a4636;
assign a7620 = a7618 & ~a4634;
assign a7622 = a7620 & ~a4632;
assign a7624 = a7622 & ~a4630;
assign a7626 = a7624 & ~a4628;
assign a7628 = a7626 & ~a4626;
assign a7630 = a7628 & ~a4624;
assign a7632 = a7630 & ~a4622;
assign a7634 = a7632 & ~a4620;
assign a7636 = a7634 & ~a4618;
assign a7638 = a7636 & ~a4616;
assign a7640 = a7638 & ~a4614;
assign a7642 = a7640 & ~a4612;
assign a7644 = a7642 & ~a4610;
assign a7646 = a7644 & ~a4608;
assign a7648 = a7646 & ~a4606;
assign a7650 = a7648 & ~a4604;
assign a7652 = a7650 & ~a4602;
assign a7654 = a7652 & ~a4600;
assign a7656 = a7654 & ~a4598;
assign a7658 = a7656 & ~a4594;
assign a7660 = a7658 & ~a4590;
assign a7662 = a7660 & ~a4586;
assign a7664 = a7662 & ~a4582;
assign a7666 = a7664 & ~a4578;
assign a7668 = a7666 & ~a4574;
assign a7670 = a7668 & ~a4570;
assign a7672 = a7670 & l798;
assign a7674 = a7672 & a4566;
assign a7678 = a7672 & i330;
assign p0 = a7678;

assert property (~p0);

endmodule
