module m139443p (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474;

output p0;

wire a1154,a1170,a1198,a1242,a1258,a1278,a1322,a1338,a1358,a1442,a1466,a1492,a1504,a1658,a1668,
a1678,a1688,a1746,a1762,a1790,a1834,a1850,a1870,a1914,a1930,a1950,a2034,a2058,a2084,a2096,
a2250,a2260,a2270,a2280,a2338,a2354,a2382,a2426,a2442,a2462,a2506,a2522,a2542,a2626,a2650,
a2676,a2688,a2842,a2852,a2862,a2872,a2930,a2946,a2974,a3018,a3034,a3054,a3098,a3114,a3134,
a3218,a3242,a3268,a3280,a3434,a3444,a3454,a3464,a3470,a3478,a3488,a3496,a3498,a11940,c1,
a1098,a1100,a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,a1124,a1126,
a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,a1156,a1158,
a1160,a1162,a1164,a1166,a1168,a1172,a1174,a1176,a1178,a1180,a1182,a1184,a1186,a1188,a1190,
a1192,a1194,a1196,a1200,a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,a1218,a1220,a1222,
a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1244,a1246,a1248,a1250,a1252,a1254,
a1256,a1260,a1262,a1264,a1266,a1268,a1270,a1272,a1274,a1276,a1280,a1282,a1284,a1286,a1288,
a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,a1310,a1312,a1314,a1316,a1318,
a1320,a1324,a1326,a1328,a1330,a1332,a1334,a1336,a1340,a1342,a1344,a1346,a1348,a1350,a1352,
a1354,a1356,a1360,a1362,a1364,a1366,a1368,a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,
a1386,a1388,a1390,a1392,a1394,a1396,a1398,a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,
a1416,a1418,a1420,a1422,a1424,a1426,a1428,a1430,a1432,a1434,a1436,a1438,a1440,a1444,a1446,
a1448,a1450,a1452,a1454,a1456,a1458,a1460,a1462,a1464,a1468,a1470,a1472,a1474,a1476,a1478,
a1480,a1482,a1484,a1486,a1488,a1490,a1494,a1496,a1498,a1500,a1502,a1506,a1508,a1510,a1512,
a1514,a1516,a1518,a1520,a1522,a1524,a1526,a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,
a1544,a1546,a1548,a1550,a1552,a1554,a1556,a1558,a1560,a1562,a1564,a1566,a1568,a1570,a1572,
a1574,a1576,a1578,a1580,a1582,a1584,a1586,a1588,a1590,a1592,a1594,a1596,a1598,a1600,a1602,
a1604,a1606,a1608,a1610,a1612,a1614,a1616,a1618,a1620,a1622,a1624,a1626,a1628,a1630,a1632,
a1634,a1636,a1638,a1640,a1642,a1644,a1646,a1648,a1650,a1652,a1654,a1656,a1660,a1662,a1664,
a1666,a1670,a1672,a1674,a1676,a1680,a1682,a1684,a1686,a1690,a1692,a1694,a1696,a1698,a1700,
a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,
a1732,a1734,a1736,a1738,a1740,a1742,a1744,a1748,a1750,a1752,a1754,a1756,a1758,a1760,a1764,
a1766,a1768,a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,a1792,a1794,a1796,
a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,a1822,a1824,a1826,
a1828,a1830,a1832,a1836,a1838,a1840,a1842,a1844,a1846,a1848,a1852,a1854,a1856,a1858,a1860,
a1862,a1864,a1866,a1868,a1872,a1874,a1876,a1878,a1880,a1882,a1884,a1886,a1888,a1890,a1892,
a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,a1910,a1912,a1916,a1918,a1920,a1922,a1924,
a1926,a1928,a1932,a1934,a1936,a1938,a1940,a1942,a1944,a1946,a1948,a1952,a1954,a1956,a1958,
a1960,a1962,a1964,a1966,a1968,a1970,a1972,a1974,a1976,a1978,a1980,a1982,a1984,a1986,a1988,
a1990,a1992,a1994,a1996,a1998,a2000,a2002,a2004,a2006,a2008,a2010,a2012,a2014,a2016,a2018,
a2020,a2022,a2024,a2026,a2028,a2030,a2032,a2036,a2038,a2040,a2042,a2044,a2046,a2048,a2050,
a2052,a2054,a2056,a2060,a2062,a2064,a2066,a2068,a2070,a2072,a2074,a2076,a2078,a2080,a2082,
a2086,a2088,a2090,a2092,a2094,a2098,a2100,a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,
a2118,a2120,a2122,a2124,a2126,a2128,a2130,a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,
a2148,a2150,a2152,a2154,a2156,a2158,a2160,a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,
a2178,a2180,a2182,a2184,a2186,a2188,a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,
a2208,a2210,a2212,a2214,a2216,a2218,a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,
a2238,a2240,a2242,a2244,a2246,a2248,a2252,a2254,a2256,a2258,a2262,a2264,a2266,a2268,a2272,
a2274,a2276,a2278,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,a2298,a2300,a2302,a2304,
a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,a2328,a2330,a2332,a2334,
a2336,a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2356,a2358,a2360,a2362,a2364,a2366,a2368,
a2370,a2372,a2374,a2376,a2378,a2380,a2384,a2386,a2388,a2390,a2392,a2394,a2396,a2398,a2400,
a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,a2420,a2422,a2424,a2428,a2430,a2432,
a2434,a2436,a2438,a2440,a2444,a2446,a2448,a2450,a2452,a2454,a2456,a2458,a2460,a2464,a2466,
a2468,a2470,a2472,a2474,a2476,a2478,a2480,a2482,a2484,a2486,a2488,a2490,a2492,a2494,a2496,
a2498,a2500,a2502,a2504,a2508,a2510,a2512,a2514,a2516,a2518,a2520,a2524,a2526,a2528,a2530,
a2532,a2534,a2536,a2538,a2540,a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,
a2564,a2566,a2568,a2570,a2572,a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,
a2594,a2596,a2598,a2600,a2602,a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,
a2624,a2628,a2630,a2632,a2634,a2636,a2638,a2640,a2642,a2644,a2646,a2648,a2652,a2654,a2656,
a2658,a2660,a2662,a2664,a2666,a2668,a2670,a2672,a2674,a2678,a2680,a2682,a2684,a2686,a2690,
a2692,a2694,a2696,a2698,a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,a2718,a2720,
a2722,a2724,a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,
a2752,a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,
a2782,a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,a2810,
a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,a2840,
a2844,a2846,a2848,a2850,a2854,a2856,a2858,a2860,a2864,a2866,a2868,a2870,a2874,a2876,a2878,
a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,a2900,a2902,a2904,a2906,a2908,
a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2932,a2934,a2936,a2938,a2940,
a2942,a2944,a2948,a2950,a2952,a2954,a2956,a2958,a2960,a2962,a2964,a2966,a2968,a2970,a2972,
a2976,a2978,a2980,a2982,a2984,a2986,a2988,a2990,a2992,a2994,a2996,a2998,a3000,a3002,a3004,
a3006,a3008,a3010,a3012,a3014,a3016,a3020,a3022,a3024,a3026,a3028,a3030,a3032,a3036,a3038,
a3040,a3042,a3044,a3046,a3048,a3050,a3052,a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,
a3072,a3074,a3076,a3078,a3080,a3082,a3084,a3086,a3088,a3090,a3092,a3094,a3096,a3100,a3102,
a3104,a3106,a3108,a3110,a3112,a3116,a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3136,
a3138,a3140,a3142,a3144,a3146,a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,
a3168,a3170,a3172,a3174,a3176,a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,
a3198,a3200,a3202,a3204,a3206,a3208,a3210,a3212,a3214,a3216,a3220,a3222,a3224,a3226,a3228,
a3230,a3232,a3234,a3236,a3238,a3240,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,
a3262,a3264,a3266,a3270,a3272,a3274,a3276,a3278,a3282,a3284,a3286,a3288,a3290,a3292,a3294,
a3296,a3298,a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,a3324,
a3326,a3328,a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,a3354,
a3356,a3358,a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3382,a3384,
a3386,a3388,a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,a3408,a3410,a3412,a3414,
a3416,a3418,a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3436,a3438,a3440,a3442,a3446,a3448,
a3450,a3452,a3456,a3458,a3460,a3462,a3466,a3468,a3472,a3474,a3476,a3480,a3482,a3484,a3486,
a3490,a3492,a3494,a3500,a3502,a3504,a3506,a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,
a3524,a3526,a3528,a3530,a3532,a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,
a3554,a3556,a3558,a3560,a3562,a3564,a3566,a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,
a3584,a3586,a3588,a3590,a3592,a3594,a3596,a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3612,
a3614,a3616,a3618,a3620,a3622,a3624,a3626,a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,
a3644,a3646,a3648,a3650,a3652,a3654,a3656,a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,
a3674,a3676,a3678,a3680,a3682,a3684,a3686,a3688,a3690,a3692,a3694,a3696,a3698,a3700,a3702,
a3704,a3706,a3708,a3710,a3712,a3714,a3716,a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,
a3734,a3736,a3738,a3740,a3742,a3744,a3746,a3748,a3750,a3752,a3754,a3756,a3758,a3760,a3762,
a3764,a3766,a3768,a3770,a3772,a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,a3790,a3792,
a3794,a3796,a3798,a3800,a3802,a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,
a3824,a3826,a3828,a3830,a3832,a3834,a3836,a3838,a3840,a3842,a3844,a3846,a3848,a3850,a3852,
a3854,a3856,a3858,a3860,a3862,a3864,a3866,a3868,a3870,a3872,a3874,a3876,a3878,a3880,a3882,
a3884,a3886,a3888,a3890,a3892,a3894,a3896,a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,
a3914,a3916,a3918,a3920,a3922,a3924,a3926,a3928,a3930,a3932,a3934,a3936,a3938,a3940,a3942,
a3944,a3946,a3948,a3950,a3952,a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,
a3974,a3976,a3978,a3980,a3982,a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,
a4004,a4006,a4008,a4010,a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,
a4034,a4036,a4038,a4040,a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,
a4064,a4066,a4068,a4070,a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,
a4094,a4096,a4098,a4100,a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,
a4124,a4126,a4128,a4130,a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,a4152,
a4154,a4156,a4158,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,
a4184,a4186,a4188,a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,
a4214,a4216,a4218,a4220,a4222,a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,
a4244,a4246,a4248,a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,
a4274,a4276,a4278,a4280,a4282,a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,
a4304,a4306,a4308,a4310,a4312,a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,
a4334,a4336,a4338,a4340,a4342,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,
a4364,a4366,a4368,a4370,a4372,a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,
a4394,a4396,a4398,a4400,a4402,a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,
a4424,a4426,a4428,a4430,a4432,a4434,a4436,a4438,a4440,a4442,a4444,a4446,a4448,a4450,a4452,
a4454,a4456,a4458,a4460,a4462,a4464,a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4482,
a4484,a4486,a4488,a4490,a4492,a4494,a4496,a4498,a4500,a4502,a4504,a4506,a4508,a4510,a4512,
a4514,a4516,a4518,a4520,a4522,a4524,a4526,a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,
a4544,a4546,a4548,a4550,a4552,a4554,a4556,a4558,a4560,a4562,a4564,a4566,a4568,a4570,a4572,
a4574,a4576,a4578,a4580,a4582,a4584,a4586,a4588,a4590,a4592,a4594,a4596,a4598,a4600,a4602,
a4604,a4606,a4608,a4610,a4612,a4614,a4616,a4618,a4620,a4622,a4624,a4626,a4628,a4630,a4632,
a4634,a4636,a4638,a4640,a4642,a4644,a4646,a4648,a4650,a4652,a4654,a4656,a4658,a4660,a4662,
a4664,a4666,a4668,a4670,a4672,a4674,a4676,a4678,a4680,a4682,a4684,a4686,a4688,a4690,a4692,
a4694,a4696,a4698,a4700,a4702,a4704,a4706,a4708,a4710,a4712,a4714,a4716,a4718,a4720,a4722,
a4724,a4726,a4728,a4730,a4732,a4734,a4736,a4738,a4740,a4742,a4744,a4746,a4748,a4750,a4752,
a4754,a4756,a4758,a4760,a4762,a4764,a4766,a4768,a4770,a4772,a4774,a4776,a4778,a4780,a4782,
a4784,a4786,a4788,a4790,a4792,a4794,a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,a4812,
a4814,a4816,a4818,a4820,a4822,a4824,a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,
a4844,a4846,a4848,a4850,a4852,a4854,a4856,a4858,a4860,a4862,a4864,a4866,a4868,a4870,a4872,
a4874,a4876,a4878,a4880,a4882,a4884,a4886,a4888,a4890,a4892,a4894,a4896,a4898,a4900,a4902,
a4904,a4906,a4908,a4910,a4912,a4914,a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,
a4934,a4936,a4938,a4940,a4942,a4944,a4946,a4948,a4950,a4952,a4954,a4956,a4958,a4960,a4962,
a4964,a4966,a4968,a4970,a4972,a4974,a4976,a4978,a4980,a4982,a4984,a4986,a4988,a4990,a4992,
a4994,a4996,a4998,a5000,a5002,a5004,a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,a5022,
a5024,a5026,a5028,a5030,a5032,a5034,a5036,a5038,a5040,a5042,a5044,a5046,a5048,a5050,a5052,
a5054,a5056,a5058,a5060,a5062,a5064,a5066,a5068,a5070,a5072,a5074,a5076,a5078,a5080,a5082,
a5084,a5086,a5088,a5090,a5092,a5094,a5096,a5098,a5100,a5102,a5104,a5106,a5108,a5110,a5112,
a5114,a5116,a5118,a5120,a5122,a5124,a5126,a5128,a5130,a5132,a5134,a5136,a5138,a5140,a5142,
a5144,a5146,a5148,a5150,a5152,a5154,a5156,a5158,a5160,a5162,a5164,a5166,a5168,a5170,a5172,
a5174,a5176,a5178,a5180,a5182,a5184,a5186,a5188,a5190,a5192,a5194,a5196,a5198,a5200,a5202,
a5204,a5206,a5208,a5210,a5212,a5214,a5216,a5218,a5220,a5222,a5224,a5226,a5228,a5230,a5232,
a5234,a5236,a5238,a5240,a5242,a5244,a5246,a5248,a5250,a5252,a5254,a5256,a5258,a5260,a5262,
a5264,a5266,a5268,a5270,a5272,a5274,a5276,a5278,a5280,a5282,a5284,a5286,a5288,a5290,a5292,
a5294,a5296,a5298,a5300,a5302,a5304,a5306,a5308,a5310,a5312,a5314,a5316,a5318,a5320,a5322,
a5324,a5326,a5328,a5330,a5332,a5334,a5336,a5338,a5340,a5342,a5344,a5346,a5348,a5350,a5352,
a5354,a5356,a5358,a5360,a5362,a5364,a5366,a5368,a5370,a5372,a5374,a5376,a5378,a5380,a5382,
a5384,a5386,a5388,a5390,a5392,a5394,a5396,a5398,a5400,a5402,a5404,a5406,a5408,a5410,a5412,
a5414,a5416,a5418,a5420,a5422,a5424,a5426,a5428,a5430,a5432,a5434,a5436,a5438,a5440,a5442,
a5444,a5446,a5448,a5450,a5452,a5454,a5456,a5458,a5460,a5462,a5464,a5466,a5468,a5470,a5472,
a5474,a5476,a5478,a5480,a5482,a5484,a5486,a5488,a5490,a5492,a5494,a5496,a5498,a5500,a5502,
a5504,a5506,a5508,a5510,a5512,a5514,a5516,a5518,a5520,a5522,a5524,a5526,a5528,a5530,a5532,
a5534,a5536,a5538,a5540,a5542,a5544,a5546,a5548,a5550,a5552,a5554,a5556,a5558,a5560,a5562,
a5564,a5566,a5568,a5570,a5572,a5574,a5576,a5578,a5580,a5582,a5584,a5586,a5588,a5590,a5592,
a5594,a5596,a5598,a5600,a5602,a5604,a5606,a5608,a5610,a5612,a5614,a5616,a5618,a5620,a5622,
a5624,a5626,a5628,a5630,a5632,a5634,a5636,a5638,a5640,a5642,a5644,a5646,a5648,a5650,a5652,
a5654,a5656,a5658,a5660,a5662,a5664,a5666,a5668,a5670,a5672,a5674,a5676,a5678,a5680,a5682,
a5684,a5686,a5688,a5690,a5692,a5694,a5696,a5698,a5700,a5702,a5704,a5706,a5708,a5710,a5712,
a5714,a5716,a5718,a5720,a5722,a5724,a5726,a5728,a5730,a5732,a5734,a5736,a5738,a5740,a5742,
a5744,a5746,a5748,a5750,a5752,a5754,a5756,a5758,a5760,a5762,a5764,a5766,a5768,a5770,a5772,
a5774,a5776,a5778,a5780,a5782,a5784,a5786,a5788,a5790,a5792,a5794,a5796,a5798,a5800,a5802,
a5804,a5806,a5808,a5810,a5812,a5814,a5816,a5818,a5820,a5822,a5824,a5826,a5828,a5830,a5832,
a5834,a5836,a5838,a5840,a5842,a5844,a5846,a5848,a5850,a5852,a5854,a5856,a5858,a5860,a5862,
a5864,a5866,a5868,a5870,a5872,a5874,a5876,a5878,a5880,a5882,a5884,a5886,a5888,a5890,a5892,
a5894,a5896,a5898,a5900,a5902,a5904,a5906,a5908,a5910,a5912,a5914,a5916,a5918,a5920,a5922,
a5924,a5926,a5928,a5930,a5932,a5934,a5936,a5938,a5940,a5942,a5944,a5946,a5948,a5950,a5952,
a5954,a5956,a5958,a5960,a5962,a5964,a5966,a5968,a5970,a5972,a5974,a5976,a5978,a5980,a5982,
a5984,a5986,a5988,a5990,a5992,a5994,a5996,a5998,a6000,a6002,a6004,a6006,a6008,a6010,a6012,
a6014,a6016,a6018,a6020,a6022,a6024,a6026,a6028,a6030,a6032,a6034,a6036,a6038,a6040,a6042,
a6044,a6046,a6048,a6050,a6052,a6054,a6056,a6058,a6060,a6062,a6064,a6066,a6068,a6070,a6072,
a6074,a6076,a6078,a6080,a6082,a6084,a6086,a6088,a6090,a6092,a6094,a6096,a6098,a6100,a6102,
a6104,a6106,a6108,a6110,a6112,a6114,a6116,a6118,a6120,a6122,a6124,a6126,a6128,a6130,a6132,
a6134,a6136,a6138,a6140,a6142,a6144,a6146,a6148,a6150,a6152,a6154,a6156,a6158,a6160,a6162,
a6164,a6166,a6168,a6170,a6172,a6174,a6176,a6178,a6180,a6182,a6184,a6186,a6188,a6190,a6192,
a6194,a6196,a6198,a6200,a6202,a6204,a6206,a6208,a6210,a6212,a6214,a6216,a6218,a6220,a6222,
a6224,a6226,a6228,a6230,a6232,a6234,a6236,a6238,a6240,a6242,a6244,a6246,a6248,a6250,a6252,
a6254,a6256,a6258,a6260,a6262,a6264,a6266,a6268,a6270,a6272,a6274,a6276,a6278,a6280,a6282,
a6284,a6286,a6288,a6290,a6292,a6294,a6296,a6298,a6300,a6302,a6304,a6306,a6308,a6310,a6312,
a6314,a6316,a6318,a6320,a6322,a6324,a6326,a6328,a6330,a6332,a6334,a6336,a6338,a6340,a6342,
a6344,a6346,a6348,a6350,a6352,a6354,a6356,a6358,a6360,a6362,a6364,a6366,a6368,a6370,a6372,
a6374,a6376,a6378,a6380,a6382,a6384,a6386,a6388,a6390,a6392,a6394,a6396,a6398,a6400,a6402,
a6404,a6406,a6408,a6410,a6412,a6414,a6416,a6418,a6420,a6422,a6424,a6426,a6428,a6430,a6432,
a6434,a6436,a6438,a6440,a6442,a6444,a6446,a6448,a6450,a6452,a6454,a6456,a6458,a6460,a6462,
a6464,a6466,a6468,a6470,a6472,a6474,a6476,a6478,a6480,a6482,a6484,a6486,a6488,a6490,a6492,
a6494,a6496,a6498,a6500,a6502,a6504,a6506,a6508,a6510,a6512,a6514,a6516,a6518,a6520,a6522,
a6524,a6526,a6528,a6530,a6532,a6534,a6536,a6538,a6540,a6542,a6544,a6546,a6548,a6550,a6552,
a6554,a6556,a6558,a6560,a6562,a6564,a6566,a6568,a6570,a6572,a6574,a6576,a6578,a6580,a6582,
a6584,a6586,a6588,a6590,a6592,a6594,a6596,a6598,a6600,a6602,a6604,a6606,a6608,a6610,a6612,
a6614,a6616,a6618,a6620,a6622,a6624,a6626,a6628,a6630,a6632,a6634,a6636,a6638,a6640,a6642,
a6644,a6646,a6648,a6650,a6652,a6654,a6656,a6658,a6660,a6662,a6664,a6666,a6668,a6670,a6672,
a6674,a6676,a6678,a6680,a6682,a6684,a6686,a6688,a6690,a6692,a6694,a6696,a6698,a6700,a6702,
a6704,a6706,a6708,a6710,a6712,a6714,a6716,a6718,a6720,a6722,a6724,a6726,a6728,a6730,a6732,
a6734,a6736,a6738,a6740,a6742,a6744,a6746,a6748,a6750,a6752,a6754,a6756,a6758,a6760,a6762,
a6764,a6766,a6768,a6770,a6772,a6774,a6776,a6778,a6780,a6782,a6784,a6786,a6788,a6790,a6792,
a6794,a6796,a6798,a6800,a6802,a6804,a6806,a6808,a6810,a6812,a6814,a6816,a6818,a6820,a6822,
a6824,a6826,a6828,a6830,a6832,a6834,a6836,a6838,a6840,a6842,a6844,a6846,a6848,a6850,a6852,
a6854,a6856,a6858,a6860,a6862,a6864,a6866,a6868,a6870,a6872,a6874,a6876,a6878,a6880,a6882,
a6884,a6886,a6888,a6890,a6892,a6894,a6896,a6898,a6900,a6902,a6904,a6906,a6908,a6910,a6912,
a6914,a6916,a6918,a6920,a6922,a6924,a6926,a6928,a6930,a6932,a6934,a6936,a6938,a6940,a6942,
a6944,a6946,a6948,a6950,a6952,a6954,a6956,a6958,a6960,a6962,a6964,a6966,a6968,a6970,a6972,
a6974,a6976,a6978,a6980,a6982,a6984,a6986,a6988,a6990,a6992,a6994,a6996,a6998,a7000,a7002,
a7004,a7006,a7008,a7010,a7012,a7014,a7016,a7018,a7020,a7022,a7024,a7026,a7028,a7030,a7032,
a7034,a7036,a7038,a7040,a7042,a7044,a7046,a7048,a7050,a7052,a7054,a7056,a7058,a7060,a7062,
a7064,a7066,a7068,a7070,a7072,a7074,a7076,a7078,a7080,a7082,a7084,a7086,a7088,a7090,a7092,
a7094,a7096,a7098,a7100,a7102,a7104,a7106,a7108,a7110,a7112,a7114,a7116,a7118,a7120,a7122,
a7124,a7126,a7128,a7130,a7132,a7134,a7136,a7138,a7140,a7142,a7144,a7146,a7148,a7150,a7152,
a7154,a7156,a7158,a7160,a7162,a7164,a7166,a7168,a7170,a7172,a7174,a7176,a7178,a7180,a7182,
a7184,a7186,a7188,a7190,a7192,a7194,a7196,a7198,a7200,a7202,a7204,a7206,a7208,a7210,a7212,
a7214,a7216,a7218,a7220,a7222,a7224,a7226,a7228,a7230,a7232,a7234,a7236,a7238,a7240,a7242,
a7244,a7246,a7248,a7250,a7252,a7254,a7256,a7258,a7260,a7262,a7264,a7266,a7268,a7270,a7272,
a7274,a7276,a7278,a7280,a7282,a7284,a7286,a7288,a7290,a7292,a7294,a7296,a7298,a7300,a7302,
a7304,a7306,a7308,a7310,a7312,a7314,a7316,a7318,a7320,a7322,a7324,a7326,a7328,a7330,a7332,
a7334,a7336,a7338,a7340,a7342,a7344,a7346,a7348,a7350,a7352,a7354,a7356,a7358,a7360,a7362,
a7364,a7366,a7368,a7370,a7372,a7374,a7376,a7378,a7380,a7382,a7384,a7386,a7388,a7390,a7392,
a7394,a7396,a7398,a7400,a7402,a7404,a7406,a7408,a7410,a7412,a7414,a7416,a7418,a7420,a7422,
a7424,a7426,a7428,a7430,a7432,a7434,a7436,a7438,a7440,a7442,a7444,a7446,a7448,a7450,a7452,
a7454,a7456,a7458,a7460,a7462,a7464,a7466,a7468,a7470,a7472,a7474,a7476,a7478,a7480,a7482,
a7484,a7486,a7488,a7490,a7492,a7494,a7496,a7498,a7500,a7502,a7504,a7506,a7508,a7510,a7512,
a7514,a7516,a7518,a7520,a7522,a7524,a7526,a7528,a7530,a7532,a7534,a7536,a7538,a7540,a7542,
a7544,a7546,a7548,a7550,a7552,a7554,a7556,a7558,a7560,a7562,a7564,a7566,a7568,a7570,a7572,
a7574,a7576,a7578,a7580,a7582,a7584,a7586,a7588,a7590,a7592,a7594,a7596,a7598,a7600,a7602,
a7604,a7606,a7608,a7610,a7612,a7614,a7616,a7618,a7620,a7622,a7624,a7626,a7628,a7630,a7632,
a7634,a7636,a7638,a7640,a7642,a7644,a7646,a7648,a7650,a7652,a7654,a7656,a7658,a7660,a7662,
a7664,a7666,a7668,a7670,a7672,a7674,a7676,a7678,a7680,a7682,a7684,a7686,a7688,a7690,a7692,
a7694,a7696,a7698,a7700,a7702,a7704,a7706,a7708,a7710,a7712,a7714,a7716,a7718,a7720,a7722,
a7724,a7726,a7728,a7730,a7732,a7734,a7736,a7738,a7740,a7742,a7744,a7746,a7748,a7750,a7752,
a7754,a7756,a7758,a7760,a7762,a7764,a7766,a7768,a7770,a7772,a7774,a7776,a7778,a7780,a7782,
a7784,a7786,a7788,a7790,a7792,a7794,a7796,a7798,a7800,a7802,a7804,a7806,a7808,a7810,a7812,
a7814,a7816,a7818,a7820,a7822,a7824,a7826,a7828,a7830,a7832,a7834,a7836,a7838,a7840,a7842,
a7844,a7846,a7848,a7850,a7852,a7854,a7856,a7858,a7860,a7862,a7864,a7866,a7868,a7870,a7872,
a7874,a7876,a7878,a7880,a7882,a7884,a7886,a7888,a7890,a7892,a7894,a7896,a7898,a7900,a7902,
a7904,a7906,a7908,a7910,a7912,a7914,a7916,a7918,a7920,a7922,a7924,a7926,a7928,a7930,a7932,
a7934,a7936,a7938,a7940,a7942,a7944,a7946,a7948,a7950,a7952,a7954,a7956,a7958,a7960,a7962,
a7964,a7966,a7968,a7970,a7972,a7974,a7976,a7978,a7980,a7982,a7984,a7986,a7988,a7990,a7992,
a7994,a7996,a7998,a8000,a8002,a8004,a8006,a8008,a8010,a8012,a8014,a8016,a8018,a8020,a8022,
a8024,a8026,a8028,a8030,a8032,a8034,a8036,a8038,a8040,a8042,a8044,a8046,a8048,a8050,a8052,
a8054,a8056,a8058,a8060,a8062,a8064,a8066,a8068,a8070,a8072,a8074,a8076,a8078,a8080,a8082,
a8084,a8086,a8088,a8090,a8092,a8094,a8096,a8098,a8100,a8102,a8104,a8106,a8108,a8110,a8112,
a8114,a8116,a8118,a8120,a8122,a8124,a8126,a8128,a8130,a8132,a8134,a8136,a8138,a8140,a8142,
a8144,a8146,a8148,a8150,a8152,a8154,a8156,a8158,a8160,a8162,a8164,a8166,a8168,a8170,a8172,
a8174,a8176,a8178,a8180,a8182,a8184,a8186,a8188,a8190,a8192,a8194,a8196,a8198,a8200,a8202,
a8204,a8206,a8208,a8210,a8212,a8214,a8216,a8218,a8220,a8222,a8224,a8226,a8228,a8230,a8232,
a8234,a8236,a8238,a8240,a8242,a8244,a8246,a8248,a8250,a8252,a8254,a8256,a8258,a8260,a8262,
a8264,a8266,a8268,a8270,a8272,a8274,a8276,a8278,a8280,a8282,a8284,a8286,a8288,a8290,a8292,
a8294,a8296,a8298,a8300,a8302,a8304,a8306,a8308,a8310,a8312,a8314,a8316,a8318,a8320,a8322,
a8324,a8326,a8328,a8330,a8332,a8334,a8336,a8338,a8340,a8342,a8344,a8346,a8348,a8350,a8352,
a8354,a8356,a8358,a8360,a8362,a8364,a8366,a8368,a8370,a8372,a8374,a8376,a8378,a8380,a8382,
a8384,a8386,a8388,a8390,a8392,a8394,a8396,a8398,a8400,a8402,a8404,a8406,a8408,a8410,a8412,
a8414,a8416,a8418,a8420,a8422,a8424,a8426,a8428,a8430,a8432,a8434,a8436,a8438,a8440,a8442,
a8444,a8446,a8448,a8450,a8452,a8454,a8456,a8458,a8460,a8462,a8464,a8466,a8468,a8470,a8472,
a8474,a8476,a8478,a8480,a8482,a8484,a8486,a8488,a8490,a8492,a8494,a8496,a8498,a8500,a8502,
a8504,a8506,a8508,a8510,a8512,a8514,a8516,a8518,a8520,a8522,a8524,a8526,a8528,a8530,a8532,
a8534,a8536,a8538,a8540,a8542,a8544,a8546,a8548,a8550,a8552,a8554,a8556,a8558,a8560,a8562,
a8564,a8566,a8568,a8570,a8572,a8574,a8576,a8578,a8580,a8582,a8584,a8586,a8588,a8590,a8592,
a8594,a8596,a8598,a8600,a8602,a8604,a8606,a8608,a8610,a8612,a8614,a8616,a8618,a8620,a8622,
a8624,a8626,a8628,a8630,a8632,a8634,a8636,a8638,a8640,a8642,a8644,a8646,a8648,a8650,a8652,
a8654,a8656,a8658,a8660,a8662,a8664,a8666,a8668,a8670,a8672,a8674,a8676,a8678,a8680,a8682,
a8684,a8686,a8688,a8690,a8692,a8694,a8696,a8698,a8700,a8702,a8704,a8706,a8708,a8710,a8712,
a8714,a8716,a8718,a8720,a8722,a8724,a8726,a8728,a8730,a8732,a8734,a8736,a8738,a8740,a8742,
a8744,a8746,a8748,a8750,a8752,a8754,a8756,a8758,a8760,a8762,a8764,a8766,a8768,a8770,a8772,
a8774,a8776,a8778,a8780,a8782,a8784,a8786,a8788,a8790,a8792,a8794,a8796,a8798,a8800,a8802,
a8804,a8806,a8808,a8810,a8812,a8814,a8816,a8818,a8820,a8822,a8824,a8826,a8828,a8830,a8832,
a8834,a8836,a8838,a8840,a8842,a8844,a8846,a8848,a8850,a8852,a8854,a8856,a8858,a8860,a8862,
a8864,a8866,a8868,a8870,a8872,a8874,a8876,a8878,a8880,a8882,a8884,a8886,a8888,a8890,a8892,
a8894,a8896,a8898,a8900,a8902,a8904,a8906,a8908,a8910,a8912,a8914,a8916,a8918,a8920,a8922,
a8924,a8926,a8928,a8930,a8932,a8934,a8936,a8938,a8940,a8942,a8944,a8946,a8948,a8950,a8952,
a8954,a8956,a8958,a8960,a8962,a8964,a8966,a8968,a8970,a8972,a8974,a8976,a8978,a8980,a8982,
a8984,a8986,a8988,a8990,a8992,a8994,a8996,a8998,a9000,a9002,a9004,a9006,a9008,a9010,a9012,
a9014,a9016,a9018,a9020,a9022,a9024,a9026,a9028,a9030,a9032,a9034,a9036,a9038,a9040,a9042,
a9044,a9046,a9048,a9050,a9052,a9054,a9056,a9058,a9060,a9062,a9064,a9066,a9068,a9070,a9072,
a9074,a9076,a9078,a9080,a9082,a9084,a9086,a9088,a9090,a9092,a9094,a9096,a9098,a9100,a9102,
a9104,a9106,a9108,a9110,a9112,a9114,a9116,a9118,a9120,a9122,a9124,a9126,a9128,a9130,a9132,
a9134,a9136,a9138,a9140,a9142,a9144,a9146,a9148,a9150,a9152,a9154,a9156,a9158,a9160,a9162,
a9164,a9166,a9168,a9170,a9172,a9174,a9176,a9178,a9180,a9182,a9184,a9186,a9188,a9190,a9192,
a9194,a9196,a9198,a9200,a9202,a9204,a9206,a9208,a9210,a9212,a9214,a9216,a9218,a9220,a9222,
a9224,a9226,a9228,a9230,a9232,a9234,a9236,a9238,a9240,a9242,a9244,a9246,a9248,a9250,a9252,
a9254,a9256,a9258,a9260,a9262,a9264,a9266,a9268,a9270,a9272,a9274,a9276,a9278,a9280,a9282,
a9284,a9286,a9288,a9290,a9292,a9294,a9296,a9298,a9300,a9302,a9304,a9306,a9308,a9310,a9312,
a9314,a9316,a9318,a9320,a9322,a9324,a9326,a9328,a9330,a9332,a9334,a9336,a9338,a9340,a9342,
a9344,a9346,a9348,a9350,a9352,a9354,a9356,a9358,a9360,a9362,a9364,a9366,a9368,a9370,a9372,
a9374,a9376,a9378,a9380,a9382,a9384,a9386,a9388,a9390,a9392,a9394,a9396,a9398,a9400,a9402,
a9404,a9406,a9408,a9410,a9412,a9414,a9416,a9418,a9420,a9422,a9424,a9426,a9428,a9430,a9432,
a9434,a9436,a9438,a9440,a9442,a9444,a9446,a9448,a9450,a9452,a9454,a9456,a9458,a9460,a9462,
a9464,a9466,a9468,a9470,a9472,a9474,a9476,a9478,a9480,a9482,a9484,a9486,a9488,a9490,a9492,
a9494,a9496,a9498,a9500,a9502,a9504,a9506,a9508,a9510,a9512,a9514,a9516,a9518,a9520,a9522,
a9524,a9526,a9528,a9530,a9532,a9534,a9536,a9538,a9540,a9542,a9544,a9546,a9548,a9550,a9552,
a9554,a9556,a9558,a9560,a9562,a9564,a9566,a9568,a9570,a9572,a9574,a9576,a9578,a9580,a9582,
a9584,a9586,a9588,a9590,a9592,a9594,a9596,a9598,a9600,a9602,a9604,a9606,a9608,a9610,a9612,
a9614,a9616,a9618,a9620,a9622,a9624,a9626,a9628,a9630,a9632,a9634,a9636,a9638,a9640,a9642,
a9644,a9646,a9648,a9650,a9652,a9654,a9656,a9658,a9660,a9662,a9664,a9666,a9668,a9670,a9672,
a9674,a9676,a9678,a9680,a9682,a9684,a9686,a9688,a9690,a9692,a9694,a9696,a9698,a9700,a9702,
a9704,a9706,a9708,a9710,a9712,a9714,a9716,a9718,a9720,a9722,a9724,a9726,a9728,a9730,a9732,
a9734,a9736,a9738,a9740,a9742,a9744,a9746,a9748,a9750,a9752,a9754,a9756,a9758,a9760,a9762,
a9764,a9766,a9768,a9770,a9772,a9774,a9776,a9778,a9780,a9782,a9784,a9786,a9788,a9790,a9792,
a9794,a9796,a9798,a9800,a9802,a9804,a9806,a9808,a9810,a9812,a9814,a9816,a9818,a9820,a9822,
a9824,a9826,a9828,a9830,a9832,a9834,a9836,a9838,a9840,a9842,a9844,a9846,a9848,a9850,a9852,
a9854,a9856,a9858,a9860,a9862,a9864,a9866,a9868,a9870,a9872,a9874,a9876,a9878,a9880,a9882,
a9884,a9886,a9888,a9890,a9892,a9894,a9896,a9898,a9900,a9902,a9904,a9906,a9908,a9910,a9912,
a9914,a9916,a9918,a9920,a9922,a9924,a9926,a9928,a9930,a9932,a9934,a9936,a9938,a9940,a9942,
a9944,a9946,a9948,a9950,a9952,a9954,a9956,a9958,a9960,a9962,a9964,a9966,a9968,a9970,a9972,
a9974,a9976,a9978,a9980,a9982,a9984,a9986,a9988,a9990,a9992,a9994,a9996,a9998,a10000,a10002,
a10004,a10006,a10008,a10010,a10012,a10014,a10016,a10018,a10020,a10022,a10024,a10026,a10028,a10030,a10032,
a10034,a10036,a10038,a10040,a10042,a10044,a10046,a10048,a10050,a10052,a10054,a10056,a10058,a10060,a10062,
a10064,a10066,a10068,a10070,a10072,a10074,a10076,a10078,a10080,a10082,a10084,a10086,a10088,a10090,a10092,
a10094,a10096,a10098,a10100,a10102,a10104,a10106,a10108,a10110,a10112,a10114,a10116,a10118,a10120,a10122,
a10124,a10126,a10128,a10130,a10132,a10134,a10136,a10138,a10140,a10142,a10144,a10146,a10148,a10150,a10152,
a10154,a10156,a10158,a10160,a10162,a10164,a10166,a10168,a10170,a10172,a10174,a10176,a10178,a10180,a10182,
a10184,a10186,a10188,a10190,a10192,a10194,a10196,a10198,a10200,a10202,a10204,a10206,a10208,a10210,a10212,
a10214,a10216,a10218,a10220,a10222,a10224,a10226,a10228,a10230,a10232,a10234,a10236,a10238,a10240,a10242,
a10244,a10246,a10248,a10250,a10252,a10254,a10256,a10258,a10260,a10262,a10264,a10266,a10268,a10270,a10272,
a10274,a10276,a10278,a10280,a10282,a10284,a10286,a10288,a10290,a10292,a10294,a10296,a10298,a10300,a10302,
a10304,a10306,a10308,a10310,a10312,a10314,a10316,a10318,a10320,a10322,a10324,a10326,a10328,a10330,a10332,
a10334,a10336,a10338,a10340,a10342,a10344,a10346,a10348,a10350,a10352,a10354,a10356,a10358,a10360,a10362,
a10364,a10366,a10368,a10370,a10372,a10374,a10376,a10378,a10380,a10382,a10384,a10386,a10388,a10390,a10392,
a10394,a10396,a10398,a10400,a10402,a10404,a10406,a10408,a10410,a10412,a10414,a10416,a10418,a10420,a10422,
a10424,a10426,a10428,a10430,a10432,a10434,a10436,a10438,a10440,a10442,a10444,a10446,a10448,a10450,a10452,
a10454,a10456,a10458,a10460,a10462,a10464,a10466,a10468,a10470,a10472,a10474,a10476,a10478,a10480,a10482,
a10484,a10486,a10488,a10490,a10492,a10494,a10496,a10498,a10500,a10502,a10504,a10506,a10508,a10510,a10512,
a10514,a10516,a10518,a10520,a10522,a10524,a10526,a10528,a10530,a10532,a10534,a10536,a10538,a10540,a10542,
a10544,a10546,a10548,a10550,a10552,a10554,a10556,a10558,a10560,a10562,a10564,a10566,a10568,a10570,a10572,
a10574,a10576,a10578,a10580,a10582,a10584,a10586,a10588,a10590,a10592,a10594,a10596,a10598,a10600,a10602,
a10604,a10606,a10608,a10610,a10612,a10614,a10616,a10618,a10620,a10622,a10624,a10626,a10628,a10630,a10632,
a10634,a10636,a10638,a10640,a10642,a10644,a10646,a10648,a10650,a10652,a10654,a10656,a10658,a10660,a10662,
a10664,a10666,a10668,a10670,a10672,a10674,a10676,a10678,a10680,a10682,a10684,a10686,a10688,a10690,a10692,
a10694,a10696,a10698,a10700,a10702,a10704,a10706,a10708,a10710,a10712,a10714,a10716,a10718,a10720,a10722,
a10724,a10726,a10728,a10730,a10732,a10734,a10736,a10738,a10740,a10742,a10744,a10746,a10748,a10750,a10752,
a10754,a10756,a10758,a10760,a10762,a10764,a10766,a10768,a10770,a10772,a10774,a10776,a10778,a10780,a10782,
a10784,a10786,a10788,a10790,a10792,a10794,a10796,a10798,a10800,a10802,a10804,a10806,a10808,a10810,a10812,
a10814,a10816,a10818,a10820,a10822,a10824,a10826,a10828,a10830,a10832,a10834,a10836,a10838,a10840,a10842,
a10844,a10846,a10848,a10850,a10852,a10854,a10856,a10858,a10860,a10862,a10864,a10866,a10868,a10870,a10872,
a10874,a10876,a10878,a10880,a10882,a10884,a10886,a10888,a10890,a10892,a10894,a10896,a10898,a10900,a10902,
a10904,a10906,a10908,a10910,a10912,a10914,a10916,a10918,a10920,a10922,a10924,a10926,a10928,a10930,a10932,
a10934,a10936,a10938,a10940,a10942,a10944,a10946,a10948,a10950,a10952,a10954,a10956,a10958,a10960,a10962,
a10964,a10966,a10968,a10970,a10972,a10974,a10976,a10978,a10980,a10982,a10984,a10986,a10988,a10990,a10992,
a10994,a10996,a10998,a11000,a11002,a11004,a11006,a11008,a11010,a11012,a11014,a11016,a11018,a11020,a11022,
a11024,a11026,a11028,a11030,a11032,a11034,a11036,a11038,a11040,a11042,a11044,a11046,a11048,a11050,a11052,
a11054,a11056,a11058,a11060,a11062,a11064,a11066,a11068,a11070,a11072,a11074,a11076,a11078,a11080,a11082,
a11084,a11086,a11088,a11090,a11092,a11094,a11096,a11098,a11100,a11102,a11104,a11106,a11108,a11110,a11112,
a11114,a11116,a11118,a11120,a11122,a11124,a11126,a11128,a11130,a11132,a11134,a11136,a11138,a11140,a11142,
a11144,a11146,a11148,a11150,a11152,a11154,a11156,a11158,a11160,a11162,a11164,a11166,a11168,a11170,a11172,
a11174,a11176,a11178,a11180,a11182,a11184,a11186,a11188,a11190,a11192,a11194,a11196,a11198,a11200,a11202,
a11204,a11206,a11208,a11210,a11212,a11214,a11216,a11218,a11220,a11222,a11224,a11226,a11228,a11230,a11232,
a11234,a11236,a11238,a11240,a11242,a11244,a11246,a11248,a11250,a11252,a11254,a11256,a11258,a11260,a11262,
a11264,a11266,a11268,a11270,a11272,a11274,a11276,a11278,a11280,a11282,a11284,a11286,a11288,a11290,a11292,
a11294,a11296,a11298,a11300,a11302,a11304,a11306,a11308,a11310,a11312,a11314,a11316,a11318,a11320,a11322,
a11324,a11326,a11328,a11330,a11332,a11334,a11336,a11338,a11340,a11342,a11344,a11346,a11348,a11350,a11352,
a11354,a11356,a11358,a11360,a11362,a11364,a11366,a11368,a11370,a11372,a11374,a11376,a11378,a11380,a11382,
a11384,a11386,a11388,a11390,a11392,a11394,a11396,a11398,a11400,a11402,a11404,a11406,a11408,a11410,a11412,
a11414,a11416,a11418,a11420,a11422,a11424,a11426,a11428,a11430,a11432,a11434,a11436,a11438,a11440,a11442,
a11444,a11446,a11448,a11450,a11452,a11454,a11456,a11458,a11460,a11462,a11464,a11466,a11468,a11470,a11472,
a11474,a11476,a11478,a11480,a11482,a11484,a11486,a11488,a11490,a11492,a11494,a11496,a11498,a11500,a11502,
a11504,a11506,a11508,a11510,a11512,a11514,a11516,a11518,a11520,a11522,a11524,a11526,a11528,a11530,a11532,
a11534,a11536,a11538,a11540,a11542,a11544,a11546,a11548,a11550,a11552,a11554,a11556,a11558,a11560,a11562,
a11564,a11566,a11568,a11570,a11572,a11574,a11576,a11578,a11580,a11582,a11584,a11586,a11588,a11590,a11592,
a11594,a11596,a11598,a11600,a11602,a11604,a11606,a11608,a11610,a11612,a11614,a11616,a11618,a11620,a11622,
a11624,a11626,a11628,a11630,a11632,a11634,a11636,a11638,a11640,a11642,a11644,a11646,a11648,a11650,a11652,
a11654,a11656,a11658,a11660,a11662,a11664,a11666,a11668,a11670,a11672,a11674,a11676,a11678,a11680,a11682,
a11684,a11686,a11688,a11690,a11692,a11694,a11696,a11698,a11700,a11702,a11704,a11706,a11708,a11710,a11712,
a11714,a11716,a11718,a11720,a11722,a11724,a11726,a11728,a11730,a11732,a11734,a11736,a11738,a11740,a11742,
a11744,a11746,a11748,a11750,a11752,a11754,a11756,a11758,a11760,a11762,a11764,a11766,a11768,a11770,a11772,
a11774,a11776,a11778,a11780,a11782,a11784,a11786,a11788,a11790,a11792,a11794,a11796,a11798,a11800,a11802,
a11804,a11806,a11808,a11810,a11812,a11814,a11816,a11818,a11820,a11822,a11824,a11826,a11828,a11830,a11832,
a11834,a11836,a11838,a11840,a11842,a11844,a11846,a11848,a11850,a11852,a11854,a11856,a11858,a11860,a11862,
a11864,a11866,a11868,a11870,a11872,a11874,a11876,a11878,a11880,a11882,a11884,a11886,a11888,a11890,a11892,
a11894,a11896,a11898,a11900,a11902,a11904,a11906,a11908,a11910,a11912,a11914,a11916,a11918,a11920,a11922,
a11924,a11926,a11928,a11930,a11932,a11934,a11936,a11938,a11942,p0;

reg l476,l478,l480,l482,l484,l486,l488,l490,l492,l494,l496,l498,l500,l502,l504,
l506,l508,l510,l512,l514,l516,l518,l520,l522,l524,l526,l528,l530,l532,l534,
l536,l538,l540,l542,l544,l546,l548,l550,l552,l554,l556,l558,l560,l562,l564,
l566,l568,l570,l572,l574,l576,l578,l580,l582,l584,l586,l588,l590,l592,l594,
l596,l598,l600,l602,l604,l606,l608,l610,l612,l614,l616,l618,l620,l622,l624,
l626,l628,l630,l632,l634,l636,l638,l640,l642,l644,l646,l648,l650,l652,l654,
l656,l658,l660,l662,l664,l666,l668,l670,l672,l674,l676,l678,l680,l682,l684,
l686,l688,l690,l692,l694,l696,l698,l700,l702,l704,l706,l708,l710,l712,l714,
l716,l718,l720,l722,l724,l726,l728,l730,l732,l734,l736,l738,l740,l742,l744,
l746,l748,l750,l752,l754,l756,l758,l760,l762,l764,l766,l768,l770,l772,l774,
l776,l778,l780,l782,l784,l786,l788,l790,l792,l794,l796,l798,l800,l802,l804,
l806,l808,l810,l812,l814,l816,l818,l820,l822,l824,l826,l828,l830,l832,l834,
l836,l838,l840,l842,l844,l846,l848,l850,l852,l854,l856,l858,l860,l862,l864,
l866,l868,l870,l872,l874,l876,l878,l880,l882,l884,l886,l888,l890,l892,l894,
l896,l898,l900,l902,l904,l906,l908,l910,l912,l914,l916,l918,l920,l922,l924,
l926,l928,l930,l932,l934,l936,l938,l940,l942,l944,l946,l948,l950,l952,l954,
l956,l958,l960,l962,l964,l966,l968,l970,l972,l974,l976,l978,l980,l982,l984,
l986,l988,l990,l992,l994,l996,l998,l1000,l1002,l1004,l1006,l1008,l1010,l1012,l1014,
l1016,l1018,l1020,l1022,l1024,l1026,l1028,l1030,l1032,l1034,l1036,l1038,l1040,l1042,l1044,
l1046,l1048,l1050,l1052,l1054,l1056,l1058,l1060,l1062,l1064,l1066,l1068,l1070,l1072,l1074,
l1076,l1078,l1080,l1082,l1084,l1086,l1088,l1090,l1092,l1094,l1096;

initial
begin
   l476 = 0;
   l478 = 0;
   l480 = 0;
   l482 = 0;
   l484 = 0;
   l486 = 0;
   l488 = 0;
   l490 = 0;
   l492 = 0;
   l494 = 0;
   l496 = 0;
   l498 = 0;
   l500 = 0;
   l502 = 0;
   l504 = 0;
   l506 = 0;
   l508 = 0;
   l510 = 0;
   l512 = 0;
   l514 = 0;
   l516 = 0;
   l518 = 0;
   l520 = 0;
   l522 = 0;
   l524 = 0;
   l526 = 0;
   l528 = 0;
   l530 = 0;
   l532 = 0;
   l534 = 0;
   l536 = 0;
   l538 = 0;
   l540 = 0;
   l542 = 0;
   l544 = 0;
   l546 = 0;
   l548 = 0;
   l550 = 0;
   l552 = 0;
   l554 = 0;
   l556 = 0;
   l558 = 0;
   l560 = 0;
   l562 = 0;
   l564 = 0;
   l566 = 0;
   l568 = 0;
   l570 = 0;
   l572 = 0;
   l574 = 0;
   l576 = 0;
   l578 = 0;
   l580 = 0;
   l582 = 0;
   l584 = 0;
   l586 = 0;
   l588 = 0;
   l590 = 0;
   l592 = 0;
   l594 = 0;
   l596 = 0;
   l598 = 0;
   l600 = 0;
   l602 = 0;
   l604 = 0;
   l606 = 0;
   l608 = 0;
   l610 = 0;
   l612 = 0;
   l614 = 0;
   l616 = 0;
   l618 = 0;
   l620 = 0;
   l622 = 0;
   l624 = 0;
   l626 = 0;
   l628 = 0;
   l630 = 0;
   l632 = 0;
   l634 = 0;
   l636 = 0;
   l638 = 0;
   l640 = 0;
   l642 = 0;
   l644 = 0;
   l646 = 0;
   l648 = 0;
   l650 = 0;
   l652 = 0;
   l654 = 0;
   l656 = 0;
   l658 = 0;
   l660 = 0;
   l662 = 0;
   l664 = 0;
   l666 = 0;
   l668 = 0;
   l670 = 0;
   l672 = 0;
   l674 = 0;
   l676 = 0;
   l678 = 0;
   l680 = 0;
   l682 = 0;
   l684 = 0;
   l686 = 0;
   l688 = 0;
   l690 = 0;
   l692 = 0;
   l694 = 0;
   l696 = 0;
   l698 = 0;
   l700 = 0;
   l702 = 0;
   l704 = 0;
   l706 = 0;
   l708 = 0;
   l710 = 0;
   l712 = 0;
   l714 = 0;
   l716 = 0;
   l718 = 0;
   l720 = 0;
   l722 = 0;
   l724 = 0;
   l726 = 0;
   l728 = 0;
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
   l802 = 0;
   l804 = 0;
   l806 = 0;
   l808 = 0;
   l810 = 0;
   l812 = 0;
   l814 = 0;
   l816 = 0;
   l818 = 0;
   l820 = 0;
   l822 = 0;
   l824 = 0;
   l826 = 0;
   l828 = 0;
   l830 = 0;
   l832 = 0;
   l834 = 0;
   l836 = 0;
   l838 = 0;
   l840 = 0;
   l842 = 0;
   l844 = 0;
   l846 = 0;
   l848 = 0;
   l850 = 0;
   l852 = 0;
   l854 = 0;
   l856 = 0;
   l858 = 0;
   l860 = 0;
   l862 = 0;
   l864 = 0;
   l866 = 0;
   l868 = 0;
   l870 = 0;
   l872 = 0;
   l874 = 0;
   l876 = 0;
   l878 = 0;
   l880 = 0;
   l882 = 0;
   l884 = 0;
   l886 = 0;
   l888 = 0;
   l890 = 0;
   l892 = 0;
   l894 = 0;
   l896 = 0;
   l898 = 0;
   l900 = 0;
   l902 = 0;
   l904 = 0;
   l906 = 0;
   l908 = 0;
   l910 = 0;
   l912 = 0;
   l914 = 0;
   l916 = 0;
   l918 = 0;
   l920 = 0;
   l922 = 0;
   l924 = 0;
   l926 = 0;
   l928 = 0;
   l930 = 0;
   l932 = 0;
   l934 = 0;
   l936 = 0;
   l938 = 0;
   l940 = 0;
   l942 = 0;
   l944 = 0;
   l946 = 0;
   l948 = 0;
   l950 = 0;
   l952 = 0;
   l954 = 0;
   l956 = 0;
   l958 = 0;
   l960 = 0;
   l962 = 0;
   l964 = 0;
   l966 = 0;
   l968 = 0;
   l970 = 0;
   l972 = 0;
   l974 = 0;
   l976 = 0;
   l978 = 0;
   l980 = 0;
   l982 = 0;
   l984 = 0;
   l986 = 0;
   l988 = 0;
   l990 = 0;
   l992 = 0;
   l994 = 0;
   l996 = 0;
   l998 = 0;
   l1000 = 0;
   l1002 = 0;
   l1004 = 0;
   l1006 = 0;
   l1008 = 0;
   l1010 = 0;
   l1012 = 0;
   l1014 = 0;
   l1016 = 0;
   l1018 = 0;
   l1020 = 0;
   l1022 = 0;
   l1024 = 0;
   l1026 = 0;
   l1028 = 0;
   l1030 = 0;
   l1032 = 0;
   l1034 = 0;
   l1036 = 0;
   l1038 = 0;
   l1040 = 0;
   l1042 = 0;
   l1044 = 0;
   l1046 = 0;
   l1048 = 0;
   l1050 = 0;
   l1052 = 0;
   l1054 = 0;
   l1056 = 0;
   l1058 = 0;
   l1060 = 0;
   l1062 = 0;
   l1064 = 0;
   l1066 = 0;
   l1068 = 0;
   l1070 = 0;
   l1072 = 0;
   l1074 = 0;
   l1076 = 0;
   l1078 = 0;
   l1080 = 0;
   l1082 = 0;
   l1084 = 0;
   l1086 = 0;
   l1088 = 0;
   l1090 = 0;
   l1092 = 0;
   l1094 = 0;
   l1096 = 0;
end

always @(posedge i2)
   l476 <= i2;

always @(posedge i4)
   l478 <= i4;

always @(posedge i6)
   l480 <= i6;

always @(posedge i8)
   l482 <= i8;

always @(posedge i10)
   l484 <= i10;

always @(posedge i12)
   l486 <= i12;

always @(posedge i14)
   l488 <= i14;

always @(posedge i16)
   l490 <= i16;

always @(posedge i18)
   l492 <= i18;

always @(posedge i20)
   l494 <= i20;

always @(posedge i22)
   l496 <= i22;

always @(posedge i24)
   l498 <= i24;

always @(posedge i26)
   l500 <= i26;

always @(posedge i28)
   l502 <= i28;

always @(posedge i30)
   l504 <= i30;

always @(posedge i32)
   l506 <= i32;

always @(posedge i34)
   l508 <= i34;

always @(posedge i36)
   l510 <= i36;

always @(posedge i38)
   l512 <= i38;

always @(posedge i40)
   l514 <= i40;

always @(posedge i42)
   l516 <= i42;

always @(posedge i44)
   l518 <= i44;

always @(posedge i46)
   l520 <= i46;

always @(posedge i48)
   l522 <= i48;

always @(posedge i50)
   l524 <= i50;

always @(posedge i52)
   l526 <= i52;

always @(posedge i54)
   l528 <= i54;

always @(posedge i56)
   l530 <= i56;

always @(posedge i58)
   l532 <= i58;

always @(posedge i60)
   l534 <= i60;

always @(posedge i62)
   l536 <= i62;

always @(posedge i64)
   l538 <= i64;

always @(posedge i66)
   l540 <= i66;

always @(posedge i68)
   l542 <= i68;

always @(posedge i70)
   l544 <= i70;

always @(posedge i72)
   l546 <= i72;

always @(posedge i74)
   l548 <= i74;

always @(posedge i76)
   l550 <= i76;

always @(posedge i78)
   l552 <= i78;

always @(posedge i80)
   l554 <= i80;

always @(posedge i82)
   l556 <= i82;

always @(posedge i84)
   l558 <= i84;

always @(posedge i86)
   l560 <= i86;

always @(posedge i88)
   l562 <= i88;

always @(posedge i90)
   l564 <= i90;

always @(posedge i92)
   l566 <= i92;

always @(posedge i94)
   l568 <= i94;

always @(posedge i96)
   l570 <= i96;

always @(posedge i98)
   l572 <= i98;

always @(posedge i100)
   l574 <= i100;

always @(posedge i102)
   l576 <= i102;

always @(posedge i104)
   l578 <= i104;

always @(posedge i106)
   l580 <= i106;

always @(posedge i108)
   l582 <= i108;

always @(posedge i110)
   l584 <= i110;

always @(posedge i112)
   l586 <= i112;

always @(posedge i114)
   l588 <= i114;

always @(posedge i116)
   l590 <= i116;

always @(posedge i118)
   l592 <= i118;

always @(posedge i120)
   l594 <= i120;

always @(posedge i122)
   l596 <= i122;

always @(posedge i124)
   l598 <= i124;

always @(posedge a1154)
   l600 <= a1154;

always @(posedge a1170)
   l602 <= a1170;

always @(posedge i126)
   l604 <= i126;

always @(posedge i128)
   l606 <= i128;

always @(posedge a1198)
   l608 <= a1198;

always @(posedge i130)
   l610 <= i130;

always @(posedge i132)
   l612 <= i132;

always @(posedge a1242)
   l614 <= a1242;

always @(posedge a1258)
   l616 <= a1258;

always @(posedge i134)
   l618 <= i134;

always @(posedge i136)
   l620 <= i136;

always @(posedge a1278)
   l622 <= a1278;

always @(posedge i138)
   l624 <= i138;

always @(posedge i140)
   l626 <= i140;

always @(posedge a1322)
   l628 <= a1322;

always @(posedge a1338)
   l630 <= a1338;

always @(posedge i142)
   l632 <= i142;

always @(posedge i144)
   l634 <= i144;

always @(posedge a1358)
   l636 <= a1358;

always @(posedge a1442)
   l638 <= a1442;

always @(posedge a1466)
   l640 <= a1466;

always @(posedge a1492)
   l642 <= a1492;

always @(posedge i146)
   l644 <= i146;

always @(posedge i148)
   l646 <= i148;

always @(posedge i150)
   l648 <= i150;

always @(posedge i152)
   l650 <= i152;

always @(posedge i154)
   l652 <= i154;

always @(posedge a1504)
   l654 <= a1504;

always @(posedge a1658)
   l656 <= a1658;

always @(posedge a1668)
   l658 <= a1668;

always @(posedge a1678)
   l660 <= a1678;

always @(posedge a1688)
   l662 <= a1688;

always @(posedge i156)
   l664 <= i156;

always @(posedge i158)
   l666 <= i158;

always @(posedge a1746)
   l668 <= a1746;

always @(posedge a1762)
   l670 <= a1762;

always @(posedge i160)
   l672 <= i160;

always @(posedge i162)
   l674 <= i162;

always @(posedge a1790)
   l676 <= a1790;

always @(posedge i164)
   l678 <= i164;

always @(posedge i166)
   l680 <= i166;

always @(posedge a1834)
   l682 <= a1834;

always @(posedge a1850)
   l684 <= a1850;

always @(posedge i168)
   l686 <= i168;

always @(posedge i170)
   l688 <= i170;

always @(posedge a1870)
   l690 <= a1870;

always @(posedge i172)
   l692 <= i172;

always @(posedge i174)
   l694 <= i174;

always @(posedge a1914)
   l696 <= a1914;

always @(posedge a1930)
   l698 <= a1930;

always @(posedge i176)
   l700 <= i176;

always @(posedge i178)
   l702 <= i178;

always @(posedge a1950)
   l704 <= a1950;

always @(posedge a2034)
   l706 <= a2034;

always @(posedge a2058)
   l708 <= a2058;

always @(posedge a2084)
   l710 <= a2084;

always @(posedge i180)
   l712 <= i180;

always @(posedge i182)
   l714 <= i182;

always @(posedge i184)
   l716 <= i184;

always @(posedge i186)
   l718 <= i186;

always @(posedge i188)
   l720 <= i188;

always @(posedge a2096)
   l722 <= a2096;

always @(posedge a2250)
   l724 <= a2250;

always @(posedge a2260)
   l726 <= a2260;

always @(posedge a2270)
   l728 <= a2270;

always @(posedge a2280)
   l730 <= a2280;

always @(posedge i190)
   l732 <= i190;

always @(posedge i192)
   l734 <= i192;

always @(posedge a2338)
   l736 <= a2338;

always @(posedge a2354)
   l738 <= a2354;

always @(posedge i194)
   l740 <= i194;

always @(posedge i196)
   l742 <= i196;

always @(posedge a2382)
   l744 <= a2382;

always @(posedge i198)
   l746 <= i198;

always @(posedge i200)
   l748 <= i200;

always @(posedge a2426)
   l750 <= a2426;

always @(posedge a2442)
   l752 <= a2442;

always @(posedge i202)
   l754 <= i202;

always @(posedge i204)
   l756 <= i204;

always @(posedge a2462)
   l758 <= a2462;

always @(posedge i206)
   l760 <= i206;

always @(posedge i208)
   l762 <= i208;

always @(posedge a2506)
   l764 <= a2506;

always @(posedge a2522)
   l766 <= a2522;

always @(posedge i210)
   l768 <= i210;

always @(posedge i212)
   l770 <= i212;

always @(posedge a2542)
   l772 <= a2542;

always @(posedge a2626)
   l774 <= a2626;

always @(posedge a2650)
   l776 <= a2650;

always @(posedge a2676)
   l778 <= a2676;

always @(posedge i214)
   l780 <= i214;

always @(posedge i216)
   l782 <= i216;

always @(posedge i218)
   l784 <= i218;

always @(posedge i220)
   l786 <= i220;

always @(posedge i222)
   l788 <= i222;

always @(posedge a2688)
   l790 <= a2688;

always @(posedge a2842)
   l792 <= a2842;

always @(posedge a2852)
   l794 <= a2852;

always @(posedge a2862)
   l796 <= a2862;

always @(posedge a2872)
   l798 <= a2872;

always @(posedge i224)
   l800 <= i224;

always @(posedge i226)
   l802 <= i226;

always @(posedge a2930)
   l804 <= a2930;

always @(posedge a2946)
   l806 <= a2946;

always @(posedge i228)
   l808 <= i228;

always @(posedge i230)
   l810 <= i230;

always @(posedge a2974)
   l812 <= a2974;

always @(posedge i232)
   l814 <= i232;

always @(posedge i234)
   l816 <= i234;

always @(posedge a3018)
   l818 <= a3018;

always @(posedge a3034)
   l820 <= a3034;

always @(posedge i236)
   l822 <= i236;

always @(posedge i238)
   l824 <= i238;

always @(posedge a3054)
   l826 <= a3054;

always @(posedge i240)
   l828 <= i240;

always @(posedge i242)
   l830 <= i242;

always @(posedge a3098)
   l832 <= a3098;

always @(posedge a3114)
   l834 <= a3114;

always @(posedge i244)
   l836 <= i244;

always @(posedge i246)
   l838 <= i246;

always @(posedge a3134)
   l840 <= a3134;

always @(posedge a3218)
   l842 <= a3218;

always @(posedge a3242)
   l844 <= a3242;

always @(posedge a3268)
   l846 <= a3268;

always @(posedge i248)
   l848 <= i248;

always @(posedge i250)
   l850 <= i250;

always @(posedge i252)
   l852 <= i252;

always @(posedge i254)
   l854 <= i254;

always @(posedge i256)
   l856 <= i256;

always @(posedge a3280)
   l858 <= a3280;

always @(posedge a3434)
   l860 <= a3434;

always @(posedge a3444)
   l862 <= a3444;

always @(posedge a3454)
   l864 <= a3454;

always @(posedge a3464)
   l866 <= a3464;

always @(posedge i258)
   l868 <= i258;

always @(posedge a3470)
   l870 <= a3470;

always @(posedge i260)
   l872 <= i260;

always @(posedge i262)
   l874 <= i262;

always @(posedge i264)
   l876 <= i264;

always @(posedge i266)
   l878 <= i266;

always @(posedge i268)
   l880 <= i268;

always @(posedge i270)
   l882 <= i270;

always @(posedge i272)
   l884 <= i272;

always @(posedge i274)
   l886 <= i274;

always @(posedge i276)
   l888 <= i276;

always @(posedge i278)
   l890 <= i278;

always @(posedge i280)
   l892 <= i280;

always @(posedge i282)
   l894 <= i282;

always @(posedge i284)
   l896 <= i284;

always @(posedge i286)
   l898 <= i286;

always @(posedge i288)
   l900 <= i288;

always @(posedge i290)
   l902 <= i290;

always @(posedge i292)
   l904 <= i292;

always @(posedge i294)
   l906 <= i294;

always @(posedge i296)
   l908 <= i296;

always @(posedge i298)
   l910 <= i298;

always @(posedge i300)
   l912 <= i300;

always @(posedge i302)
   l914 <= i302;

always @(posedge i304)
   l916 <= i304;

always @(posedge i306)
   l918 <= i306;

always @(posedge i308)
   l920 <= i308;

always @(posedge i310)
   l922 <= i310;

always @(posedge i312)
   l924 <= i312;

always @(posedge i314)
   l926 <= i314;

always @(posedge i316)
   l928 <= i316;

always @(posedge i318)
   l930 <= i318;

always @(posedge i320)
   l932 <= i320;

always @(posedge i322)
   l934 <= i322;

always @(posedge i324)
   l936 <= i324;

always @(posedge i326)
   l938 <= i326;

always @(posedge i328)
   l940 <= i328;

always @(posedge i330)
   l942 <= i330;

always @(posedge i332)
   l944 <= i332;

always @(posedge i334)
   l946 <= i334;

always @(posedge i336)
   l948 <= i336;

always @(posedge i338)
   l950 <= i338;

always @(posedge i340)
   l952 <= i340;

always @(posedge i342)
   l954 <= i342;

always @(posedge i344)
   l956 <= i344;

always @(posedge i346)
   l958 <= i346;

always @(posedge i348)
   l960 <= i348;

always @(posedge i350)
   l962 <= i350;

always @(posedge i352)
   l964 <= i352;

always @(posedge i354)
   l966 <= i354;

always @(posedge i356)
   l968 <= i356;

always @(posedge i358)
   l970 <= i358;

always @(posedge i360)
   l972 <= i360;

always @(posedge i362)
   l974 <= i362;

always @(posedge i364)
   l976 <= i364;

always @(posedge i366)
   l978 <= i366;

always @(posedge i368)
   l980 <= i368;

always @(posedge i370)
   l982 <= i370;

always @(posedge i372)
   l984 <= i372;

always @(posedge i374)
   l986 <= i374;

always @(posedge i376)
   l988 <= i376;

always @(posedge i378)
   l990 <= i378;

always @(posedge i380)
   l992 <= i380;

always @(posedge i382)
   l994 <= i382;

always @(posedge i384)
   l996 <= i384;

always @(posedge i386)
   l998 <= i386;

always @(posedge i388)
   l1000 <= i388;

always @(posedge i390)
   l1002 <= i390;

always @(posedge i392)
   l1004 <= i392;

always @(posedge i394)
   l1006 <= i394;

always @(posedge i396)
   l1008 <= i396;

always @(posedge i398)
   l1010 <= i398;

always @(posedge i400)
   l1012 <= i400;

always @(posedge i402)
   l1014 <= i402;

always @(posedge i404)
   l1016 <= i404;

always @(posedge i406)
   l1018 <= i406;

always @(posedge i408)
   l1020 <= i408;

always @(posedge i410)
   l1022 <= i410;

always @(posedge i412)
   l1024 <= i412;

always @(posedge i414)
   l1026 <= i414;

always @(posedge i416)
   l1028 <= i416;

always @(posedge i418)
   l1030 <= i418;

always @(posedge i420)
   l1032 <= i420;

always @(posedge i422)
   l1034 <= i422;

always @(posedge i424)
   l1036 <= i424;

always @(posedge i426)
   l1038 <= i426;

always @(posedge i428)
   l1040 <= i428;

always @(posedge i430)
   l1042 <= i430;

always @(posedge i432)
   l1044 <= i432;

always @(posedge i434)
   l1046 <= i434;

always @(posedge i436)
   l1048 <= i436;

always @(posedge i438)
   l1050 <= i438;

always @(posedge i440)
   l1052 <= i440;

always @(posedge i442)
   l1054 <= i442;

always @(posedge i444)
   l1056 <= i444;

always @(posedge i446)
   l1058 <= i446;

always @(posedge i448)
   l1060 <= i448;

always @(posedge i450)
   l1062 <= i450;

always @(posedge i452)
   l1064 <= i452;

always @(posedge i454)
   l1066 <= i454;

always @(posedge i456)
   l1068 <= i456;

always @(posedge i458)
   l1070 <= i458;

always @(posedge i460)
   l1072 <= i460;

always @(posedge i462)
   l1074 <= i462;

always @(posedge a3478)
   l1076 <= a3478;

always @(posedge a3488)
   l1078 <= a3488;

always @(posedge a3496)
   l1080 <= a3496;

always @(posedge i464)
   l1082 <= i464;

always @(posedge a3498)
   l1084 <= a3498;

always @(posedge i468)
   l1086 <= i468;

always @(posedge i470)
   l1088 <= i470;

always @(posedge i472)
   l1090 <= i472;

always @(posedge i474)
   l1092 <= i474;

always @(posedge a11940)
   l1094 <= a11940;

always @(posedge c1)
   l1096 <= c1;


assign a1154 = a1152 & l1096;
assign a1170 = ~a1168 & l1096;
assign a1198 = ~a1196 & l1096;
assign a1242 = a1240 & l1096;
assign a1258 = ~a1256 & l1096;
assign a1278 = ~a1276 & l1096;
assign a1322 = a1320 & l1096;
assign a1338 = ~a1336 & l1096;
assign a1358 = ~a1356 & l1096;
assign a1442 = a1440 & l1096;
assign a1466 = ~a1464 & l1096;
assign a1492 = ~a1490 & l1096;
assign a1504 = ~a1502 & l1096;
assign a1658 = a1656 & l1096;
assign a1668 = a1666 & l1096;
assign a1678 = a1676 & l1096;
assign a1688 = a1686 & l1096;
assign a1746 = a1744 & l1096;
assign a1762 = ~a1760 & l1096;
assign a1790 = ~a1788 & l1096;
assign a1834 = a1832 & l1096;
assign a1850 = ~a1848 & l1096;
assign a1870 = ~a1868 & l1096;
assign a1914 = a1912 & l1096;
assign a1930 = ~a1928 & l1096;
assign a1950 = ~a1948 & l1096;
assign a2034 = a2032 & l1096;
assign a2058 = ~a2056 & l1096;
assign a2084 = ~a2082 & l1096;
assign a2096 = ~a2094 & l1096;
assign a2250 = a2248 & l1096;
assign a2260 = a2258 & l1096;
assign a2270 = a2268 & l1096;
assign a2280 = a2278 & l1096;
assign a2338 = a2336 & l1096;
assign a2354 = ~a2352 & l1096;
assign a2382 = ~a2380 & l1096;
assign a2426 = a2424 & l1096;
assign a2442 = ~a2440 & l1096;
assign a2462 = ~a2460 & l1096;
assign a2506 = a2504 & l1096;
assign a2522 = ~a2520 & l1096;
assign a2542 = ~a2540 & l1096;
assign a2626 = a2624 & l1096;
assign a2650 = ~a2648 & l1096;
assign a2676 = ~a2674 & l1096;
assign a2688 = ~a2686 & l1096;
assign a2842 = a2840 & l1096;
assign a2852 = a2850 & l1096;
assign a2862 = a2860 & l1096;
assign a2872 = a2870 & l1096;
assign a2930 = a2928 & l1096;
assign a2946 = ~a2944 & l1096;
assign a2974 = ~a2972 & l1096;
assign a3018 = a3016 & l1096;
assign a3034 = ~a3032 & l1096;
assign a3054 = ~a3052 & l1096;
assign a3098 = a3096 & l1096;
assign a3114 = ~a3112 & l1096;
assign a3134 = ~a3132 & l1096;
assign a3218 = a3216 & l1096;
assign a3242 = ~a3240 & l1096;
assign a3268 = ~a3266 & l1096;
assign a3280 = ~a3278 & l1096;
assign a3434 = a3432 & l1096;
assign a3444 = a3442 & l1096;
assign a3454 = a3452 & l1096;
assign a3464 = a3462 & l1096;
assign a3470 = ~a3468 & l1096;
assign a3478 = ~a3476 & l1096;
assign a3488 = ~a3486 & l1096;
assign a3496 = ~a3494 & l1096;
assign a3498 = ~a3472 & l1096;
assign a11940 = a11938 & l1096;
assign c1 = 1;
assign a1098 = l608 & ~l606;
assign a1100 = l642 & l640;
assign a1102 = a1100 & ~l638;
assign a1104 = a1102 & a1098;
assign a1106 = ~l608 & l606;
assign a1108 = a1106 & a1102;
assign a1110 = l642 & ~l640;
assign a1112 = a1110 & l638;
assign a1114 = a1112 & a1106;
assign a1116 = l598 & ~l596;
assign a1118 = a1100 & l638;
assign a1120 = a1118 & a1106;
assign a1122 = a1120 & a1116;
assign a1124 = ~l598 & ~l596;
assign a1126 = l608 & l606;
assign a1128 = a1110 & ~l638;
assign a1130 = a1128 & a1126;
assign a1132 = a1130 & a1124;
assign a1134 = a1128 & a1098;
assign a1136 = a1134 & a1116;
assign a1138 = a1128 & l644;
assign a1140 = ~a1138 & l600;
assign a1142 = a1140 & ~a1136;
assign a1144 = a1142 & ~a1132;
assign a1146 = ~a1144 & ~a1122;
assign a1148 = ~a1146 & ~a1114;
assign a1150 = ~a1148 & ~a1108;
assign a1152 = ~a1150 & ~a1104;
assign a1156 = ~a1138 & l602;
assign a1158 = a1156 & ~a1136;
assign a1160 = a1158 & ~a1132;
assign a1162 = ~a1160 & ~a1122;
assign a1164 = ~a1162 & ~a1114;
assign a1166 = ~a1164 & ~a1108;
assign a1168 = a1166 & ~a1104;
assign a1172 = ~l598 & l596;
assign a1174 = ~l642 & ~l640;
assign a1176 = a1174 & ~l638;
assign a1178 = a1176 & a1106;
assign a1180 = a1178 & a1172;
assign a1182 = ~l642 & l640;
assign a1184 = a1182 & ~l638;
assign a1186 = a1184 & a1106;
assign a1188 = a1186 & a1124;
assign a1190 = a1172 & a1120;
assign a1192 = ~a1190 & ~l608;
assign a1194 = a1192 & ~a1188;
assign a1196 = a1194 & ~a1180;
assign a1200 = l622 & ~l620;
assign a1202 = a1200 & a1102;
assign a1204 = ~l622 & l620;
assign a1206 = a1204 & a1102;
assign a1208 = a1204 & a1112;
assign a1210 = l612 & ~l610;
assign a1212 = a1204 & a1118;
assign a1214 = a1212 & a1210;
assign a1216 = ~l612 & ~l610;
assign a1218 = l622 & l620;
assign a1220 = a1218 & a1128;
assign a1222 = a1220 & a1216;
assign a1224 = a1200 & a1128;
assign a1226 = a1224 & a1210;
assign a1228 = ~a1138 & l614;
assign a1230 = a1228 & ~a1226;
assign a1232 = a1230 & ~a1222;
assign a1234 = ~a1232 & ~a1214;
assign a1236 = ~a1234 & ~a1208;
assign a1238 = ~a1236 & ~a1206;
assign a1240 = ~a1238 & ~a1202;
assign a1244 = ~a1138 & l616;
assign a1246 = a1244 & ~a1226;
assign a1248 = a1246 & ~a1222;
assign a1250 = ~a1248 & ~a1214;
assign a1252 = ~a1250 & ~a1208;
assign a1254 = ~a1252 & ~a1206;
assign a1256 = a1254 & ~a1202;
assign a1260 = ~l612 & l610;
assign a1262 = a1204 & a1176;
assign a1264 = a1262 & a1260;
assign a1266 = a1204 & a1184;
assign a1268 = a1266 & a1216;
assign a1270 = a1260 & a1212;
assign a1272 = ~a1270 & ~l622;
assign a1274 = a1272 & ~a1268;
assign a1276 = a1274 & ~a1264;
assign a1280 = l636 & ~l634;
assign a1282 = a1280 & a1102;
assign a1284 = ~l636 & l634;
assign a1286 = a1284 & a1102;
assign a1288 = a1284 & a1112;
assign a1290 = l626 & ~l624;
assign a1292 = a1284 & a1118;
assign a1294 = a1292 & a1290;
assign a1296 = ~l626 & ~l624;
assign a1298 = l636 & l634;
assign a1300 = a1298 & a1128;
assign a1302 = a1300 & a1296;
assign a1304 = a1280 & a1128;
assign a1306 = a1304 & a1290;
assign a1308 = ~a1138 & l628;
assign a1310 = a1308 & ~a1306;
assign a1312 = a1310 & ~a1302;
assign a1314 = ~a1312 & ~a1294;
assign a1316 = ~a1314 & ~a1288;
assign a1318 = ~a1316 & ~a1286;
assign a1320 = ~a1318 & ~a1282;
assign a1324 = ~a1138 & l630;
assign a1326 = a1324 & ~a1306;
assign a1328 = a1326 & ~a1302;
assign a1330 = ~a1328 & ~a1294;
assign a1332 = ~a1330 & ~a1288;
assign a1334 = ~a1332 & ~a1286;
assign a1336 = a1334 & ~a1282;
assign a1340 = ~l626 & l624;
assign a1342 = a1284 & a1176;
assign a1344 = a1342 & a1340;
assign a1346 = a1284 & a1184;
assign a1348 = a1346 & a1296;
assign a1350 = a1340 & a1292;
assign a1352 = ~a1350 & ~l636;
assign a1354 = a1352 & ~a1348;
assign a1356 = a1354 & ~a1344;
assign a1360 = ~l656 & l650;
assign a1362 = ~a1204 & ~a1106;
assign a1364 = a1204 & a1106;
assign a1366 = ~a1364 & ~a1284;
assign a1368 = ~a1366 & ~a1362;
assign a1370 = ~a1368 & a1176;
assign a1372 = a1370 & ~a1360;
assign a1374 = ~a1116 & a1098;
assign a1376 = ~a1374 & a1102;
assign a1378 = ~a1210 & a1200;
assign a1380 = ~a1378 & a1376;
assign a1382 = ~a1290 & a1280;
assign a1384 = ~a1382 & a1380;
assign a1386 = ~a1124 & a1106;
assign a1388 = ~a1386 & a1184;
assign a1390 = ~a1216 & a1204;
assign a1392 = ~a1390 & a1388;
assign a1394 = ~a1296 & a1284;
assign a1396 = ~a1394 & a1392;
assign a1398 = ~a1340 & a1284;
assign a1400 = ~a1260 & a1204;
assign a1402 = ~a1172 & a1106;
assign a1404 = ~a1402 & a1184;
assign a1406 = a1404 & ~a1400;
assign a1408 = a1406 & ~a1398;
assign a1410 = ~a1290 & a1284;
assign a1412 = ~a1116 & a1106;
assign a1414 = ~a1210 & a1204;
assign a1416 = ~a1414 & ~a1412;
assign a1418 = a1416 & ~a1410;
assign a1420 = ~a1402 & ~a1400;
assign a1422 = a1420 & ~a1398;
assign a1424 = ~a1422 & ~a1418;
assign a1426 = ~a1424 & ~a1110;
assign a1428 = a1426 & a1118;
assign a1430 = a1428 & ~a1174;
assign a1432 = ~a1430 & l638;
assign a1434 = ~a1432 & ~a1408;
assign a1436 = ~a1434 & ~a1396;
assign a1438 = a1436 & ~a1384;
assign a1440 = a1438 & ~a1372;
assign a1444 = a1112 & ~l652;
assign a1446 = a1174 & l638;
assign a1448 = l642 & l638;
assign a1450 = a1448 & l652;
assign a1452 = ~a1450 & a1446;
assign a1454 = ~a1452 & ~l640;
assign a1456 = a1454 & ~a1444;
assign a1458 = ~a1456 & ~a1408;
assign a1460 = a1458 & ~a1396;
assign a1462 = ~a1460 & ~a1384;
assign a1464 = a1462 & ~a1372;
assign a1468 = a1112 & l652;
assign a1470 = ~a1414 & ~a1410;
assign a1472 = a1470 & ~a1412;
assign a1474 = a1472 & a1118;
assign a1476 = ~a1474 & l642;
assign a1478 = ~a1476 & ~a1446;
assign a1480 = ~a1478 & ~a1468;
assign a1482 = ~a1480 & ~a1444;
assign a1484 = a1482 & ~a1408;
assign a1486 = a1484 & ~a1396;
assign a1488 = ~a1486 & ~a1384;
assign a1490 = ~a1488 & ~a1372;
assign a1494 = ~l662 & ~l660;
assign a1496 = ~a1494 & l658;
assign a1498 = a1496 & l656;
assign a1500 = a1498 & a1176;
assign a1502 = ~a1500 & ~l654;
assign a1506 = ~l660 & ~l658;
assign a1508 = a1506 & ~l656;
assign a1510 = l662 & ~l660;
assign a1512 = a1510 & ~l658;
assign a1514 = a1512 & ~l656;
assign a1516 = l660 & ~l658;
assign a1518 = a1516 & ~l656;
assign a1520 = l662 & l660;
assign a1522 = a1520 & ~l658;
assign a1524 = a1522 & ~l656;
assign a1526 = ~l660 & l658;
assign a1528 = a1526 & ~l656;
assign a1530 = a1510 & l658;
assign a1532 = a1530 & ~l656;
assign a1534 = l660 & l658;
assign a1536 = a1534 & ~l656;
assign a1538 = a1512 & l656;
assign a1540 = a1522 & l656;
assign a1542 = ~a1540 & a1526;
assign a1544 = ~a1542 & ~a1516;
assign a1546 = ~a1544 & ~a1538;
assign a1548 = ~a1546 & ~a1506;
assign a1550 = ~a1548 & l656;
assign a1552 = ~a1550 & ~a1536;
assign a1554 = ~a1552 & ~a1532;
assign a1556 = ~a1554 & ~a1528;
assign a1558 = ~a1556 & ~a1524;
assign a1560 = ~a1558 & ~a1518;
assign a1562 = ~a1560 & ~a1514;
assign a1564 = ~a1562 & ~a1508;
assign a1566 = ~a1564 & ~l662;
assign a1568 = a1494 & ~l658;
assign a1570 = a1568 & ~l656;
assign a1572 = l662 & ~l658;
assign a1574 = a1572 & ~l656;
assign a1576 = a1494 & l658;
assign a1578 = a1576 & ~l656;
assign a1580 = l662 & l658;
assign a1582 = a1580 & ~l656;
assign a1584 = a1568 & l656;
assign a1586 = ~l658 & l656;
assign a1588 = a1586 & ~a1510;
assign a1590 = a1588 & ~a1584;
assign a1592 = ~a1590 & ~a1582;
assign a1594 = ~l662 & l658;
assign a1596 = a1594 & ~l656;
assign a1598 = ~a1596 & a1592;
assign a1600 = ~a1598 & ~a1532;
assign a1602 = a1600 & ~a1578;
assign a1604 = ~a1602 & ~a1574;
assign a1606 = ~l662 & ~l658;
assign a1608 = a1606 & ~l656;
assign a1610 = ~a1608 & a1604;
assign a1612 = ~a1610 & l660;
assign a1614 = a1612 & ~a1514;
assign a1616 = a1614 & ~a1570;
assign a1618 = a1616 & a1566;
assign a1620 = ~l662 & l660;
assign a1622 = ~a1520 & ~l656;
assign a1624 = a1622 & ~a1620;
assign a1626 = a1510 & ~l656;
assign a1628 = ~a1626 & a1624;
assign a1630 = a1494 & ~l656;
assign a1632 = ~a1630 & a1628;
assign a1634 = ~a1632 & ~l658;
assign a1636 = ~a1634 & a1618;
assign a1638 = ~a1520 & ~l658;
assign a1640 = a1638 & ~a1620;
assign a1642 = a1640 & ~a1512;
assign a1644 = a1642 & ~a1568;
assign a1646 = ~a1644 & ~l656;
assign a1648 = ~a1646 & a1636;
assign a1650 = ~a1648 & l656;
assign a1652 = ~a1650 & a1176;
assign a1654 = ~a1176 & ~l656;
assign a1656 = ~a1654 & ~a1652;
assign a1660 = ~a1648 & l658;
assign a1662 = ~a1660 & a1176;
assign a1664 = ~a1176 & ~l658;
assign a1666 = ~a1664 & ~a1662;
assign a1670 = ~a1648 & l660;
assign a1672 = ~a1670 & a1176;
assign a1674 = ~a1176 & ~l660;
assign a1676 = ~a1674 & ~a1672;
assign a1680 = ~a1648 & ~l662;
assign a1682 = ~a1680 & a1176;
assign a1684 = ~a1176 & ~l662;
assign a1686 = ~a1684 & ~a1682;
assign a1690 = l676 & ~l674;
assign a1692 = l710 & l708;
assign a1694 = a1692 & ~l706;
assign a1696 = a1694 & a1690;
assign a1698 = ~l676 & l674;
assign a1700 = a1698 & a1694;
assign a1702 = l710 & ~l708;
assign a1704 = a1702 & l706;
assign a1706 = a1704 & a1698;
assign a1708 = l666 & ~l664;
assign a1710 = a1692 & l706;
assign a1712 = a1710 & a1698;
assign a1714 = a1712 & a1708;
assign a1716 = ~l666 & ~l664;
assign a1718 = l676 & l674;
assign a1720 = a1702 & ~l706;
assign a1722 = a1720 & a1718;
assign a1724 = a1722 & a1716;
assign a1726 = a1720 & a1690;
assign a1728 = a1726 & a1708;
assign a1730 = a1720 & l712;
assign a1732 = ~a1730 & l668;
assign a1734 = a1732 & ~a1728;
assign a1736 = a1734 & ~a1724;
assign a1738 = ~a1736 & ~a1714;
assign a1740 = ~a1738 & ~a1706;
assign a1742 = ~a1740 & ~a1700;
assign a1744 = ~a1742 & ~a1696;
assign a1748 = ~a1730 & l670;
assign a1750 = a1748 & ~a1728;
assign a1752 = a1750 & ~a1724;
assign a1754 = ~a1752 & ~a1714;
assign a1756 = ~a1754 & ~a1706;
assign a1758 = ~a1756 & ~a1700;
assign a1760 = a1758 & ~a1696;
assign a1764 = ~l666 & l664;
assign a1766 = ~l710 & ~l708;
assign a1768 = a1766 & ~l706;
assign a1770 = a1768 & a1698;
assign a1772 = a1770 & a1764;
assign a1774 = ~l710 & l708;
assign a1776 = a1774 & ~l706;
assign a1778 = a1776 & a1698;
assign a1780 = a1778 & a1716;
assign a1782 = a1764 & a1712;
assign a1784 = ~a1782 & ~l676;
assign a1786 = a1784 & ~a1780;
assign a1788 = a1786 & ~a1772;
assign a1792 = l690 & ~l688;
assign a1794 = a1792 & a1694;
assign a1796 = ~l690 & l688;
assign a1798 = a1796 & a1694;
assign a1800 = a1796 & a1704;
assign a1802 = l680 & ~l678;
assign a1804 = a1796 & a1710;
assign a1806 = a1804 & a1802;
assign a1808 = ~l680 & ~l678;
assign a1810 = l690 & l688;
assign a1812 = a1810 & a1720;
assign a1814 = a1812 & a1808;
assign a1816 = a1792 & a1720;
assign a1818 = a1816 & a1802;
assign a1820 = ~a1730 & l682;
assign a1822 = a1820 & ~a1818;
assign a1824 = a1822 & ~a1814;
assign a1826 = ~a1824 & ~a1806;
assign a1828 = ~a1826 & ~a1800;
assign a1830 = ~a1828 & ~a1798;
assign a1832 = ~a1830 & ~a1794;
assign a1836 = ~a1730 & l684;
assign a1838 = a1836 & ~a1818;
assign a1840 = a1838 & ~a1814;
assign a1842 = ~a1840 & ~a1806;
assign a1844 = ~a1842 & ~a1800;
assign a1846 = ~a1844 & ~a1798;
assign a1848 = a1846 & ~a1794;
assign a1852 = ~l680 & l678;
assign a1854 = a1796 & a1768;
assign a1856 = a1854 & a1852;
assign a1858 = a1796 & a1776;
assign a1860 = a1858 & a1808;
assign a1862 = a1852 & a1804;
assign a1864 = ~a1862 & ~l690;
assign a1866 = a1864 & ~a1860;
assign a1868 = a1866 & ~a1856;
assign a1872 = l704 & ~l702;
assign a1874 = a1872 & a1694;
assign a1876 = ~l704 & l702;
assign a1878 = a1876 & a1694;
assign a1880 = a1876 & a1704;
assign a1882 = l694 & ~l692;
assign a1884 = a1876 & a1710;
assign a1886 = a1884 & a1882;
assign a1888 = ~l694 & ~l692;
assign a1890 = l704 & l702;
assign a1892 = a1890 & a1720;
assign a1894 = a1892 & a1888;
assign a1896 = a1872 & a1720;
assign a1898 = a1896 & a1882;
assign a1900 = ~a1730 & l696;
assign a1902 = a1900 & ~a1898;
assign a1904 = a1902 & ~a1894;
assign a1906 = ~a1904 & ~a1886;
assign a1908 = ~a1906 & ~a1880;
assign a1910 = ~a1908 & ~a1878;
assign a1912 = ~a1910 & ~a1874;
assign a1916 = ~a1730 & l698;
assign a1918 = a1916 & ~a1898;
assign a1920 = a1918 & ~a1894;
assign a1922 = ~a1920 & ~a1886;
assign a1924 = ~a1922 & ~a1880;
assign a1926 = ~a1924 & ~a1878;
assign a1928 = a1926 & ~a1874;
assign a1932 = ~l694 & l692;
assign a1934 = a1876 & a1768;
assign a1936 = a1934 & a1932;
assign a1938 = a1876 & a1776;
assign a1940 = a1938 & a1888;
assign a1942 = a1932 & a1884;
assign a1944 = ~a1942 & ~l704;
assign a1946 = a1944 & ~a1940;
assign a1948 = a1946 & ~a1936;
assign a1952 = ~l724 & l718;
assign a1954 = ~a1796 & ~a1698;
assign a1956 = a1796 & a1698;
assign a1958 = ~a1956 & ~a1876;
assign a1960 = ~a1958 & ~a1954;
assign a1962 = ~a1960 & a1768;
assign a1964 = a1962 & ~a1952;
assign a1966 = ~a1708 & a1690;
assign a1968 = ~a1966 & a1694;
assign a1970 = ~a1802 & a1792;
assign a1972 = ~a1970 & a1968;
assign a1974 = ~a1882 & a1872;
assign a1976 = ~a1974 & a1972;
assign a1978 = ~a1716 & a1698;
assign a1980 = ~a1978 & a1776;
assign a1982 = ~a1808 & a1796;
assign a1984 = ~a1982 & a1980;
assign a1986 = ~a1888 & a1876;
assign a1988 = ~a1986 & a1984;
assign a1990 = ~a1932 & a1876;
assign a1992 = ~a1852 & a1796;
assign a1994 = ~a1764 & a1698;
assign a1996 = ~a1994 & a1776;
assign a1998 = a1996 & ~a1992;
assign a2000 = a1998 & ~a1990;
assign a2002 = ~a1882 & a1876;
assign a2004 = ~a1708 & a1698;
assign a2006 = ~a1802 & a1796;
assign a2008 = ~a2006 & ~a2004;
assign a2010 = a2008 & ~a2002;
assign a2012 = ~a1994 & ~a1992;
assign a2014 = a2012 & ~a1990;
assign a2016 = ~a2014 & ~a2010;
assign a2018 = ~a2016 & ~a1702;
assign a2020 = a2018 & a1710;
assign a2022 = a2020 & ~a1766;
assign a2024 = ~a2022 & l706;
assign a2026 = ~a2024 & ~a2000;
assign a2028 = ~a2026 & ~a1988;
assign a2030 = a2028 & ~a1976;
assign a2032 = a2030 & ~a1964;
assign a2036 = a1704 & ~l720;
assign a2038 = a1766 & l706;
assign a2040 = l710 & l706;
assign a2042 = a2040 & l720;
assign a2044 = ~a2042 & a2038;
assign a2046 = ~a2044 & ~l708;
assign a2048 = a2046 & ~a2036;
assign a2050 = ~a2048 & ~a2000;
assign a2052 = a2050 & ~a1988;
assign a2054 = ~a2052 & ~a1976;
assign a2056 = a2054 & ~a1964;
assign a2060 = a1704 & l720;
assign a2062 = ~a2006 & ~a2002;
assign a2064 = a2062 & ~a2004;
assign a2066 = a2064 & a1710;
assign a2068 = ~a2066 & l710;
assign a2070 = ~a2068 & ~a2038;
assign a2072 = ~a2070 & ~a2060;
assign a2074 = ~a2072 & ~a2036;
assign a2076 = a2074 & ~a2000;
assign a2078 = a2076 & ~a1988;
assign a2080 = ~a2078 & ~a1976;
assign a2082 = ~a2080 & ~a1964;
assign a2086 = ~l730 & ~l728;
assign a2088 = ~a2086 & l726;
assign a2090 = a2088 & l724;
assign a2092 = a2090 & a1768;
assign a2094 = ~a2092 & ~l722;
assign a2098 = ~l728 & ~l726;
assign a2100 = a2098 & ~l724;
assign a2102 = l730 & ~l728;
assign a2104 = a2102 & ~l726;
assign a2106 = a2104 & ~l724;
assign a2108 = l728 & ~l726;
assign a2110 = a2108 & ~l724;
assign a2112 = l730 & l728;
assign a2114 = a2112 & ~l726;
assign a2116 = a2114 & ~l724;
assign a2118 = ~l728 & l726;
assign a2120 = a2118 & ~l724;
assign a2122 = a2102 & l726;
assign a2124 = a2122 & ~l724;
assign a2126 = l728 & l726;
assign a2128 = a2126 & ~l724;
assign a2130 = a2104 & l724;
assign a2132 = a2114 & l724;
assign a2134 = ~a2132 & a2118;
assign a2136 = ~a2134 & ~a2108;
assign a2138 = ~a2136 & ~a2130;
assign a2140 = ~a2138 & ~a2098;
assign a2142 = ~a2140 & l724;
assign a2144 = ~a2142 & ~a2128;
assign a2146 = ~a2144 & ~a2124;
assign a2148 = ~a2146 & ~a2120;
assign a2150 = ~a2148 & ~a2116;
assign a2152 = ~a2150 & ~a2110;
assign a2154 = ~a2152 & ~a2106;
assign a2156 = ~a2154 & ~a2100;
assign a2158 = ~a2156 & ~l730;
assign a2160 = a2086 & ~l726;
assign a2162 = a2160 & ~l724;
assign a2164 = l730 & ~l726;
assign a2166 = a2164 & ~l724;
assign a2168 = a2086 & l726;
assign a2170 = a2168 & ~l724;
assign a2172 = l730 & l726;
assign a2174 = a2172 & ~l724;
assign a2176 = a2160 & l724;
assign a2178 = ~l726 & l724;
assign a2180 = a2178 & ~a2102;
assign a2182 = a2180 & ~a2176;
assign a2184 = ~a2182 & ~a2174;
assign a2186 = ~l730 & l726;
assign a2188 = a2186 & ~l724;
assign a2190 = ~a2188 & a2184;
assign a2192 = ~a2190 & ~a2124;
assign a2194 = a2192 & ~a2170;
assign a2196 = ~a2194 & ~a2166;
assign a2198 = ~l730 & ~l726;
assign a2200 = a2198 & ~l724;
assign a2202 = ~a2200 & a2196;
assign a2204 = ~a2202 & l728;
assign a2206 = a2204 & ~a2106;
assign a2208 = a2206 & ~a2162;
assign a2210 = a2208 & a2158;
assign a2212 = ~l730 & l728;
assign a2214 = ~a2112 & ~l724;
assign a2216 = a2214 & ~a2212;
assign a2218 = a2102 & ~l724;
assign a2220 = ~a2218 & a2216;
assign a2222 = a2086 & ~l724;
assign a2224 = ~a2222 & a2220;
assign a2226 = ~a2224 & ~l726;
assign a2228 = ~a2226 & a2210;
assign a2230 = ~a2112 & ~l726;
assign a2232 = a2230 & ~a2212;
assign a2234 = a2232 & ~a2104;
assign a2236 = a2234 & ~a2160;
assign a2238 = ~a2236 & ~l724;
assign a2240 = ~a2238 & a2228;
assign a2242 = ~a2240 & l724;
assign a2244 = ~a2242 & a1768;
assign a2246 = ~a1768 & ~l724;
assign a2248 = ~a2246 & ~a2244;
assign a2252 = ~a2240 & l726;
assign a2254 = ~a2252 & a1768;
assign a2256 = ~a1768 & ~l726;
assign a2258 = ~a2256 & ~a2254;
assign a2262 = ~a2240 & l728;
assign a2264 = ~a2262 & a1768;
assign a2266 = ~a1768 & ~l728;
assign a2268 = ~a2266 & ~a2264;
assign a2272 = ~a2240 & ~l730;
assign a2274 = ~a2272 & a1768;
assign a2276 = ~a1768 & ~l730;
assign a2278 = ~a2276 & ~a2274;
assign a2282 = l744 & ~l742;
assign a2284 = l778 & l776;
assign a2286 = a2284 & ~l774;
assign a2288 = a2286 & a2282;
assign a2290 = ~l744 & l742;
assign a2292 = a2290 & a2286;
assign a2294 = l778 & ~l776;
assign a2296 = a2294 & l774;
assign a2298 = a2296 & a2290;
assign a2300 = l734 & ~l732;
assign a2302 = a2284 & l774;
assign a2304 = a2302 & a2290;
assign a2306 = a2304 & a2300;
assign a2308 = ~l734 & ~l732;
assign a2310 = l744 & l742;
assign a2312 = a2294 & ~l774;
assign a2314 = a2312 & a2310;
assign a2316 = a2314 & a2308;
assign a2318 = a2312 & a2282;
assign a2320 = a2318 & a2300;
assign a2322 = a2312 & l780;
assign a2324 = ~a2322 & l736;
assign a2326 = a2324 & ~a2320;
assign a2328 = a2326 & ~a2316;
assign a2330 = ~a2328 & ~a2306;
assign a2332 = ~a2330 & ~a2298;
assign a2334 = ~a2332 & ~a2292;
assign a2336 = ~a2334 & ~a2288;
assign a2340 = ~a2322 & l738;
assign a2342 = a2340 & ~a2320;
assign a2344 = a2342 & ~a2316;
assign a2346 = ~a2344 & ~a2306;
assign a2348 = ~a2346 & ~a2298;
assign a2350 = ~a2348 & ~a2292;
assign a2352 = a2350 & ~a2288;
assign a2356 = ~l734 & l732;
assign a2358 = ~l778 & ~l776;
assign a2360 = a2358 & ~l774;
assign a2362 = a2360 & a2290;
assign a2364 = a2362 & a2356;
assign a2366 = ~l778 & l776;
assign a2368 = a2366 & ~l774;
assign a2370 = a2368 & a2290;
assign a2372 = a2370 & a2308;
assign a2374 = a2356 & a2304;
assign a2376 = ~a2374 & ~l744;
assign a2378 = a2376 & ~a2372;
assign a2380 = a2378 & ~a2364;
assign a2384 = l758 & ~l756;
assign a2386 = a2384 & a2286;
assign a2388 = ~l758 & l756;
assign a2390 = a2388 & a2286;
assign a2392 = a2388 & a2296;
assign a2394 = l748 & ~l746;
assign a2396 = a2388 & a2302;
assign a2398 = a2396 & a2394;
assign a2400 = ~l748 & ~l746;
assign a2402 = l758 & l756;
assign a2404 = a2402 & a2312;
assign a2406 = a2404 & a2400;
assign a2408 = a2384 & a2312;
assign a2410 = a2408 & a2394;
assign a2412 = ~a2322 & l750;
assign a2414 = a2412 & ~a2410;
assign a2416 = a2414 & ~a2406;
assign a2418 = ~a2416 & ~a2398;
assign a2420 = ~a2418 & ~a2392;
assign a2422 = ~a2420 & ~a2390;
assign a2424 = ~a2422 & ~a2386;
assign a2428 = ~a2322 & l752;
assign a2430 = a2428 & ~a2410;
assign a2432 = a2430 & ~a2406;
assign a2434 = ~a2432 & ~a2398;
assign a2436 = ~a2434 & ~a2392;
assign a2438 = ~a2436 & ~a2390;
assign a2440 = a2438 & ~a2386;
assign a2444 = ~l748 & l746;
assign a2446 = a2388 & a2360;
assign a2448 = a2446 & a2444;
assign a2450 = a2388 & a2368;
assign a2452 = a2450 & a2400;
assign a2454 = a2444 & a2396;
assign a2456 = ~a2454 & ~l758;
assign a2458 = a2456 & ~a2452;
assign a2460 = a2458 & ~a2448;
assign a2464 = l772 & ~l770;
assign a2466 = a2464 & a2286;
assign a2468 = ~l772 & l770;
assign a2470 = a2468 & a2286;
assign a2472 = a2468 & a2296;
assign a2474 = l762 & ~l760;
assign a2476 = a2468 & a2302;
assign a2478 = a2476 & a2474;
assign a2480 = ~l762 & ~l760;
assign a2482 = l772 & l770;
assign a2484 = a2482 & a2312;
assign a2486 = a2484 & a2480;
assign a2488 = a2464 & a2312;
assign a2490 = a2488 & a2474;
assign a2492 = ~a2322 & l764;
assign a2494 = a2492 & ~a2490;
assign a2496 = a2494 & ~a2486;
assign a2498 = ~a2496 & ~a2478;
assign a2500 = ~a2498 & ~a2472;
assign a2502 = ~a2500 & ~a2470;
assign a2504 = ~a2502 & ~a2466;
assign a2508 = ~a2322 & l766;
assign a2510 = a2508 & ~a2490;
assign a2512 = a2510 & ~a2486;
assign a2514 = ~a2512 & ~a2478;
assign a2516 = ~a2514 & ~a2472;
assign a2518 = ~a2516 & ~a2470;
assign a2520 = a2518 & ~a2466;
assign a2524 = ~l762 & l760;
assign a2526 = a2468 & a2360;
assign a2528 = a2526 & a2524;
assign a2530 = a2468 & a2368;
assign a2532 = a2530 & a2480;
assign a2534 = a2524 & a2476;
assign a2536 = ~a2534 & ~l772;
assign a2538 = a2536 & ~a2532;
assign a2540 = a2538 & ~a2528;
assign a2544 = ~l792 & l786;
assign a2546 = ~a2388 & ~a2290;
assign a2548 = a2388 & a2290;
assign a2550 = ~a2548 & ~a2468;
assign a2552 = ~a2550 & ~a2546;
assign a2554 = ~a2552 & a2360;
assign a2556 = a2554 & ~a2544;
assign a2558 = ~a2300 & a2282;
assign a2560 = ~a2558 & a2286;
assign a2562 = ~a2394 & a2384;
assign a2564 = ~a2562 & a2560;
assign a2566 = ~a2474 & a2464;
assign a2568 = ~a2566 & a2564;
assign a2570 = ~a2308 & a2290;
assign a2572 = ~a2570 & a2368;
assign a2574 = ~a2400 & a2388;
assign a2576 = ~a2574 & a2572;
assign a2578 = ~a2480 & a2468;
assign a2580 = ~a2578 & a2576;
assign a2582 = ~a2524 & a2468;
assign a2584 = ~a2444 & a2388;
assign a2586 = ~a2356 & a2290;
assign a2588 = ~a2586 & a2368;
assign a2590 = a2588 & ~a2584;
assign a2592 = a2590 & ~a2582;
assign a2594 = ~a2474 & a2468;
assign a2596 = ~a2300 & a2290;
assign a2598 = ~a2394 & a2388;
assign a2600 = ~a2598 & ~a2596;
assign a2602 = a2600 & ~a2594;
assign a2604 = ~a2586 & ~a2584;
assign a2606 = a2604 & ~a2582;
assign a2608 = ~a2606 & ~a2602;
assign a2610 = ~a2608 & ~a2294;
assign a2612 = a2610 & a2302;
assign a2614 = a2612 & ~a2358;
assign a2616 = ~a2614 & l774;
assign a2618 = ~a2616 & ~a2592;
assign a2620 = ~a2618 & ~a2580;
assign a2622 = a2620 & ~a2568;
assign a2624 = a2622 & ~a2556;
assign a2628 = a2296 & ~l788;
assign a2630 = a2358 & l774;
assign a2632 = l778 & l774;
assign a2634 = a2632 & l788;
assign a2636 = ~a2634 & a2630;
assign a2638 = ~a2636 & ~l776;
assign a2640 = a2638 & ~a2628;
assign a2642 = ~a2640 & ~a2592;
assign a2644 = a2642 & ~a2580;
assign a2646 = ~a2644 & ~a2568;
assign a2648 = a2646 & ~a2556;
assign a2652 = a2296 & l788;
assign a2654 = ~a2598 & ~a2594;
assign a2656 = a2654 & ~a2596;
assign a2658 = a2656 & a2302;
assign a2660 = ~a2658 & l778;
assign a2662 = ~a2660 & ~a2630;
assign a2664 = ~a2662 & ~a2652;
assign a2666 = ~a2664 & ~a2628;
assign a2668 = a2666 & ~a2592;
assign a2670 = a2668 & ~a2580;
assign a2672 = ~a2670 & ~a2568;
assign a2674 = ~a2672 & ~a2556;
assign a2678 = ~l798 & ~l796;
assign a2680 = ~a2678 & l794;
assign a2682 = a2680 & l792;
assign a2684 = a2682 & a2360;
assign a2686 = ~a2684 & ~l790;
assign a2690 = ~l796 & ~l794;
assign a2692 = a2690 & ~l792;
assign a2694 = l798 & ~l796;
assign a2696 = a2694 & ~l794;
assign a2698 = a2696 & ~l792;
assign a2700 = l796 & ~l794;
assign a2702 = a2700 & ~l792;
assign a2704 = l798 & l796;
assign a2706 = a2704 & ~l794;
assign a2708 = a2706 & ~l792;
assign a2710 = ~l796 & l794;
assign a2712 = a2710 & ~l792;
assign a2714 = a2694 & l794;
assign a2716 = a2714 & ~l792;
assign a2718 = l796 & l794;
assign a2720 = a2718 & ~l792;
assign a2722 = a2696 & l792;
assign a2724 = a2706 & l792;
assign a2726 = ~a2724 & a2710;
assign a2728 = ~a2726 & ~a2700;
assign a2730 = ~a2728 & ~a2722;
assign a2732 = ~a2730 & ~a2690;
assign a2734 = ~a2732 & l792;
assign a2736 = ~a2734 & ~a2720;
assign a2738 = ~a2736 & ~a2716;
assign a2740 = ~a2738 & ~a2712;
assign a2742 = ~a2740 & ~a2708;
assign a2744 = ~a2742 & ~a2702;
assign a2746 = ~a2744 & ~a2698;
assign a2748 = ~a2746 & ~a2692;
assign a2750 = ~a2748 & ~l798;
assign a2752 = a2678 & ~l794;
assign a2754 = a2752 & ~l792;
assign a2756 = l798 & ~l794;
assign a2758 = a2756 & ~l792;
assign a2760 = a2678 & l794;
assign a2762 = a2760 & ~l792;
assign a2764 = l798 & l794;
assign a2766 = a2764 & ~l792;
assign a2768 = a2752 & l792;
assign a2770 = ~l794 & l792;
assign a2772 = a2770 & ~a2694;
assign a2774 = a2772 & ~a2768;
assign a2776 = ~a2774 & ~a2766;
assign a2778 = ~l798 & l794;
assign a2780 = a2778 & ~l792;
assign a2782 = ~a2780 & a2776;
assign a2784 = ~a2782 & ~a2716;
assign a2786 = a2784 & ~a2762;
assign a2788 = ~a2786 & ~a2758;
assign a2790 = ~l798 & ~l794;
assign a2792 = a2790 & ~l792;
assign a2794 = ~a2792 & a2788;
assign a2796 = ~a2794 & l796;
assign a2798 = a2796 & ~a2698;
assign a2800 = a2798 & ~a2754;
assign a2802 = a2800 & a2750;
assign a2804 = ~l798 & l796;
assign a2806 = ~a2704 & ~l792;
assign a2808 = a2806 & ~a2804;
assign a2810 = a2694 & ~l792;
assign a2812 = ~a2810 & a2808;
assign a2814 = a2678 & ~l792;
assign a2816 = ~a2814 & a2812;
assign a2818 = ~a2816 & ~l794;
assign a2820 = ~a2818 & a2802;
assign a2822 = ~a2704 & ~l794;
assign a2824 = a2822 & ~a2804;
assign a2826 = a2824 & ~a2696;
assign a2828 = a2826 & ~a2752;
assign a2830 = ~a2828 & ~l792;
assign a2832 = ~a2830 & a2820;
assign a2834 = ~a2832 & l792;
assign a2836 = ~a2834 & a2360;
assign a2838 = ~a2360 & ~l792;
assign a2840 = ~a2838 & ~a2836;
assign a2844 = ~a2832 & l794;
assign a2846 = ~a2844 & a2360;
assign a2848 = ~a2360 & ~l794;
assign a2850 = ~a2848 & ~a2846;
assign a2854 = ~a2832 & l796;
assign a2856 = ~a2854 & a2360;
assign a2858 = ~a2360 & ~l796;
assign a2860 = ~a2858 & ~a2856;
assign a2864 = ~a2832 & ~l798;
assign a2866 = ~a2864 & a2360;
assign a2868 = ~a2360 & ~l798;
assign a2870 = ~a2868 & ~a2866;
assign a2874 = l812 & ~l810;
assign a2876 = l846 & l844;
assign a2878 = a2876 & ~l842;
assign a2880 = a2878 & a2874;
assign a2882 = ~l812 & l810;
assign a2884 = a2882 & a2878;
assign a2886 = l846 & ~l844;
assign a2888 = a2886 & l842;
assign a2890 = a2888 & a2882;
assign a2892 = l802 & ~l800;
assign a2894 = a2876 & l842;
assign a2896 = a2894 & a2882;
assign a2898 = a2896 & a2892;
assign a2900 = ~l802 & ~l800;
assign a2902 = l812 & l810;
assign a2904 = a2886 & ~l842;
assign a2906 = a2904 & a2902;
assign a2908 = a2906 & a2900;
assign a2910 = a2904 & a2874;
assign a2912 = a2910 & a2892;
assign a2914 = a2904 & l848;
assign a2916 = ~a2914 & l804;
assign a2918 = a2916 & ~a2912;
assign a2920 = a2918 & ~a2908;
assign a2922 = ~a2920 & ~a2898;
assign a2924 = ~a2922 & ~a2890;
assign a2926 = ~a2924 & ~a2884;
assign a2928 = ~a2926 & ~a2880;
assign a2932 = ~a2914 & l806;
assign a2934 = a2932 & ~a2912;
assign a2936 = a2934 & ~a2908;
assign a2938 = ~a2936 & ~a2898;
assign a2940 = ~a2938 & ~a2890;
assign a2942 = ~a2940 & ~a2884;
assign a2944 = a2942 & ~a2880;
assign a2948 = ~l802 & l800;
assign a2950 = ~l846 & ~l844;
assign a2952 = a2950 & ~l842;
assign a2954 = a2952 & a2882;
assign a2956 = a2954 & a2948;
assign a2958 = ~l846 & l844;
assign a2960 = a2958 & ~l842;
assign a2962 = a2960 & a2882;
assign a2964 = a2962 & a2900;
assign a2966 = a2948 & a2896;
assign a2968 = ~a2966 & ~l812;
assign a2970 = a2968 & ~a2964;
assign a2972 = a2970 & ~a2956;
assign a2976 = l826 & ~l824;
assign a2978 = a2976 & a2878;
assign a2980 = ~l826 & l824;
assign a2982 = a2980 & a2878;
assign a2984 = a2980 & a2888;
assign a2986 = l816 & ~l814;
assign a2988 = a2980 & a2894;
assign a2990 = a2988 & a2986;
assign a2992 = ~l816 & ~l814;
assign a2994 = l826 & l824;
assign a2996 = a2994 & a2904;
assign a2998 = a2996 & a2992;
assign a3000 = a2976 & a2904;
assign a3002 = a3000 & a2986;
assign a3004 = ~a2914 & l818;
assign a3006 = a3004 & ~a3002;
assign a3008 = a3006 & ~a2998;
assign a3010 = ~a3008 & ~a2990;
assign a3012 = ~a3010 & ~a2984;
assign a3014 = ~a3012 & ~a2982;
assign a3016 = ~a3014 & ~a2978;
assign a3020 = ~a2914 & l820;
assign a3022 = a3020 & ~a3002;
assign a3024 = a3022 & ~a2998;
assign a3026 = ~a3024 & ~a2990;
assign a3028 = ~a3026 & ~a2984;
assign a3030 = ~a3028 & ~a2982;
assign a3032 = a3030 & ~a2978;
assign a3036 = ~l816 & l814;
assign a3038 = a2980 & a2952;
assign a3040 = a3038 & a3036;
assign a3042 = a2980 & a2960;
assign a3044 = a3042 & a2992;
assign a3046 = a3036 & a2988;
assign a3048 = ~a3046 & ~l826;
assign a3050 = a3048 & ~a3044;
assign a3052 = a3050 & ~a3040;
assign a3056 = l840 & ~l838;
assign a3058 = a3056 & a2878;
assign a3060 = ~l840 & l838;
assign a3062 = a3060 & a2878;
assign a3064 = a3060 & a2888;
assign a3066 = l830 & ~l828;
assign a3068 = a3060 & a2894;
assign a3070 = a3068 & a3066;
assign a3072 = ~l830 & ~l828;
assign a3074 = l840 & l838;
assign a3076 = a3074 & a2904;
assign a3078 = a3076 & a3072;
assign a3080 = a3056 & a2904;
assign a3082 = a3080 & a3066;
assign a3084 = ~a2914 & l832;
assign a3086 = a3084 & ~a3082;
assign a3088 = a3086 & ~a3078;
assign a3090 = ~a3088 & ~a3070;
assign a3092 = ~a3090 & ~a3064;
assign a3094 = ~a3092 & ~a3062;
assign a3096 = ~a3094 & ~a3058;
assign a3100 = ~a2914 & l834;
assign a3102 = a3100 & ~a3082;
assign a3104 = a3102 & ~a3078;
assign a3106 = ~a3104 & ~a3070;
assign a3108 = ~a3106 & ~a3064;
assign a3110 = ~a3108 & ~a3062;
assign a3112 = a3110 & ~a3058;
assign a3116 = ~l830 & l828;
assign a3118 = a3060 & a2952;
assign a3120 = a3118 & a3116;
assign a3122 = a3060 & a2960;
assign a3124 = a3122 & a3072;
assign a3126 = a3116 & a3068;
assign a3128 = ~a3126 & ~l840;
assign a3130 = a3128 & ~a3124;
assign a3132 = a3130 & ~a3120;
assign a3136 = ~l860 & l854;
assign a3138 = ~a2980 & ~a2882;
assign a3140 = a2980 & a2882;
assign a3142 = ~a3140 & ~a3060;
assign a3144 = ~a3142 & ~a3138;
assign a3146 = ~a3144 & a2952;
assign a3148 = a3146 & ~a3136;
assign a3150 = ~a2892 & a2874;
assign a3152 = ~a3150 & a2878;
assign a3154 = ~a2986 & a2976;
assign a3156 = ~a3154 & a3152;
assign a3158 = ~a3066 & a3056;
assign a3160 = ~a3158 & a3156;
assign a3162 = ~a2900 & a2882;
assign a3164 = ~a3162 & a2960;
assign a3166 = ~a2992 & a2980;
assign a3168 = ~a3166 & a3164;
assign a3170 = ~a3072 & a3060;
assign a3172 = ~a3170 & a3168;
assign a3174 = ~a3116 & a3060;
assign a3176 = ~a3036 & a2980;
assign a3178 = ~a2948 & a2882;
assign a3180 = ~a3178 & a2960;
assign a3182 = a3180 & ~a3176;
assign a3184 = a3182 & ~a3174;
assign a3186 = ~a3066 & a3060;
assign a3188 = ~a2892 & a2882;
assign a3190 = ~a2986 & a2980;
assign a3192 = ~a3190 & ~a3188;
assign a3194 = a3192 & ~a3186;
assign a3196 = ~a3178 & ~a3176;
assign a3198 = a3196 & ~a3174;
assign a3200 = ~a3198 & ~a3194;
assign a3202 = ~a3200 & ~a2886;
assign a3204 = a3202 & a2894;
assign a3206 = a3204 & ~a2950;
assign a3208 = ~a3206 & l842;
assign a3210 = ~a3208 & ~a3184;
assign a3212 = ~a3210 & ~a3172;
assign a3214 = a3212 & ~a3160;
assign a3216 = a3214 & ~a3148;
assign a3220 = a2888 & ~l856;
assign a3222 = a2950 & l842;
assign a3224 = l846 & l842;
assign a3226 = a3224 & l856;
assign a3228 = ~a3226 & a3222;
assign a3230 = ~a3228 & ~l844;
assign a3232 = a3230 & ~a3220;
assign a3234 = ~a3232 & ~a3184;
assign a3236 = a3234 & ~a3172;
assign a3238 = ~a3236 & ~a3160;
assign a3240 = a3238 & ~a3148;
assign a3244 = a2888 & l856;
assign a3246 = ~a3190 & ~a3186;
assign a3248 = a3246 & ~a3188;
assign a3250 = a3248 & a2894;
assign a3252 = ~a3250 & l846;
assign a3254 = ~a3252 & ~a3222;
assign a3256 = ~a3254 & ~a3244;
assign a3258 = ~a3256 & ~a3220;
assign a3260 = a3258 & ~a3184;
assign a3262 = a3260 & ~a3172;
assign a3264 = ~a3262 & ~a3160;
assign a3266 = ~a3264 & ~a3148;
assign a3270 = ~l866 & ~l864;
assign a3272 = ~a3270 & l862;
assign a3274 = a3272 & l860;
assign a3276 = a3274 & a2952;
assign a3278 = ~a3276 & ~l858;
assign a3282 = ~l864 & ~l862;
assign a3284 = a3282 & ~l860;
assign a3286 = l866 & ~l864;
assign a3288 = a3286 & ~l862;
assign a3290 = a3288 & ~l860;
assign a3292 = l864 & ~l862;
assign a3294 = a3292 & ~l860;
assign a3296 = l866 & l864;
assign a3298 = a3296 & ~l862;
assign a3300 = a3298 & ~l860;
assign a3302 = ~l864 & l862;
assign a3304 = a3302 & ~l860;
assign a3306 = a3286 & l862;
assign a3308 = a3306 & ~l860;
assign a3310 = l864 & l862;
assign a3312 = a3310 & ~l860;
assign a3314 = a3288 & l860;
assign a3316 = a3298 & l860;
assign a3318 = ~a3316 & a3302;
assign a3320 = ~a3318 & ~a3292;
assign a3322 = ~a3320 & ~a3314;
assign a3324 = ~a3322 & ~a3282;
assign a3326 = ~a3324 & l860;
assign a3328 = ~a3326 & ~a3312;
assign a3330 = ~a3328 & ~a3308;
assign a3332 = ~a3330 & ~a3304;
assign a3334 = ~a3332 & ~a3300;
assign a3336 = ~a3334 & ~a3294;
assign a3338 = ~a3336 & ~a3290;
assign a3340 = ~a3338 & ~a3284;
assign a3342 = ~a3340 & ~l866;
assign a3344 = a3270 & ~l862;
assign a3346 = a3344 & ~l860;
assign a3348 = l866 & ~l862;
assign a3350 = a3348 & ~l860;
assign a3352 = a3270 & l862;
assign a3354 = a3352 & ~l860;
assign a3356 = l866 & l862;
assign a3358 = a3356 & ~l860;
assign a3360 = a3344 & l860;
assign a3362 = ~l862 & l860;
assign a3364 = a3362 & ~a3286;
assign a3366 = a3364 & ~a3360;
assign a3368 = ~a3366 & ~a3358;
assign a3370 = ~l866 & l862;
assign a3372 = a3370 & ~l860;
assign a3374 = ~a3372 & a3368;
assign a3376 = ~a3374 & ~a3308;
assign a3378 = a3376 & ~a3354;
assign a3380 = ~a3378 & ~a3350;
assign a3382 = ~l866 & ~l862;
assign a3384 = a3382 & ~l860;
assign a3386 = ~a3384 & a3380;
assign a3388 = ~a3386 & l864;
assign a3390 = a3388 & ~a3290;
assign a3392 = a3390 & ~a3346;
assign a3394 = a3392 & a3342;
assign a3396 = ~l866 & l864;
assign a3398 = ~a3296 & ~l860;
assign a3400 = a3398 & ~a3396;
assign a3402 = a3286 & ~l860;
assign a3404 = ~a3402 & a3400;
assign a3406 = a3270 & ~l860;
assign a3408 = ~a3406 & a3404;
assign a3410 = ~a3408 & ~l862;
assign a3412 = ~a3410 & a3394;
assign a3414 = ~a3296 & ~l862;
assign a3416 = a3414 & ~a3396;
assign a3418 = a3416 & ~a3288;
assign a3420 = a3418 & ~a3344;
assign a3422 = ~a3420 & ~l860;
assign a3424 = ~a3422 & a3412;
assign a3426 = ~a3424 & l860;
assign a3428 = ~a3426 & a2952;
assign a3430 = ~a2952 & ~l860;
assign a3432 = ~a3430 & ~a3428;
assign a3436 = ~a3424 & l862;
assign a3438 = ~a3436 & a2952;
assign a3440 = ~a2952 & ~l862;
assign a3442 = ~a3440 & ~a3438;
assign a3446 = ~a3424 & l864;
assign a3448 = ~a3446 & a2952;
assign a3450 = ~a2952 & ~l864;
assign a3452 = ~a3450 & ~a3448;
assign a3456 = ~a3424 & ~l866;
assign a3458 = ~a3456 & a2952;
assign a3460 = ~a2952 & ~l866;
assign a3462 = ~a3460 & ~a3458;
assign a3466 = ~a2038 & l870;
assign a3468 = ~a3466 & ~a1446;
assign a3472 = ~l1084 & ~l1082;
assign a3474 = ~a3472 & l868;
assign a3476 = ~a3474 & ~l1076;
assign a3480 = ~l872 & l712;
assign a3482 = ~a3480 & l874;
assign a3484 = ~a3482 & ~a3472;
assign a3486 = ~a3484 & ~l1078;
assign a3490 = l872 & l712;
assign a3492 = ~a3490 & ~a3472;
assign a3494 = ~a3492 & ~l1080;
assign a3500 = ~l872 & ~l712;
assign a3502 = l868 & ~i258;
assign a3504 = a3480 & ~l874;
assign a3506 = ~a3504 & ~a3502;
assign a3508 = a3506 & ~a3500;
assign a3510 = l476 & ~i2;
assign a3512 = ~l476 & i2;
assign a3514 = ~a3512 & ~a3510;
assign a3516 = a3514 & a3508;
assign a3518 = l478 & ~i4;
assign a3520 = ~l478 & i4;
assign a3522 = ~a3520 & ~a3518;
assign a3524 = a3522 & a3516;
assign a3526 = l480 & ~i6;
assign a3528 = ~l480 & i6;
assign a3530 = ~a3528 & ~a3526;
assign a3532 = a3530 & a3524;
assign a3534 = l482 & ~i8;
assign a3536 = ~l482 & i8;
assign a3538 = ~a3536 & ~a3534;
assign a3540 = a3538 & a3532;
assign a3542 = l484 & ~i10;
assign a3544 = ~l484 & i10;
assign a3546 = ~a3544 & ~a3542;
assign a3548 = a3546 & a3540;
assign a3550 = l486 & ~i12;
assign a3552 = ~l486 & i12;
assign a3554 = ~a3552 & ~a3550;
assign a3556 = a3554 & a3548;
assign a3558 = l488 & ~i14;
assign a3560 = ~l488 & i14;
assign a3562 = ~a3560 & ~a3558;
assign a3564 = a3562 & a3556;
assign a3566 = l490 & ~i16;
assign a3568 = ~l490 & i16;
assign a3570 = ~a3568 & ~a3566;
assign a3572 = a3570 & a3564;
assign a3574 = l492 & ~i18;
assign a3576 = ~l492 & i18;
assign a3578 = ~a3576 & ~a3574;
assign a3580 = a3578 & a3572;
assign a3582 = l494 & ~i20;
assign a3584 = ~l494 & i20;
assign a3586 = ~a3584 & ~a3582;
assign a3588 = a3586 & a3580;
assign a3590 = l496 & ~i22;
assign a3592 = ~l496 & i22;
assign a3594 = ~a3592 & ~a3590;
assign a3596 = a3594 & a3588;
assign a3598 = l498 & ~i24;
assign a3600 = ~l498 & i24;
assign a3602 = ~a3600 & ~a3598;
assign a3604 = a3602 & a3596;
assign a3606 = l500 & ~i26;
assign a3608 = ~l500 & i26;
assign a3610 = ~a3608 & ~a3606;
assign a3612 = a3610 & a3604;
assign a3614 = l502 & ~i28;
assign a3616 = ~l502 & i28;
assign a3618 = ~a3616 & ~a3614;
assign a3620 = a3618 & a3612;
assign a3622 = l504 & ~i30;
assign a3624 = ~l504 & i30;
assign a3626 = ~a3624 & ~a3622;
assign a3628 = a3626 & a3620;
assign a3630 = l506 & ~i32;
assign a3632 = ~l506 & i32;
assign a3634 = ~a3632 & ~a3630;
assign a3636 = a3634 & a3628;
assign a3638 = l508 & ~i34;
assign a3640 = ~l508 & i34;
assign a3642 = ~a3640 & ~a3638;
assign a3644 = a3642 & a3636;
assign a3646 = l510 & ~i36;
assign a3648 = ~l510 & i36;
assign a3650 = ~a3648 & ~a3646;
assign a3652 = a3650 & a3644;
assign a3654 = l512 & ~i38;
assign a3656 = ~l512 & i38;
assign a3658 = ~a3656 & ~a3654;
assign a3660 = a3658 & a3652;
assign a3662 = l514 & ~i40;
assign a3664 = ~l514 & i40;
assign a3666 = ~a3664 & ~a3662;
assign a3668 = a3666 & a3660;
assign a3670 = l516 & ~i42;
assign a3672 = ~l516 & i42;
assign a3674 = ~a3672 & ~a3670;
assign a3676 = a3674 & a3668;
assign a3678 = l518 & ~i44;
assign a3680 = ~l518 & i44;
assign a3682 = ~a3680 & ~a3678;
assign a3684 = a3682 & a3676;
assign a3686 = l520 & ~i46;
assign a3688 = ~l520 & i46;
assign a3690 = ~a3688 & ~a3686;
assign a3692 = a3690 & a3684;
assign a3694 = l522 & ~i48;
assign a3696 = ~l522 & i48;
assign a3698 = ~a3696 & ~a3694;
assign a3700 = a3698 & a3692;
assign a3702 = l524 & ~i50;
assign a3704 = ~l524 & i50;
assign a3706 = ~a3704 & ~a3702;
assign a3708 = a3706 & a3700;
assign a3710 = l526 & ~i52;
assign a3712 = ~l526 & i52;
assign a3714 = ~a3712 & ~a3710;
assign a3716 = a3714 & a3708;
assign a3718 = l528 & ~i54;
assign a3720 = ~l528 & i54;
assign a3722 = ~a3720 & ~a3718;
assign a3724 = a3722 & a3716;
assign a3726 = l530 & ~i56;
assign a3728 = ~l530 & i56;
assign a3730 = ~a3728 & ~a3726;
assign a3732 = a3730 & a3724;
assign a3734 = l532 & ~i58;
assign a3736 = ~l532 & i58;
assign a3738 = ~a3736 & ~a3734;
assign a3740 = a3738 & a3732;
assign a3742 = l534 & ~i60;
assign a3744 = ~l534 & i60;
assign a3746 = ~a3744 & ~a3742;
assign a3748 = a3746 & a3740;
assign a3750 = l536 & ~i62;
assign a3752 = ~l536 & i62;
assign a3754 = ~a3752 & ~a3750;
assign a3756 = a3754 & a3748;
assign a3758 = l538 & ~i64;
assign a3760 = ~l538 & i64;
assign a3762 = ~a3760 & ~a3758;
assign a3764 = a3762 & a3756;
assign a3766 = l540 & ~i66;
assign a3768 = ~l540 & i66;
assign a3770 = ~a3768 & ~a3766;
assign a3772 = a3770 & a3764;
assign a3774 = l542 & ~i68;
assign a3776 = ~l542 & i68;
assign a3778 = ~a3776 & ~a3774;
assign a3780 = a3778 & a3772;
assign a3782 = l544 & ~i70;
assign a3784 = ~l544 & i70;
assign a3786 = ~a3784 & ~a3782;
assign a3788 = a3786 & a3780;
assign a3790 = l546 & ~i72;
assign a3792 = ~l546 & i72;
assign a3794 = ~a3792 & ~a3790;
assign a3796 = a3794 & a3788;
assign a3798 = l548 & ~i74;
assign a3800 = ~l548 & i74;
assign a3802 = ~a3800 & ~a3798;
assign a3804 = a3802 & a3796;
assign a3806 = l550 & ~i76;
assign a3808 = ~l550 & i76;
assign a3810 = ~a3808 & ~a3806;
assign a3812 = a3810 & a3804;
assign a3814 = l552 & ~i78;
assign a3816 = ~l552 & i78;
assign a3818 = ~a3816 & ~a3814;
assign a3820 = a3818 & a3812;
assign a3822 = l554 & ~i80;
assign a3824 = ~l554 & i80;
assign a3826 = ~a3824 & ~a3822;
assign a3828 = a3826 & a3820;
assign a3830 = l556 & ~i82;
assign a3832 = ~l556 & i82;
assign a3834 = ~a3832 & ~a3830;
assign a3836 = a3834 & a3828;
assign a3838 = l558 & ~i84;
assign a3840 = ~l558 & i84;
assign a3842 = ~a3840 & ~a3838;
assign a3844 = a3842 & a3836;
assign a3846 = l560 & ~i86;
assign a3848 = ~l560 & i86;
assign a3850 = ~a3848 & ~a3846;
assign a3852 = a3850 & a3844;
assign a3854 = l562 & ~i88;
assign a3856 = ~l562 & i88;
assign a3858 = ~a3856 & ~a3854;
assign a3860 = a3858 & a3852;
assign a3862 = l564 & ~i90;
assign a3864 = ~l564 & i90;
assign a3866 = ~a3864 & ~a3862;
assign a3868 = a3866 & a3860;
assign a3870 = l566 & ~i92;
assign a3872 = ~l566 & i92;
assign a3874 = ~a3872 & ~a3870;
assign a3876 = a3874 & a3868;
assign a3878 = l568 & ~i94;
assign a3880 = ~l568 & i94;
assign a3882 = ~a3880 & ~a3878;
assign a3884 = a3882 & a3876;
assign a3886 = l570 & ~i96;
assign a3888 = ~l570 & i96;
assign a3890 = ~a3888 & ~a3886;
assign a3892 = a3890 & a3884;
assign a3894 = l572 & ~i98;
assign a3896 = ~l572 & i98;
assign a3898 = ~a3896 & ~a3894;
assign a3900 = a3898 & a3892;
assign a3902 = l574 & ~i100;
assign a3904 = ~l574 & i100;
assign a3906 = ~a3904 & ~a3902;
assign a3908 = a3906 & a3900;
assign a3910 = l576 & ~i102;
assign a3912 = ~l576 & i102;
assign a3914 = ~a3912 & ~a3910;
assign a3916 = a3914 & a3908;
assign a3918 = l578 & ~i104;
assign a3920 = ~l578 & i104;
assign a3922 = ~a3920 & ~a3918;
assign a3924 = a3922 & a3916;
assign a3926 = l580 & ~i106;
assign a3928 = ~l580 & i106;
assign a3930 = ~a3928 & ~a3926;
assign a3932 = a3930 & a3924;
assign a3934 = l582 & ~i108;
assign a3936 = ~l582 & i108;
assign a3938 = ~a3936 & ~a3934;
assign a3940 = a3938 & a3932;
assign a3942 = l584 & ~i110;
assign a3944 = ~l584 & i110;
assign a3946 = ~a3944 & ~a3942;
assign a3948 = a3946 & a3940;
assign a3950 = l586 & ~i112;
assign a3952 = ~l586 & i112;
assign a3954 = ~a3952 & ~a3950;
assign a3956 = a3954 & a3948;
assign a3958 = l588 & ~i114;
assign a3960 = ~l588 & i114;
assign a3962 = ~a3960 & ~a3958;
assign a3964 = a3962 & a3956;
assign a3966 = l590 & ~i116;
assign a3968 = ~l590 & i116;
assign a3970 = ~a3968 & ~a3966;
assign a3972 = a3970 & a3964;
assign a3974 = l592 & ~i118;
assign a3976 = ~l592 & i118;
assign a3978 = ~a3976 & ~a3974;
assign a3980 = a3978 & a3972;
assign a3982 = l594 & ~i120;
assign a3984 = ~l594 & i120;
assign a3986 = ~a3984 & ~a3982;
assign a3988 = a3986 & a3980;
assign a3990 = l604 & ~i126;
assign a3992 = ~l604 & i126;
assign a3994 = ~a3992 & ~a3990;
assign a3996 = a3994 & a3988;
assign a3998 = a1184 & ~l608;
assign a4000 = a3998 & a1124;
assign a4002 = ~a4000 & a1190;
assign a4004 = ~a4002 & l606;
assign a4006 = a4004 & ~a1180;
assign a4008 = a4006 & ~i128;
assign a4010 = ~a4006 & i128;
assign a4012 = ~a4010 & ~a4008;
assign a4014 = a4012 & a3996;
assign a4016 = l618 & ~i134;
assign a4018 = ~l618 & i134;
assign a4020 = ~a4018 & ~a4016;
assign a4022 = a4020 & a4014;
assign a4024 = a1184 & ~l622;
assign a4026 = a4024 & a1216;
assign a4028 = ~a4026 & a1270;
assign a4030 = ~a4028 & l620;
assign a4032 = a4030 & ~a1264;
assign a4034 = a4032 & ~i136;
assign a4036 = ~a4032 & i136;
assign a4038 = ~a4036 & ~a4034;
assign a4040 = a4038 & a4022;
assign a4042 = l632 & ~i142;
assign a4044 = ~l632 & i142;
assign a4046 = ~a4044 & ~a4042;
assign a4048 = a4046 & a4040;
assign a4050 = a1184 & ~l636;
assign a4052 = a4050 & a1296;
assign a4054 = ~a4052 & a1350;
assign a4056 = ~a4054 & l634;
assign a4058 = a4056 & ~a1344;
assign a4060 = a4058 & ~i144;
assign a4062 = ~a4058 & i144;
assign a4064 = ~a4062 & ~a4060;
assign a4066 = a4064 & a4048;
assign a4068 = a1362 & ~a1284;
assign a4070 = ~a4068 & a1102;
assign a4072 = ~a1102 & ~l644;
assign a4074 = ~a4072 & ~a4070;
assign a4076 = a4074 & ~i146;
assign a4078 = ~a4074 & i146;
assign a4080 = ~a4078 & ~a4076;
assign a4082 = a4080 & a4066;
assign a4084 = ~a1286 & ~l646;
assign a4086 = ~a4084 & ~a1206;
assign a4088 = a4086 & ~a1108;
assign a4090 = a4088 & ~i148;
assign a4092 = ~a4088 & i148;
assign a4094 = ~a4092 & ~a4090;
assign a4096 = a4094 & a4082;
assign a4098 = ~a1286 & l648;
assign a4100 = ~a4098 & ~a1206;
assign a4102 = ~a4100 & ~a1108;
assign a4104 = a4102 & ~i150;
assign a4106 = ~a4102 & i150;
assign a4108 = ~a4106 & ~a4104;
assign a4110 = a4108 & a4096;
assign a4112 = l650 & ~i152;
assign a4114 = ~l650 & i152;
assign a4116 = ~a4114 & ~a4112;
assign a4118 = a4116 & a4110;
assign a4120 = a1184 & l1086;
assign a4122 = ~a1184 & ~l652;
assign a4124 = ~a4122 & ~a4120;
assign a4126 = a4124 & ~i154;
assign a4128 = ~a4124 & i154;
assign a4130 = ~a4128 & ~a4126;
assign a4132 = a4130 & a4118;
assign a4134 = l672 & ~i160;
assign a4136 = ~l672 & i160;
assign a4138 = ~a4136 & ~a4134;
assign a4140 = a4138 & a4132;
assign a4142 = a1776 & ~l676;
assign a4144 = a4142 & a1716;
assign a4146 = ~a4144 & a1782;
assign a4148 = ~a4146 & l674;
assign a4150 = a4148 & ~a1772;
assign a4152 = a4150 & ~i162;
assign a4154 = ~a4150 & i162;
assign a4156 = ~a4154 & ~a4152;
assign a4158 = a4156 & a4140;
assign a4160 = l686 & ~i168;
assign a4162 = ~l686 & i168;
assign a4164 = ~a4162 & ~a4160;
assign a4166 = a4164 & a4158;
assign a4168 = a1776 & ~l690;
assign a4170 = a4168 & a1808;
assign a4172 = ~a4170 & a1862;
assign a4174 = ~a4172 & l688;
assign a4176 = a4174 & ~a1856;
assign a4178 = a4176 & ~i170;
assign a4180 = ~a4176 & i170;
assign a4182 = ~a4180 & ~a4178;
assign a4184 = a4182 & a4166;
assign a4186 = l700 & ~i176;
assign a4188 = ~l700 & i176;
assign a4190 = ~a4188 & ~a4186;
assign a4192 = a4190 & a4184;
assign a4194 = a1776 & ~l704;
assign a4196 = a4194 & a1888;
assign a4198 = ~a4196 & a1942;
assign a4200 = ~a4198 & l702;
assign a4202 = a4200 & ~a1936;
assign a4204 = a4202 & ~i178;
assign a4206 = ~a4202 & i178;
assign a4208 = ~a4206 & ~a4204;
assign a4210 = a4208 & a4192;
assign a4212 = a1954 & ~a1876;
assign a4214 = ~a4212 & a1694;
assign a4216 = ~a1694 & ~l712;
assign a4218 = ~a4216 & ~a4214;
assign a4220 = a4218 & ~i180;
assign a4222 = ~a4218 & i180;
assign a4224 = ~a4222 & ~a4220;
assign a4226 = a4224 & a4210;
assign a4228 = ~a1878 & ~l714;
assign a4230 = ~a4228 & ~a1798;
assign a4232 = a4230 & ~a1700;
assign a4234 = a4232 & ~i182;
assign a4236 = ~a4232 & i182;
assign a4238 = ~a4236 & ~a4234;
assign a4240 = a4238 & a4226;
assign a4242 = ~a1878 & l716;
assign a4244 = ~a4242 & ~a1798;
assign a4246 = ~a4244 & ~a1700;
assign a4248 = a4246 & ~i184;
assign a4250 = ~a4246 & i184;
assign a4252 = ~a4250 & ~a4248;
assign a4254 = a4252 & a4240;
assign a4256 = l718 & ~i186;
assign a4258 = ~l718 & i186;
assign a4260 = ~a4258 & ~a4256;
assign a4262 = a4260 & a4254;
assign a4264 = a1776 & l1088;
assign a4266 = ~a1776 & ~l720;
assign a4268 = ~a4266 & ~a4264;
assign a4270 = a4268 & ~i188;
assign a4272 = ~a4268 & i188;
assign a4274 = ~a4272 & ~a4270;
assign a4276 = a4274 & a4262;
assign a4278 = l740 & ~i194;
assign a4280 = ~l740 & i194;
assign a4282 = ~a4280 & ~a4278;
assign a4284 = a4282 & a4276;
assign a4286 = a2368 & ~l744;
assign a4288 = a4286 & a2308;
assign a4290 = ~a4288 & a2374;
assign a4292 = ~a4290 & l742;
assign a4294 = a4292 & ~a2364;
assign a4296 = a4294 & ~i196;
assign a4298 = ~a4294 & i196;
assign a4300 = ~a4298 & ~a4296;
assign a4302 = a4300 & a4284;
assign a4304 = l754 & ~i202;
assign a4306 = ~l754 & i202;
assign a4308 = ~a4306 & ~a4304;
assign a4310 = a4308 & a4302;
assign a4312 = a2368 & ~l758;
assign a4314 = a4312 & a2400;
assign a4316 = ~a4314 & a2454;
assign a4318 = ~a4316 & l756;
assign a4320 = a4318 & ~a2448;
assign a4322 = a4320 & ~i204;
assign a4324 = ~a4320 & i204;
assign a4326 = ~a4324 & ~a4322;
assign a4328 = a4326 & a4310;
assign a4330 = l768 & ~i210;
assign a4332 = ~l768 & i210;
assign a4334 = ~a4332 & ~a4330;
assign a4336 = a4334 & a4328;
assign a4338 = a2368 & ~l772;
assign a4340 = a4338 & a2480;
assign a4342 = ~a4340 & a2534;
assign a4344 = ~a4342 & l770;
assign a4346 = a4344 & ~a2528;
assign a4348 = a4346 & ~i212;
assign a4350 = ~a4346 & i212;
assign a4352 = ~a4350 & ~a4348;
assign a4354 = a4352 & a4336;
assign a4356 = a2546 & ~a2468;
assign a4358 = ~a4356 & a2286;
assign a4360 = ~a2286 & ~l780;
assign a4362 = ~a4360 & ~a4358;
assign a4364 = a4362 & ~i214;
assign a4366 = ~a4362 & i214;
assign a4368 = ~a4366 & ~a4364;
assign a4370 = a4368 & a4354;
assign a4372 = ~a2470 & ~l782;
assign a4374 = ~a4372 & ~a2390;
assign a4376 = a4374 & ~a2292;
assign a4378 = a4376 & ~i216;
assign a4380 = ~a4376 & i216;
assign a4382 = ~a4380 & ~a4378;
assign a4384 = a4382 & a4370;
assign a4386 = ~a2470 & l784;
assign a4388 = ~a4386 & ~a2390;
assign a4390 = ~a4388 & ~a2292;
assign a4392 = a4390 & ~i218;
assign a4394 = ~a4390 & i218;
assign a4396 = ~a4394 & ~a4392;
assign a4398 = a4396 & a4384;
assign a4400 = l786 & ~i220;
assign a4402 = ~l786 & i220;
assign a4404 = ~a4402 & ~a4400;
assign a4406 = a4404 & a4398;
assign a4408 = a2368 & l1090;
assign a4410 = ~a2368 & ~l788;
assign a4412 = ~a4410 & ~a4408;
assign a4414 = a4412 & ~i222;
assign a4416 = ~a4412 & i222;
assign a4418 = ~a4416 & ~a4414;
assign a4420 = a4418 & a4406;
assign a4422 = l808 & ~i228;
assign a4424 = ~l808 & i228;
assign a4426 = ~a4424 & ~a4422;
assign a4428 = a4426 & a4420;
assign a4430 = a2960 & ~l812;
assign a4432 = a4430 & a2900;
assign a4434 = ~a4432 & a2966;
assign a4436 = ~a4434 & l810;
assign a4438 = a4436 & ~a2956;
assign a4440 = a4438 & ~i230;
assign a4442 = ~a4438 & i230;
assign a4444 = ~a4442 & ~a4440;
assign a4446 = a4444 & a4428;
assign a4448 = l822 & ~i236;
assign a4450 = ~l822 & i236;
assign a4452 = ~a4450 & ~a4448;
assign a4454 = a4452 & a4446;
assign a4456 = a2960 & ~l826;
assign a4458 = a4456 & a2992;
assign a4460 = ~a4458 & a3046;
assign a4462 = ~a4460 & l824;
assign a4464 = a4462 & ~a3040;
assign a4466 = a4464 & ~i238;
assign a4468 = ~a4464 & i238;
assign a4470 = ~a4468 & ~a4466;
assign a4472 = a4470 & a4454;
assign a4474 = l836 & ~i244;
assign a4476 = ~l836 & i244;
assign a4478 = ~a4476 & ~a4474;
assign a4480 = a4478 & a4472;
assign a4482 = a2960 & ~l840;
assign a4484 = a4482 & a3072;
assign a4486 = ~a4484 & a3126;
assign a4488 = ~a4486 & l838;
assign a4490 = a4488 & ~a3120;
assign a4492 = a4490 & ~i246;
assign a4494 = ~a4490 & i246;
assign a4496 = ~a4494 & ~a4492;
assign a4498 = a4496 & a4480;
assign a4500 = a3138 & ~a3060;
assign a4502 = ~a4500 & a2878;
assign a4504 = ~a2878 & ~l848;
assign a4506 = ~a4504 & ~a4502;
assign a4508 = a4506 & ~i248;
assign a4510 = ~a4506 & i248;
assign a4512 = ~a4510 & ~a4508;
assign a4514 = a4512 & a4498;
assign a4516 = ~a3062 & ~l850;
assign a4518 = ~a4516 & ~a2982;
assign a4520 = a4518 & ~a2884;
assign a4522 = a4520 & ~i250;
assign a4524 = ~a4520 & i250;
assign a4526 = ~a4524 & ~a4522;
assign a4528 = a4526 & a4514;
assign a4530 = ~a3062 & l852;
assign a4532 = ~a4530 & ~a2982;
assign a4534 = ~a4532 & ~a2884;
assign a4536 = a4534 & ~i252;
assign a4538 = ~a4534 & i252;
assign a4540 = ~a4538 & ~a4536;
assign a4542 = a4540 & a4528;
assign a4544 = l854 & ~i254;
assign a4546 = ~l854 & i254;
assign a4548 = ~a4546 & ~a4544;
assign a4550 = a4548 & a4542;
assign a4552 = a2960 & l1092;
assign a4554 = ~a2960 & ~l856;
assign a4556 = ~a4554 & ~a4552;
assign a4558 = a4556 & ~i256;
assign a4560 = ~a4556 & i256;
assign a4562 = ~a4560 & ~a4558;
assign a4564 = a4562 & a4550;
assign a4566 = ~l1084 & l1082;
assign a4568 = a4566 & ~l600;
assign a4570 = ~a4566 & ~l876;
assign a4572 = ~a4570 & ~a4568;
assign a4574 = a4572 & ~i264;
assign a4576 = ~a4572 & i264;
assign a4578 = ~a4576 & ~a4574;
assign a4580 = a4578 & a4564;
assign a4582 = ~a4566 & ~l878;
assign a4584 = a4566 & l602;
assign a4586 = ~a4584 & ~a4582;
assign a4588 = a4586 & ~i266;
assign a4590 = ~a4586 & i266;
assign a4592 = ~a4590 & ~a4588;
assign a4594 = a4592 & a4580;
assign a4596 = a4566 & ~l606;
assign a4598 = ~a4566 & ~l880;
assign a4600 = ~a4598 & ~a4596;
assign a4602 = a4600 & ~i268;
assign a4604 = ~a4600 & i268;
assign a4606 = ~a4604 & ~a4602;
assign a4608 = a4606 & a4594;
assign a4610 = ~a4566 & ~l882;
assign a4612 = a4566 & l608;
assign a4614 = ~a4612 & ~a4610;
assign a4616 = a4614 & ~i270;
assign a4618 = ~a4614 & i270;
assign a4620 = ~a4618 & ~a4616;
assign a4622 = a4620 & a4608;
assign a4624 = a4566 & ~l614;
assign a4626 = ~a4566 & ~l884;
assign a4628 = ~a4626 & ~a4624;
assign a4630 = a4628 & ~i272;
assign a4632 = ~a4628 & i272;
assign a4634 = ~a4632 & ~a4630;
assign a4636 = a4634 & a4622;
assign a4638 = ~a4566 & ~l886;
assign a4640 = a4566 & l616;
assign a4642 = ~a4640 & ~a4638;
assign a4644 = a4642 & ~i274;
assign a4646 = ~a4642 & i274;
assign a4648 = ~a4646 & ~a4644;
assign a4650 = a4648 & a4636;
assign a4652 = a4566 & ~l620;
assign a4654 = ~a4566 & ~l888;
assign a4656 = ~a4654 & ~a4652;
assign a4658 = a4656 & ~i276;
assign a4660 = ~a4656 & i276;
assign a4662 = ~a4660 & ~a4658;
assign a4664 = a4662 & a4650;
assign a4666 = ~a4566 & ~l890;
assign a4668 = a4566 & l622;
assign a4670 = ~a4668 & ~a4666;
assign a4672 = a4670 & ~i278;
assign a4674 = ~a4670 & i278;
assign a4676 = ~a4674 & ~a4672;
assign a4678 = a4676 & a4664;
assign a4680 = a4566 & ~l628;
assign a4682 = ~a4566 & ~l892;
assign a4684 = ~a4682 & ~a4680;
assign a4686 = a4684 & ~i280;
assign a4688 = ~a4684 & i280;
assign a4690 = ~a4688 & ~a4686;
assign a4692 = a4690 & a4678;
assign a4694 = ~a4566 & ~l894;
assign a4696 = a4566 & l630;
assign a4698 = ~a4696 & ~a4694;
assign a4700 = a4698 & ~i282;
assign a4702 = ~a4698 & i282;
assign a4704 = ~a4702 & ~a4700;
assign a4706 = a4704 & a4692;
assign a4708 = a4566 & ~l634;
assign a4710 = ~a4566 & ~l896;
assign a4712 = ~a4710 & ~a4708;
assign a4714 = a4712 & ~i284;
assign a4716 = ~a4712 & i284;
assign a4718 = ~a4716 & ~a4714;
assign a4720 = a4718 & a4706;
assign a4722 = ~a4566 & ~l898;
assign a4724 = a4566 & l636;
assign a4726 = ~a4724 & ~a4722;
assign a4728 = a4726 & ~i286;
assign a4730 = ~a4726 & i286;
assign a4732 = ~a4730 & ~a4728;
assign a4734 = a4732 & a4720;
assign a4736 = a4566 & ~l638;
assign a4738 = ~a4566 & ~l900;
assign a4740 = ~a4738 & ~a4736;
assign a4742 = a4740 & ~i288;
assign a4744 = ~a4740 & i288;
assign a4746 = ~a4744 & ~a4742;
assign a4748 = a4746 & a4734;
assign a4750 = a4566 & ~l640;
assign a4752 = ~a4566 & ~l902;
assign a4754 = ~a4752 & ~a4750;
assign a4756 = a4754 & ~i290;
assign a4758 = ~a4754 & i290;
assign a4760 = ~a4758 & ~a4756;
assign a4762 = a4760 & a4748;
assign a4764 = ~a4566 & ~l904;
assign a4766 = a4566 & l642;
assign a4768 = ~a4766 & ~a4764;
assign a4770 = a4768 & ~i292;
assign a4772 = ~a4768 & i292;
assign a4774 = ~a4772 & ~a4770;
assign a4776 = a4774 & a4762;
assign a4778 = a4566 & ~l644;
assign a4780 = ~a4566 & ~l906;
assign a4782 = ~a4780 & ~a4778;
assign a4784 = a4782 & ~i294;
assign a4786 = ~a4782 & i294;
assign a4788 = ~a4786 & ~a4784;
assign a4790 = a4788 & a4776;
assign a4792 = a4566 & ~l646;
assign a4794 = ~a4566 & ~l908;
assign a4796 = ~a4794 & ~a4792;
assign a4798 = a4796 & ~i296;
assign a4800 = ~a4796 & i296;
assign a4802 = ~a4800 & ~a4798;
assign a4804 = a4802 & a4790;
assign a4806 = a4566 & ~l648;
assign a4808 = ~a4566 & ~l910;
assign a4810 = ~a4808 & ~a4806;
assign a4812 = a4810 & ~i298;
assign a4814 = ~a4810 & i298;
assign a4816 = ~a4814 & ~a4812;
assign a4818 = a4816 & a4804;
assign a4820 = a4566 & ~l652;
assign a4822 = ~a4566 & ~l912;
assign a4824 = ~a4822 & ~a4820;
assign a4826 = a4824 & ~i300;
assign a4828 = ~a4824 & i300;
assign a4830 = ~a4828 & ~a4826;
assign a4832 = a4830 & a4818;
assign a4834 = a4566 & ~l654;
assign a4836 = ~a4566 & ~l914;
assign a4838 = ~a4836 & ~a4834;
assign a4840 = a4838 & ~i302;
assign a4842 = ~a4838 & i302;
assign a4844 = ~a4842 & ~a4840;
assign a4846 = a4844 & a4832;
assign a4848 = a4566 & ~l656;
assign a4850 = ~a4566 & ~l916;
assign a4852 = ~a4850 & ~a4848;
assign a4854 = a4852 & ~i304;
assign a4856 = ~a4852 & i304;
assign a4858 = ~a4856 & ~a4854;
assign a4860 = a4858 & a4846;
assign a4862 = a4566 & ~l658;
assign a4864 = ~a4566 & ~l918;
assign a4866 = ~a4864 & ~a4862;
assign a4868 = a4866 & ~i306;
assign a4870 = ~a4866 & i306;
assign a4872 = ~a4870 & ~a4868;
assign a4874 = a4872 & a4860;
assign a4876 = a4566 & ~l660;
assign a4878 = ~a4566 & ~l920;
assign a4880 = ~a4878 & ~a4876;
assign a4882 = a4880 & ~i308;
assign a4884 = ~a4880 & i308;
assign a4886 = ~a4884 & ~a4882;
assign a4888 = a4886 & a4874;
assign a4890 = a4566 & ~l662;
assign a4892 = ~a4566 & ~l922;
assign a4894 = ~a4892 & ~a4890;
assign a4896 = a4894 & ~i310;
assign a4898 = ~a4894 & i310;
assign a4900 = ~a4898 & ~a4896;
assign a4902 = a4900 & a4888;
assign a4904 = a4566 & ~l668;
assign a4906 = ~a4566 & ~l924;
assign a4908 = ~a4906 & ~a4904;
assign a4910 = a4908 & ~i312;
assign a4912 = ~a4908 & i312;
assign a4914 = ~a4912 & ~a4910;
assign a4916 = a4914 & a4902;
assign a4918 = ~a4566 & ~l926;
assign a4920 = a4566 & l670;
assign a4922 = ~a4920 & ~a4918;
assign a4924 = a4922 & ~i314;
assign a4926 = ~a4922 & i314;
assign a4928 = ~a4926 & ~a4924;
assign a4930 = a4928 & a4916;
assign a4932 = a4566 & ~l674;
assign a4934 = ~a4566 & ~l928;
assign a4936 = ~a4934 & ~a4932;
assign a4938 = a4936 & ~i316;
assign a4940 = ~a4936 & i316;
assign a4942 = ~a4940 & ~a4938;
assign a4944 = a4942 & a4930;
assign a4946 = ~a4566 & ~l930;
assign a4948 = a4566 & l676;
assign a4950 = ~a4948 & ~a4946;
assign a4952 = a4950 & ~i318;
assign a4954 = ~a4950 & i318;
assign a4956 = ~a4954 & ~a4952;
assign a4958 = a4956 & a4944;
assign a4960 = a4566 & ~l682;
assign a4962 = ~a4566 & ~l932;
assign a4964 = ~a4962 & ~a4960;
assign a4966 = a4964 & ~i320;
assign a4968 = ~a4964 & i320;
assign a4970 = ~a4968 & ~a4966;
assign a4972 = a4970 & a4958;
assign a4974 = ~a4566 & ~l934;
assign a4976 = a4566 & l684;
assign a4978 = ~a4976 & ~a4974;
assign a4980 = a4978 & ~i322;
assign a4982 = ~a4978 & i322;
assign a4984 = ~a4982 & ~a4980;
assign a4986 = a4984 & a4972;
assign a4988 = a4566 & ~l688;
assign a4990 = ~a4566 & ~l936;
assign a4992 = ~a4990 & ~a4988;
assign a4994 = a4992 & ~i324;
assign a4996 = ~a4992 & i324;
assign a4998 = ~a4996 & ~a4994;
assign a5000 = a4998 & a4986;
assign a5002 = ~a4566 & ~l938;
assign a5004 = a4566 & l690;
assign a5006 = ~a5004 & ~a5002;
assign a5008 = a5006 & ~i326;
assign a5010 = ~a5006 & i326;
assign a5012 = ~a5010 & ~a5008;
assign a5014 = a5012 & a5000;
assign a5016 = a4566 & ~l696;
assign a5018 = ~a4566 & ~l940;
assign a5020 = ~a5018 & ~a5016;
assign a5022 = a5020 & ~i328;
assign a5024 = ~a5020 & i328;
assign a5026 = ~a5024 & ~a5022;
assign a5028 = a5026 & a5014;
assign a5030 = ~a4566 & ~l942;
assign a5032 = a4566 & l698;
assign a5034 = ~a5032 & ~a5030;
assign a5036 = a5034 & ~i330;
assign a5038 = ~a5034 & i330;
assign a5040 = ~a5038 & ~a5036;
assign a5042 = a5040 & a5028;
assign a5044 = a4566 & ~l702;
assign a5046 = ~a4566 & ~l944;
assign a5048 = ~a5046 & ~a5044;
assign a5050 = a5048 & ~i332;
assign a5052 = ~a5048 & i332;
assign a5054 = ~a5052 & ~a5050;
assign a5056 = a5054 & a5042;
assign a5058 = ~a4566 & ~l946;
assign a5060 = a4566 & l704;
assign a5062 = ~a5060 & ~a5058;
assign a5064 = a5062 & ~i334;
assign a5066 = ~a5062 & i334;
assign a5068 = ~a5066 & ~a5064;
assign a5070 = a5068 & a5056;
assign a5072 = a4566 & ~l706;
assign a5074 = ~a4566 & ~l948;
assign a5076 = ~a5074 & ~a5072;
assign a5078 = a5076 & ~i336;
assign a5080 = ~a5076 & i336;
assign a5082 = ~a5080 & ~a5078;
assign a5084 = a5082 & a5070;
assign a5086 = a4566 & ~l708;
assign a5088 = ~a4566 & ~l950;
assign a5090 = ~a5088 & ~a5086;
assign a5092 = a5090 & ~i338;
assign a5094 = ~a5090 & i338;
assign a5096 = ~a5094 & ~a5092;
assign a5098 = a5096 & a5084;
assign a5100 = ~a4566 & ~l952;
assign a5102 = a4566 & l710;
assign a5104 = ~a5102 & ~a5100;
assign a5106 = a5104 & ~i340;
assign a5108 = ~a5104 & i340;
assign a5110 = ~a5108 & ~a5106;
assign a5112 = a5110 & a5098;
assign a5114 = a4566 & ~l712;
assign a5116 = ~a4566 & ~l954;
assign a5118 = ~a5116 & ~a5114;
assign a5120 = a5118 & ~i342;
assign a5122 = ~a5118 & i342;
assign a5124 = ~a5122 & ~a5120;
assign a5126 = a5124 & a5112;
assign a5128 = a4566 & ~l714;
assign a5130 = ~a4566 & ~l956;
assign a5132 = ~a5130 & ~a5128;
assign a5134 = a5132 & ~i344;
assign a5136 = ~a5132 & i344;
assign a5138 = ~a5136 & ~a5134;
assign a5140 = a5138 & a5126;
assign a5142 = a4566 & ~l716;
assign a5144 = ~a4566 & ~l958;
assign a5146 = ~a5144 & ~a5142;
assign a5148 = a5146 & ~i346;
assign a5150 = ~a5146 & i346;
assign a5152 = ~a5150 & ~a5148;
assign a5154 = a5152 & a5140;
assign a5156 = a4566 & ~l720;
assign a5158 = ~a4566 & ~l960;
assign a5160 = ~a5158 & ~a5156;
assign a5162 = a5160 & ~i348;
assign a5164 = ~a5160 & i348;
assign a5166 = ~a5164 & ~a5162;
assign a5168 = a5166 & a5154;
assign a5170 = a4566 & ~l722;
assign a5172 = ~a4566 & ~l962;
assign a5174 = ~a5172 & ~a5170;
assign a5176 = a5174 & ~i350;
assign a5178 = ~a5174 & i350;
assign a5180 = ~a5178 & ~a5176;
assign a5182 = a5180 & a5168;
assign a5184 = a4566 & ~l724;
assign a5186 = ~a4566 & ~l964;
assign a5188 = ~a5186 & ~a5184;
assign a5190 = a5188 & ~i352;
assign a5192 = ~a5188 & i352;
assign a5194 = ~a5192 & ~a5190;
assign a5196 = a5194 & a5182;
assign a5198 = a4566 & ~l726;
assign a5200 = ~a4566 & ~l966;
assign a5202 = ~a5200 & ~a5198;
assign a5204 = a5202 & ~i354;
assign a5206 = ~a5202 & i354;
assign a5208 = ~a5206 & ~a5204;
assign a5210 = a5208 & a5196;
assign a5212 = a4566 & ~l728;
assign a5214 = ~a4566 & ~l968;
assign a5216 = ~a5214 & ~a5212;
assign a5218 = a5216 & ~i356;
assign a5220 = ~a5216 & i356;
assign a5222 = ~a5220 & ~a5218;
assign a5224 = a5222 & a5210;
assign a5226 = a4566 & ~l730;
assign a5228 = ~a4566 & ~l970;
assign a5230 = ~a5228 & ~a5226;
assign a5232 = a5230 & ~i358;
assign a5234 = ~a5230 & i358;
assign a5236 = ~a5234 & ~a5232;
assign a5238 = a5236 & a5224;
assign a5240 = a4566 & ~l736;
assign a5242 = ~a4566 & ~l972;
assign a5244 = ~a5242 & ~a5240;
assign a5246 = a5244 & ~i360;
assign a5248 = ~a5244 & i360;
assign a5250 = ~a5248 & ~a5246;
assign a5252 = a5250 & a5238;
assign a5254 = ~a4566 & ~l974;
assign a5256 = a4566 & l738;
assign a5258 = ~a5256 & ~a5254;
assign a5260 = a5258 & ~i362;
assign a5262 = ~a5258 & i362;
assign a5264 = ~a5262 & ~a5260;
assign a5266 = a5264 & a5252;
assign a5268 = a4566 & ~l742;
assign a5270 = ~a4566 & ~l976;
assign a5272 = ~a5270 & ~a5268;
assign a5274 = a5272 & ~i364;
assign a5276 = ~a5272 & i364;
assign a5278 = ~a5276 & ~a5274;
assign a5280 = a5278 & a5266;
assign a5282 = ~a4566 & ~l978;
assign a5284 = a4566 & l744;
assign a5286 = ~a5284 & ~a5282;
assign a5288 = a5286 & ~i366;
assign a5290 = ~a5286 & i366;
assign a5292 = ~a5290 & ~a5288;
assign a5294 = a5292 & a5280;
assign a5296 = a4566 & ~l750;
assign a5298 = ~a4566 & ~l980;
assign a5300 = ~a5298 & ~a5296;
assign a5302 = a5300 & ~i368;
assign a5304 = ~a5300 & i368;
assign a5306 = ~a5304 & ~a5302;
assign a5308 = a5306 & a5294;
assign a5310 = ~a4566 & ~l982;
assign a5312 = a4566 & l752;
assign a5314 = ~a5312 & ~a5310;
assign a5316 = a5314 & ~i370;
assign a5318 = ~a5314 & i370;
assign a5320 = ~a5318 & ~a5316;
assign a5322 = a5320 & a5308;
assign a5324 = a4566 & ~l756;
assign a5326 = ~a4566 & ~l984;
assign a5328 = ~a5326 & ~a5324;
assign a5330 = a5328 & ~i372;
assign a5332 = ~a5328 & i372;
assign a5334 = ~a5332 & ~a5330;
assign a5336 = a5334 & a5322;
assign a5338 = ~a4566 & ~l986;
assign a5340 = a4566 & l758;
assign a5342 = ~a5340 & ~a5338;
assign a5344 = a5342 & ~i374;
assign a5346 = ~a5342 & i374;
assign a5348 = ~a5346 & ~a5344;
assign a5350 = a5348 & a5336;
assign a5352 = a4566 & ~l764;
assign a5354 = ~a4566 & ~l988;
assign a5356 = ~a5354 & ~a5352;
assign a5358 = a5356 & ~i376;
assign a5360 = ~a5356 & i376;
assign a5362 = ~a5360 & ~a5358;
assign a5364 = a5362 & a5350;
assign a5366 = ~a4566 & ~l990;
assign a5368 = a4566 & l766;
assign a5370 = ~a5368 & ~a5366;
assign a5372 = a5370 & ~i378;
assign a5374 = ~a5370 & i378;
assign a5376 = ~a5374 & ~a5372;
assign a5378 = a5376 & a5364;
assign a5380 = a4566 & ~l770;
assign a5382 = ~a4566 & ~l992;
assign a5384 = ~a5382 & ~a5380;
assign a5386 = a5384 & ~i380;
assign a5388 = ~a5384 & i380;
assign a5390 = ~a5388 & ~a5386;
assign a5392 = a5390 & a5378;
assign a5394 = ~a4566 & ~l994;
assign a5396 = a4566 & l772;
assign a5398 = ~a5396 & ~a5394;
assign a5400 = a5398 & ~i382;
assign a5402 = ~a5398 & i382;
assign a5404 = ~a5402 & ~a5400;
assign a5406 = a5404 & a5392;
assign a5408 = a4566 & ~l774;
assign a5410 = ~a4566 & ~l996;
assign a5412 = ~a5410 & ~a5408;
assign a5414 = a5412 & ~i384;
assign a5416 = ~a5412 & i384;
assign a5418 = ~a5416 & ~a5414;
assign a5420 = a5418 & a5406;
assign a5422 = a4566 & ~l776;
assign a5424 = ~a4566 & ~l998;
assign a5426 = ~a5424 & ~a5422;
assign a5428 = a5426 & ~i386;
assign a5430 = ~a5426 & i386;
assign a5432 = ~a5430 & ~a5428;
assign a5434 = a5432 & a5420;
assign a5436 = ~a4566 & ~l1000;
assign a5438 = a4566 & l778;
assign a5440 = ~a5438 & ~a5436;
assign a5442 = a5440 & ~i388;
assign a5444 = ~a5440 & i388;
assign a5446 = ~a5444 & ~a5442;
assign a5448 = a5446 & a5434;
assign a5450 = a4566 & ~l780;
assign a5452 = ~a4566 & ~l1002;
assign a5454 = ~a5452 & ~a5450;
assign a5456 = a5454 & ~i390;
assign a5458 = ~a5454 & i390;
assign a5460 = ~a5458 & ~a5456;
assign a5462 = a5460 & a5448;
assign a5464 = a4566 & ~l782;
assign a5466 = ~a4566 & ~l1004;
assign a5468 = ~a5466 & ~a5464;
assign a5470 = a5468 & ~i392;
assign a5472 = ~a5468 & i392;
assign a5474 = ~a5472 & ~a5470;
assign a5476 = a5474 & a5462;
assign a5478 = a4566 & ~l784;
assign a5480 = ~a4566 & ~l1006;
assign a5482 = ~a5480 & ~a5478;
assign a5484 = a5482 & ~i394;
assign a5486 = ~a5482 & i394;
assign a5488 = ~a5486 & ~a5484;
assign a5490 = a5488 & a5476;
assign a5492 = a4566 & ~l788;
assign a5494 = ~a4566 & ~l1008;
assign a5496 = ~a5494 & ~a5492;
assign a5498 = a5496 & ~i396;
assign a5500 = ~a5496 & i396;
assign a5502 = ~a5500 & ~a5498;
assign a5504 = a5502 & a5490;
assign a5506 = a4566 & ~l790;
assign a5508 = ~a4566 & ~l1010;
assign a5510 = ~a5508 & ~a5506;
assign a5512 = a5510 & ~i398;
assign a5514 = ~a5510 & i398;
assign a5516 = ~a5514 & ~a5512;
assign a5518 = a5516 & a5504;
assign a5520 = a4566 & ~l792;
assign a5522 = ~a4566 & ~l1012;
assign a5524 = ~a5522 & ~a5520;
assign a5526 = a5524 & ~i400;
assign a5528 = ~a5524 & i400;
assign a5530 = ~a5528 & ~a5526;
assign a5532 = a5530 & a5518;
assign a5534 = a4566 & ~l794;
assign a5536 = ~a4566 & ~l1014;
assign a5538 = ~a5536 & ~a5534;
assign a5540 = a5538 & ~i402;
assign a5542 = ~a5538 & i402;
assign a5544 = ~a5542 & ~a5540;
assign a5546 = a5544 & a5532;
assign a5548 = a4566 & ~l796;
assign a5550 = ~a4566 & ~l1016;
assign a5552 = ~a5550 & ~a5548;
assign a5554 = a5552 & ~i404;
assign a5556 = ~a5552 & i404;
assign a5558 = ~a5556 & ~a5554;
assign a5560 = a5558 & a5546;
assign a5562 = a4566 & ~l798;
assign a5564 = ~a4566 & ~l1018;
assign a5566 = ~a5564 & ~a5562;
assign a5568 = a5566 & ~i406;
assign a5570 = ~a5566 & i406;
assign a5572 = ~a5570 & ~a5568;
assign a5574 = a5572 & a5560;
assign a5576 = a4566 & ~l804;
assign a5578 = ~a4566 & ~l1020;
assign a5580 = ~a5578 & ~a5576;
assign a5582 = a5580 & ~i408;
assign a5584 = ~a5580 & i408;
assign a5586 = ~a5584 & ~a5582;
assign a5588 = a5586 & a5574;
assign a5590 = ~a4566 & ~l1022;
assign a5592 = a4566 & l806;
assign a5594 = ~a5592 & ~a5590;
assign a5596 = a5594 & ~i410;
assign a5598 = ~a5594 & i410;
assign a5600 = ~a5598 & ~a5596;
assign a5602 = a5600 & a5588;
assign a5604 = a4566 & ~l810;
assign a5606 = ~a4566 & ~l1024;
assign a5608 = ~a5606 & ~a5604;
assign a5610 = a5608 & ~i412;
assign a5612 = ~a5608 & i412;
assign a5614 = ~a5612 & ~a5610;
assign a5616 = a5614 & a5602;
assign a5618 = ~a4566 & ~l1026;
assign a5620 = a4566 & l812;
assign a5622 = ~a5620 & ~a5618;
assign a5624 = a5622 & ~i414;
assign a5626 = ~a5622 & i414;
assign a5628 = ~a5626 & ~a5624;
assign a5630 = a5628 & a5616;
assign a5632 = a4566 & ~l818;
assign a5634 = ~a4566 & ~l1028;
assign a5636 = ~a5634 & ~a5632;
assign a5638 = a5636 & ~i416;
assign a5640 = ~a5636 & i416;
assign a5642 = ~a5640 & ~a5638;
assign a5644 = a5642 & a5630;
assign a5646 = ~a4566 & ~l1030;
assign a5648 = a4566 & l820;
assign a5650 = ~a5648 & ~a5646;
assign a5652 = a5650 & ~i418;
assign a5654 = ~a5650 & i418;
assign a5656 = ~a5654 & ~a5652;
assign a5658 = a5656 & a5644;
assign a5660 = a4566 & ~l824;
assign a5662 = ~a4566 & ~l1032;
assign a5664 = ~a5662 & ~a5660;
assign a5666 = a5664 & ~i420;
assign a5668 = ~a5664 & i420;
assign a5670 = ~a5668 & ~a5666;
assign a5672 = a5670 & a5658;
assign a5674 = ~a4566 & ~l1034;
assign a5676 = a4566 & l826;
assign a5678 = ~a5676 & ~a5674;
assign a5680 = a5678 & ~i422;
assign a5682 = ~a5678 & i422;
assign a5684 = ~a5682 & ~a5680;
assign a5686 = a5684 & a5672;
assign a5688 = a4566 & ~l832;
assign a5690 = ~a4566 & ~l1036;
assign a5692 = ~a5690 & ~a5688;
assign a5694 = a5692 & ~i424;
assign a5696 = ~a5692 & i424;
assign a5698 = ~a5696 & ~a5694;
assign a5700 = a5698 & a5686;
assign a5702 = ~a4566 & ~l1038;
assign a5704 = a4566 & l834;
assign a5706 = ~a5704 & ~a5702;
assign a5708 = a5706 & ~i426;
assign a5710 = ~a5706 & i426;
assign a5712 = ~a5710 & ~a5708;
assign a5714 = a5712 & a5700;
assign a5716 = a4566 & ~l838;
assign a5718 = ~a4566 & ~l1040;
assign a5720 = ~a5718 & ~a5716;
assign a5722 = a5720 & ~i428;
assign a5724 = ~a5720 & i428;
assign a5726 = ~a5724 & ~a5722;
assign a5728 = a5726 & a5714;
assign a5730 = ~a4566 & ~l1042;
assign a5732 = a4566 & l840;
assign a5734 = ~a5732 & ~a5730;
assign a5736 = a5734 & ~i430;
assign a5738 = ~a5734 & i430;
assign a5740 = ~a5738 & ~a5736;
assign a5742 = a5740 & a5728;
assign a5744 = a4566 & ~l842;
assign a5746 = ~a4566 & ~l1044;
assign a5748 = ~a5746 & ~a5744;
assign a5750 = a5748 & ~i432;
assign a5752 = ~a5748 & i432;
assign a5754 = ~a5752 & ~a5750;
assign a5756 = a5754 & a5742;
assign a5758 = a4566 & ~l844;
assign a5760 = ~a4566 & ~l1046;
assign a5762 = ~a5760 & ~a5758;
assign a5764 = a5762 & ~i434;
assign a5766 = ~a5762 & i434;
assign a5768 = ~a5766 & ~a5764;
assign a5770 = a5768 & a5756;
assign a5772 = ~a4566 & ~l1048;
assign a5774 = a4566 & l846;
assign a5776 = ~a5774 & ~a5772;
assign a5778 = a5776 & ~i436;
assign a5780 = ~a5776 & i436;
assign a5782 = ~a5780 & ~a5778;
assign a5784 = a5782 & a5770;
assign a5786 = a4566 & ~l848;
assign a5788 = ~a4566 & ~l1050;
assign a5790 = ~a5788 & ~a5786;
assign a5792 = a5790 & ~i438;
assign a5794 = ~a5790 & i438;
assign a5796 = ~a5794 & ~a5792;
assign a5798 = a5796 & a5784;
assign a5800 = a4566 & ~l850;
assign a5802 = ~a4566 & ~l1052;
assign a5804 = ~a5802 & ~a5800;
assign a5806 = a5804 & ~i440;
assign a5808 = ~a5804 & i440;
assign a5810 = ~a5808 & ~a5806;
assign a5812 = a5810 & a5798;
assign a5814 = a4566 & ~l852;
assign a5816 = ~a4566 & ~l1054;
assign a5818 = ~a5816 & ~a5814;
assign a5820 = a5818 & ~i442;
assign a5822 = ~a5818 & i442;
assign a5824 = ~a5822 & ~a5820;
assign a5826 = a5824 & a5812;
assign a5828 = a4566 & ~l856;
assign a5830 = ~a4566 & ~l1056;
assign a5832 = ~a5830 & ~a5828;
assign a5834 = a5832 & ~i444;
assign a5836 = ~a5832 & i444;
assign a5838 = ~a5836 & ~a5834;
assign a5840 = a5838 & a5826;
assign a5842 = a4566 & ~l858;
assign a5844 = ~a4566 & ~l1058;
assign a5846 = ~a5844 & ~a5842;
assign a5848 = a5846 & ~i446;
assign a5850 = ~a5846 & i446;
assign a5852 = ~a5850 & ~a5848;
assign a5854 = a5852 & a5840;
assign a5856 = a4566 & ~l860;
assign a5858 = ~a4566 & ~l1060;
assign a5860 = ~a5858 & ~a5856;
assign a5862 = a5860 & ~i448;
assign a5864 = ~a5860 & i448;
assign a5866 = ~a5864 & ~a5862;
assign a5868 = a5866 & a5854;
assign a5870 = a4566 & ~l862;
assign a5872 = ~a4566 & ~l1062;
assign a5874 = ~a5872 & ~a5870;
assign a5876 = a5874 & ~i450;
assign a5878 = ~a5874 & i450;
assign a5880 = ~a5878 & ~a5876;
assign a5882 = a5880 & a5868;
assign a5884 = a4566 & ~l864;
assign a5886 = ~a4566 & ~l1064;
assign a5888 = ~a5886 & ~a5884;
assign a5890 = a5888 & ~i452;
assign a5892 = ~a5888 & i452;
assign a5894 = ~a5892 & ~a5890;
assign a5896 = a5894 & a5882;
assign a5898 = a4566 & ~l866;
assign a5900 = ~a4566 & ~l1066;
assign a5902 = ~a5900 & ~a5898;
assign a5904 = a5902 & ~i454;
assign a5906 = ~a5902 & i454;
assign a5908 = ~a5906 & ~a5904;
assign a5910 = a5908 & a5896;
assign a5912 = a4566 & ~l868;
assign a5914 = ~a4566 & ~l1068;
assign a5916 = ~a5914 & ~a5912;
assign a5918 = a5916 & ~i456;
assign a5920 = ~a5916 & i456;
assign a5922 = ~a5920 & ~a5918;
assign a5924 = a5922 & a5910;
assign a5926 = a4566 & ~l870;
assign a5928 = ~a4566 & ~l1070;
assign a5930 = ~a5928 & ~a5926;
assign a5932 = a5930 & ~i458;
assign a5934 = ~a5930 & i458;
assign a5936 = ~a5934 & ~a5932;
assign a5938 = a5936 & a5924;
assign a5940 = a4566 & ~l872;
assign a5942 = ~a4566 & ~l1072;
assign a5944 = ~a5942 & ~a5940;
assign a5946 = a5944 & ~i460;
assign a5948 = ~a5944 & i460;
assign a5950 = ~a5948 & ~a5946;
assign a5952 = a5950 & a5938;
assign a5954 = a4566 & ~l874;
assign a5956 = ~a4566 & ~l1074;
assign a5958 = ~a5956 & ~a5954;
assign a5960 = a5958 & ~i462;
assign a5962 = ~a5958 & i462;
assign a5964 = ~a5962 & ~a5960;
assign a5966 = a5964 & a5952;
assign a5968 = ~l480 & ~l478;
assign a5970 = ~a5968 & l476;
assign a5972 = l484 & l482;
assign a5974 = ~l490 & ~l488;
assign a5976 = ~a5974 & l486;
assign a5978 = l494 & l492;
assign a5980 = ~l500 & ~l498;
assign a5982 = ~a5980 & l496;
assign a5984 = l504 & l502;
assign a5986 = ~l510 & ~l508;
assign a5988 = ~a5986 & l506;
assign a5990 = l514 & l512;
assign a5992 = ~l520 & ~l518;
assign a5994 = ~a5992 & l516;
assign a5996 = l524 & l522;
assign a5998 = ~l530 & ~l528;
assign a6000 = ~a5998 & l526;
assign a6002 = l534 & l532;
assign a6004 = ~l540 & ~l538;
assign a6006 = ~a6004 & l536;
assign a6008 = l544 & l542;
assign a6010 = ~l550 & ~l548;
assign a6012 = ~a6010 & l546;
assign a6014 = l554 & l552;
assign a6016 = ~l560 & ~l558;
assign a6018 = ~a6016 & l556;
assign a6020 = l564 & l562;
assign a6022 = ~l570 & ~l568;
assign a6024 = ~a6022 & l566;
assign a6026 = l574 & l572;
assign a6028 = ~l580 & ~l578;
assign a6030 = ~a6028 & l576;
assign a6032 = l584 & l582;
assign a6034 = ~l590 & ~l588;
assign a6036 = ~a6034 & l586;
assign a6038 = l594 & l592;
assign a6040 = l598 & l596;
assign a6042 = ~l602 & l600;
assign a6044 = l612 & l610;
assign a6046 = ~l616 & l614;
assign a6048 = l626 & l624;
assign a6050 = ~l630 & l628;
assign a6052 = a1182 & l638;
assign a6054 = l648 & l646;
assign a6056 = a1534 & l656;
assign a6058 = l666 & l664;
assign a6060 = ~l670 & l668;
assign a6062 = l680 & l678;
assign a6064 = ~l684 & l682;
assign a6066 = l694 & l692;
assign a6068 = ~l698 & l696;
assign a6070 = a1774 & l706;
assign a6072 = l716 & l714;
assign a6074 = a2126 & l724;
assign a6076 = l734 & l732;
assign a6078 = ~l738 & l736;
assign a6080 = l748 & l746;
assign a6082 = ~l752 & l750;
assign a6084 = l762 & l760;
assign a6086 = ~l766 & l764;
assign a6088 = a2366 & l774;
assign a6090 = l784 & l782;
assign a6092 = a2718 & l792;
assign a6094 = l802 & l800;
assign a6096 = ~l806 & l804;
assign a6098 = l816 & l814;
assign a6100 = ~l820 & l818;
assign a6102 = l830 & l828;
assign a6104 = ~l834 & l832;
assign a6106 = a2958 & l842;
assign a6108 = l852 & l850;
assign a6110 = a3310 & l860;
assign a6112 = l878 & l876;
assign a6114 = l886 & l884;
assign a6116 = l894 & l892;
assign a6118 = l904 & l902;
assign a6120 = a6118 & l900;
assign a6122 = l910 & l908;
assign a6124 = l920 & l918;
assign a6126 = a6124 & l916;
assign a6128 = l926 & l924;
assign a6130 = l934 & l932;
assign a6132 = l942 & l940;
assign a6134 = l952 & l950;
assign a6136 = a6134 & l948;
assign a6138 = l958 & l956;
assign a6140 = l968 & l966;
assign a6142 = a6140 & l964;
assign a6144 = l974 & l972;
assign a6146 = l982 & l980;
assign a6148 = l990 & l988;
assign a6150 = l1000 & l998;
assign a6152 = a6150 & l996;
assign a6154 = l1006 & l1004;
assign a6156 = l1016 & l1014;
assign a6158 = a6156 & l1012;
assign a6160 = l1022 & l1020;
assign a6162 = l1030 & l1028;
assign a6164 = l1038 & l1036;
assign a6166 = l1048 & l1046;
assign a6168 = a6166 & l1044;
assign a6170 = l1054 & l1052;
assign a6172 = l1064 & l1062;
assign a6174 = a6172 & l1060;
assign a6176 = ~l788 & ~l720;
assign a6178 = l788 & l720;
assign a6180 = ~a6178 & ~a6176;
assign a6182 = a2296 & a1704;
assign a6184 = a6182 & ~a6180;
assign a6186 = ~l720 & ~l652;
assign a6188 = l720 & l652;
assign a6190 = ~a6188 & ~a6186;
assign a6192 = ~a6190 & a1704;
assign a6194 = ~l788 & ~l652;
assign a6196 = l788 & l652;
assign a6198 = ~a6196 & ~a6194;
assign a6200 = ~a6198 & a2296;
assign a6202 = ~l856 & ~l652;
assign a6204 = l856 & l652;
assign a6206 = ~a6204 & ~a6202;
assign a6208 = ~a6206 & a2888;
assign a6210 = ~a6208 & ~a6200;
assign a6212 = a6210 & ~a6192;
assign a6214 = ~a6212 & a1112;
assign a6216 = ~l856 & ~l720;
assign a6218 = l856 & l720;
assign a6220 = ~a6218 & ~a6216;
assign a6222 = a2888 & a1704;
assign a6224 = a6222 & ~a6220;
assign a6226 = ~l856 & ~l788;
assign a6228 = l856 & l788;
assign a6230 = ~a6228 & ~a6226;
assign a6232 = a2888 & a2296;
assign a6234 = a6232 & ~a6230;
assign a6236 = ~a6234 & ~a6224;
assign a6238 = a6236 & ~a6214;
assign a6240 = a6238 & ~a6184;
assign a6242 = ~a6240 & l868;
assign a6244 = a5968 & ~l476;
assign a6246 = l480 & ~l478;
assign a6248 = a6246 & ~l476;
assign a6250 = ~l480 & l478;
assign a6252 = a6250 & ~l476;
assign a6254 = l480 & l478;
assign a6256 = a6254 & ~l476;
assign a6258 = a5968 & l476;
assign a6260 = ~l804 & ~l484;
assign a6262 = ~l818 & l484;
assign a6264 = ~a6262 & ~a6260;
assign a6266 = ~a6264 & ~l482;
assign a6268 = ~l484 & l482;
assign a6270 = a6268 & ~l832;
assign a6272 = ~a6270 & ~a6266;
assign a6274 = ~a6272 & a6258;
assign a6276 = a6274 & ~a6256;
assign a6278 = ~l736 & ~l484;
assign a6280 = ~l750 & l484;
assign a6282 = ~a6280 & ~a6278;
assign a6284 = ~a6282 & ~l482;
assign a6286 = a6268 & ~l764;
assign a6288 = ~a6286 & ~a6284;
assign a6290 = ~a6288 & a6256;
assign a6292 = ~a6290 & ~a6276;
assign a6294 = ~a6292 & ~a6252;
assign a6296 = ~l668 & ~l484;
assign a6298 = ~l682 & l484;
assign a6300 = ~a6298 & ~a6296;
assign a6302 = ~a6300 & ~l482;
assign a6304 = a6268 & ~l696;
assign a6306 = ~a6304 & ~a6302;
assign a6308 = ~a6306 & a6252;
assign a6310 = ~a6308 & ~a6294;
assign a6312 = ~a6310 & ~a6248;
assign a6314 = ~l600 & ~l484;
assign a6316 = ~l614 & l484;
assign a6318 = ~a6316 & ~a6314;
assign a6320 = ~a6318 & ~l482;
assign a6322 = a6268 & ~l628;
assign a6324 = ~a6322 & ~a6320;
assign a6326 = ~a6324 & a6248;
assign a6328 = ~a6326 & ~a6312;
assign a6330 = a6328 & ~l596;
assign a6332 = ~a6328 & l596;
assign a6334 = ~a6332 & ~a6330;
assign a6336 = l806 & ~l484;
assign a6338 = l820 & l484;
assign a6340 = ~a6338 & ~a6336;
assign a6342 = ~a6340 & ~l482;
assign a6344 = a6268 & l834;
assign a6346 = ~a6344 & ~a6342;
assign a6348 = ~a6346 & a6258;
assign a6350 = a6348 & ~a6256;
assign a6352 = l738 & ~l484;
assign a6354 = l752 & l484;
assign a6356 = ~a6354 & ~a6352;
assign a6358 = ~a6356 & ~l482;
assign a6360 = a6268 & l766;
assign a6362 = ~a6360 & ~a6358;
assign a6364 = ~a6362 & a6256;
assign a6366 = ~a6364 & ~a6350;
assign a6368 = ~a6366 & ~a6252;
assign a6370 = l670 & ~l484;
assign a6372 = l684 & l484;
assign a6374 = ~a6372 & ~a6370;
assign a6376 = ~a6374 & ~l482;
assign a6378 = a6268 & l698;
assign a6380 = ~a6378 & ~a6376;
assign a6382 = ~a6380 & a6252;
assign a6384 = ~a6382 & ~a6368;
assign a6386 = ~a6384 & ~a6248;
assign a6388 = l602 & ~l484;
assign a6390 = l616 & l484;
assign a6392 = ~a6390 & ~a6388;
assign a6394 = ~a6392 & ~l482;
assign a6396 = a6268 & l630;
assign a6398 = ~a6396 & ~a6394;
assign a6400 = ~a6398 & a6248;
assign a6402 = ~a6400 & ~a6386;
assign a6404 = a6402 & ~l598;
assign a6406 = ~a6402 & l598;
assign a6408 = ~a6406 & ~a6404;
assign a6410 = a6408 & a6334;
assign a6412 = ~a6410 & ~a6244;
assign a6414 = a5974 & ~l486;
assign a6416 = l490 & ~l488;
assign a6418 = a6416 & ~l486;
assign a6420 = ~l490 & l488;
assign a6422 = a6420 & ~l486;
assign a6424 = l490 & l488;
assign a6426 = a6424 & ~l486;
assign a6428 = a5974 & l486;
assign a6430 = ~l804 & ~l494;
assign a6432 = ~l818 & l494;
assign a6434 = ~a6432 & ~a6430;
assign a6436 = ~a6434 & ~l492;
assign a6438 = ~l494 & l492;
assign a6440 = a6438 & ~l832;
assign a6442 = ~a6440 & ~a6436;
assign a6444 = ~a6442 & a6428;
assign a6446 = a6444 & ~a6426;
assign a6448 = ~l736 & ~l494;
assign a6450 = ~l750 & l494;
assign a6452 = ~a6450 & ~a6448;
assign a6454 = ~a6452 & ~l492;
assign a6456 = a6438 & ~l764;
assign a6458 = ~a6456 & ~a6454;
assign a6460 = ~a6458 & a6426;
assign a6462 = ~a6460 & ~a6446;
assign a6464 = ~a6462 & ~a6422;
assign a6466 = ~l668 & ~l494;
assign a6468 = ~l682 & l494;
assign a6470 = ~a6468 & ~a6466;
assign a6472 = ~a6470 & ~l492;
assign a6474 = a6438 & ~l696;
assign a6476 = ~a6474 & ~a6472;
assign a6478 = ~a6476 & a6422;
assign a6480 = ~a6478 & ~a6464;
assign a6482 = ~a6480 & ~a6418;
assign a6484 = ~l600 & ~l494;
assign a6486 = ~l614 & l494;
assign a6488 = ~a6486 & ~a6484;
assign a6490 = ~a6488 & ~l492;
assign a6492 = a6438 & ~l628;
assign a6494 = ~a6492 & ~a6490;
assign a6496 = ~a6494 & a6418;
assign a6498 = ~a6496 & ~a6482;
assign a6500 = a6498 & ~l610;
assign a6502 = ~a6498 & l610;
assign a6504 = ~a6502 & ~a6500;
assign a6506 = l806 & ~l494;
assign a6508 = l820 & l494;
assign a6510 = ~a6508 & ~a6506;
assign a6512 = ~a6510 & ~l492;
assign a6514 = a6438 & l834;
assign a6516 = ~a6514 & ~a6512;
assign a6518 = ~a6516 & a6428;
assign a6520 = a6518 & ~a6426;
assign a6522 = l738 & ~l494;
assign a6524 = l752 & l494;
assign a6526 = ~a6524 & ~a6522;
assign a6528 = ~a6526 & ~l492;
assign a6530 = a6438 & l766;
assign a6532 = ~a6530 & ~a6528;
assign a6534 = ~a6532 & a6426;
assign a6536 = ~a6534 & ~a6520;
assign a6538 = ~a6536 & ~a6422;
assign a6540 = l670 & ~l494;
assign a6542 = l684 & l494;
assign a6544 = ~a6542 & ~a6540;
assign a6546 = ~a6544 & ~l492;
assign a6548 = a6438 & l698;
assign a6550 = ~a6548 & ~a6546;
assign a6552 = ~a6550 & a6422;
assign a6554 = ~a6552 & ~a6538;
assign a6556 = ~a6554 & ~a6418;
assign a6558 = l602 & ~l494;
assign a6560 = l616 & l494;
assign a6562 = ~a6560 & ~a6558;
assign a6564 = ~a6562 & ~l492;
assign a6566 = a6438 & l630;
assign a6568 = ~a6566 & ~a6564;
assign a6570 = ~a6568 & a6418;
assign a6572 = ~a6570 & ~a6556;
assign a6574 = a6572 & ~l612;
assign a6576 = ~a6572 & l612;
assign a6578 = ~a6576 & ~a6574;
assign a6580 = a6578 & a6504;
assign a6582 = ~a6580 & ~a6414;
assign a6584 = a5980 & ~l496;
assign a6586 = l500 & ~l498;
assign a6588 = a6586 & ~l496;
assign a6590 = ~l500 & l498;
assign a6592 = a6590 & ~l496;
assign a6594 = l500 & l498;
assign a6596 = a6594 & ~l496;
assign a6598 = a5980 & l496;
assign a6600 = ~l804 & ~l504;
assign a6602 = ~l818 & l504;
assign a6604 = ~a6602 & ~a6600;
assign a6606 = ~a6604 & ~l502;
assign a6608 = ~l504 & l502;
assign a6610 = a6608 & ~l832;
assign a6612 = ~a6610 & ~a6606;
assign a6614 = ~a6612 & a6598;
assign a6616 = a6614 & ~a6596;
assign a6618 = ~l736 & ~l504;
assign a6620 = ~l750 & l504;
assign a6622 = ~a6620 & ~a6618;
assign a6624 = ~a6622 & ~l502;
assign a6626 = a6608 & ~l764;
assign a6628 = ~a6626 & ~a6624;
assign a6630 = ~a6628 & a6596;
assign a6632 = ~a6630 & ~a6616;
assign a6634 = ~a6632 & ~a6592;
assign a6636 = ~l668 & ~l504;
assign a6638 = ~l682 & l504;
assign a6640 = ~a6638 & ~a6636;
assign a6642 = ~a6640 & ~l502;
assign a6644 = a6608 & ~l696;
assign a6646 = ~a6644 & ~a6642;
assign a6648 = ~a6646 & a6592;
assign a6650 = ~a6648 & ~a6634;
assign a6652 = ~a6650 & ~a6588;
assign a6654 = ~l600 & ~l504;
assign a6656 = ~l614 & l504;
assign a6658 = ~a6656 & ~a6654;
assign a6660 = ~a6658 & ~l502;
assign a6662 = a6608 & ~l628;
assign a6664 = ~a6662 & ~a6660;
assign a6666 = ~a6664 & a6588;
assign a6668 = ~a6666 & ~a6652;
assign a6670 = a6668 & ~l624;
assign a6672 = ~a6668 & l624;
assign a6674 = ~a6672 & ~a6670;
assign a6676 = l806 & ~l504;
assign a6678 = l820 & l504;
assign a6680 = ~a6678 & ~a6676;
assign a6682 = ~a6680 & ~l502;
assign a6684 = a6608 & l834;
assign a6686 = ~a6684 & ~a6682;
assign a6688 = ~a6686 & a6598;
assign a6690 = a6688 & ~a6596;
assign a6692 = l738 & ~l504;
assign a6694 = l752 & l504;
assign a6696 = ~a6694 & ~a6692;
assign a6698 = ~a6696 & ~l502;
assign a6700 = a6608 & l766;
assign a6702 = ~a6700 & ~a6698;
assign a6704 = ~a6702 & a6596;
assign a6706 = ~a6704 & ~a6690;
assign a6708 = ~a6706 & ~a6592;
assign a6710 = l670 & ~l504;
assign a6712 = l684 & l504;
assign a6714 = ~a6712 & ~a6710;
assign a6716 = ~a6714 & ~l502;
assign a6718 = a6608 & l698;
assign a6720 = ~a6718 & ~a6716;
assign a6722 = ~a6720 & a6592;
assign a6724 = ~a6722 & ~a6708;
assign a6726 = ~a6724 & ~a6588;
assign a6728 = l602 & ~l504;
assign a6730 = l616 & l504;
assign a6732 = ~a6730 & ~a6728;
assign a6734 = ~a6732 & ~l502;
assign a6736 = a6608 & l630;
assign a6738 = ~a6736 & ~a6734;
assign a6740 = ~a6738 & a6588;
assign a6742 = ~a6740 & ~a6726;
assign a6744 = a6742 & ~l626;
assign a6746 = ~a6742 & l626;
assign a6748 = ~a6746 & ~a6744;
assign a6750 = a6748 & a6674;
assign a6752 = ~a6750 & ~a6584;
assign a6754 = a5986 & ~l506;
assign a6756 = l510 & ~l508;
assign a6758 = a6756 & ~l506;
assign a6760 = ~l510 & l508;
assign a6762 = a6760 & ~l506;
assign a6764 = l510 & l508;
assign a6766 = a6764 & ~l506;
assign a6768 = a5986 & l506;
assign a6770 = ~l804 & ~l514;
assign a6772 = ~l818 & l514;
assign a6774 = ~a6772 & ~a6770;
assign a6776 = ~a6774 & ~l512;
assign a6778 = ~l514 & l512;
assign a6780 = a6778 & ~l832;
assign a6782 = ~a6780 & ~a6776;
assign a6784 = ~a6782 & a6768;
assign a6786 = a6784 & ~a6766;
assign a6788 = ~l736 & ~l514;
assign a6790 = ~l750 & l514;
assign a6792 = ~a6790 & ~a6788;
assign a6794 = ~a6792 & ~l512;
assign a6796 = a6778 & ~l764;
assign a6798 = ~a6796 & ~a6794;
assign a6800 = ~a6798 & a6766;
assign a6802 = ~a6800 & ~a6786;
assign a6804 = ~a6802 & ~a6762;
assign a6806 = ~l668 & ~l514;
assign a6808 = ~l682 & l514;
assign a6810 = ~a6808 & ~a6806;
assign a6812 = ~a6810 & ~l512;
assign a6814 = a6778 & ~l696;
assign a6816 = ~a6814 & ~a6812;
assign a6818 = ~a6816 & a6762;
assign a6820 = ~a6818 & ~a6804;
assign a6822 = ~a6820 & ~a6758;
assign a6824 = ~l600 & ~l514;
assign a6826 = ~l614 & l514;
assign a6828 = ~a6826 & ~a6824;
assign a6830 = ~a6828 & ~l512;
assign a6832 = a6778 & ~l628;
assign a6834 = ~a6832 & ~a6830;
assign a6836 = ~a6834 & a6758;
assign a6838 = ~a6836 & ~a6822;
assign a6840 = a6838 & ~l664;
assign a6842 = ~a6838 & l664;
assign a6844 = ~a6842 & ~a6840;
assign a6846 = l806 & ~l514;
assign a6848 = l820 & l514;
assign a6850 = ~a6848 & ~a6846;
assign a6852 = ~a6850 & ~l512;
assign a6854 = a6778 & l834;
assign a6856 = ~a6854 & ~a6852;
assign a6858 = ~a6856 & a6768;
assign a6860 = a6858 & ~a6766;
assign a6862 = l738 & ~l514;
assign a6864 = l752 & l514;
assign a6866 = ~a6864 & ~a6862;
assign a6868 = ~a6866 & ~l512;
assign a6870 = a6778 & l766;
assign a6872 = ~a6870 & ~a6868;
assign a6874 = ~a6872 & a6766;
assign a6876 = ~a6874 & ~a6860;
assign a6878 = ~a6876 & ~a6762;
assign a6880 = l670 & ~l514;
assign a6882 = l684 & l514;
assign a6884 = ~a6882 & ~a6880;
assign a6886 = ~a6884 & ~l512;
assign a6888 = a6778 & l698;
assign a6890 = ~a6888 & ~a6886;
assign a6892 = ~a6890 & a6762;
assign a6894 = ~a6892 & ~a6878;
assign a6896 = ~a6894 & ~a6758;
assign a6898 = l602 & ~l514;
assign a6900 = l616 & l514;
assign a6902 = ~a6900 & ~a6898;
assign a6904 = ~a6902 & ~l512;
assign a6906 = a6778 & l630;
assign a6908 = ~a6906 & ~a6904;
assign a6910 = ~a6908 & a6758;
assign a6912 = ~a6910 & ~a6896;
assign a6914 = a6912 & ~l666;
assign a6916 = ~a6912 & l666;
assign a6918 = ~a6916 & ~a6914;
assign a6920 = a6918 & a6844;
assign a6922 = ~a6920 & ~a6754;
assign a6924 = a5992 & ~l516;
assign a6926 = l520 & ~l518;
assign a6928 = a6926 & ~l516;
assign a6930 = ~l520 & l518;
assign a6932 = a6930 & ~l516;
assign a6934 = l520 & l518;
assign a6936 = a6934 & ~l516;
assign a6938 = a5992 & l516;
assign a6940 = ~l804 & ~l524;
assign a6942 = ~l818 & l524;
assign a6944 = ~a6942 & ~a6940;
assign a6946 = ~a6944 & ~l522;
assign a6948 = ~l524 & l522;
assign a6950 = a6948 & ~l832;
assign a6952 = ~a6950 & ~a6946;
assign a6954 = ~a6952 & a6938;
assign a6956 = a6954 & ~a6936;
assign a6958 = ~l736 & ~l524;
assign a6960 = ~l750 & l524;
assign a6962 = ~a6960 & ~a6958;
assign a6964 = ~a6962 & ~l522;
assign a6966 = a6948 & ~l764;
assign a6968 = ~a6966 & ~a6964;
assign a6970 = ~a6968 & a6936;
assign a6972 = ~a6970 & ~a6956;
assign a6974 = ~a6972 & ~a6932;
assign a6976 = ~l668 & ~l524;
assign a6978 = ~l682 & l524;
assign a6980 = ~a6978 & ~a6976;
assign a6982 = ~a6980 & ~l522;
assign a6984 = a6948 & ~l696;
assign a6986 = ~a6984 & ~a6982;
assign a6988 = ~a6986 & a6932;
assign a6990 = ~a6988 & ~a6974;
assign a6992 = ~a6990 & ~a6928;
assign a6994 = ~l600 & ~l524;
assign a6996 = ~l614 & l524;
assign a6998 = ~a6996 & ~a6994;
assign a7000 = ~a6998 & ~l522;
assign a7002 = a6948 & ~l628;
assign a7004 = ~a7002 & ~a7000;
assign a7006 = ~a7004 & a6928;
assign a7008 = ~a7006 & ~a6992;
assign a7010 = a7008 & ~l678;
assign a7012 = ~a7008 & l678;
assign a7014 = ~a7012 & ~a7010;
assign a7016 = l806 & ~l524;
assign a7018 = l820 & l524;
assign a7020 = ~a7018 & ~a7016;
assign a7022 = ~a7020 & ~l522;
assign a7024 = a6948 & l834;
assign a7026 = ~a7024 & ~a7022;
assign a7028 = ~a7026 & a6938;
assign a7030 = a7028 & ~a6936;
assign a7032 = l738 & ~l524;
assign a7034 = l752 & l524;
assign a7036 = ~a7034 & ~a7032;
assign a7038 = ~a7036 & ~l522;
assign a7040 = a6948 & l766;
assign a7042 = ~a7040 & ~a7038;
assign a7044 = ~a7042 & a6936;
assign a7046 = ~a7044 & ~a7030;
assign a7048 = ~a7046 & ~a6932;
assign a7050 = l670 & ~l524;
assign a7052 = l684 & l524;
assign a7054 = ~a7052 & ~a7050;
assign a7056 = ~a7054 & ~l522;
assign a7058 = a6948 & l698;
assign a7060 = ~a7058 & ~a7056;
assign a7062 = ~a7060 & a6932;
assign a7064 = ~a7062 & ~a7048;
assign a7066 = ~a7064 & ~a6928;
assign a7068 = l602 & ~l524;
assign a7070 = l616 & l524;
assign a7072 = ~a7070 & ~a7068;
assign a7074 = ~a7072 & ~l522;
assign a7076 = a6948 & l630;
assign a7078 = ~a7076 & ~a7074;
assign a7080 = ~a7078 & a6928;
assign a7082 = ~a7080 & ~a7066;
assign a7084 = a7082 & ~l680;
assign a7086 = ~a7082 & l680;
assign a7088 = ~a7086 & ~a7084;
assign a7090 = a7088 & a7014;
assign a7092 = ~a7090 & ~a6924;
assign a7094 = a5998 & ~l526;
assign a7096 = l530 & ~l528;
assign a7098 = a7096 & ~l526;
assign a7100 = ~l530 & l528;
assign a7102 = a7100 & ~l526;
assign a7104 = l530 & l528;
assign a7106 = a7104 & ~l526;
assign a7108 = a5998 & l526;
assign a7110 = ~l804 & ~l534;
assign a7112 = ~l818 & l534;
assign a7114 = ~a7112 & ~a7110;
assign a7116 = ~a7114 & ~l532;
assign a7118 = ~l534 & l532;
assign a7120 = a7118 & ~l832;
assign a7122 = ~a7120 & ~a7116;
assign a7124 = ~a7122 & a7108;
assign a7126 = a7124 & ~a7106;
assign a7128 = ~l736 & ~l534;
assign a7130 = ~l750 & l534;
assign a7132 = ~a7130 & ~a7128;
assign a7134 = ~a7132 & ~l532;
assign a7136 = a7118 & ~l764;
assign a7138 = ~a7136 & ~a7134;
assign a7140 = ~a7138 & a7106;
assign a7142 = ~a7140 & ~a7126;
assign a7144 = ~a7142 & ~a7102;
assign a7146 = ~l668 & ~l534;
assign a7148 = ~l682 & l534;
assign a7150 = ~a7148 & ~a7146;
assign a7152 = ~a7150 & ~l532;
assign a7154 = a7118 & ~l696;
assign a7156 = ~a7154 & ~a7152;
assign a7158 = ~a7156 & a7102;
assign a7160 = ~a7158 & ~a7144;
assign a7162 = ~a7160 & ~a7098;
assign a7164 = ~l600 & ~l534;
assign a7166 = ~l614 & l534;
assign a7168 = ~a7166 & ~a7164;
assign a7170 = ~a7168 & ~l532;
assign a7172 = a7118 & ~l628;
assign a7174 = ~a7172 & ~a7170;
assign a7176 = ~a7174 & a7098;
assign a7178 = ~a7176 & ~a7162;
assign a7180 = a7178 & ~l692;
assign a7182 = ~a7178 & l692;
assign a7184 = ~a7182 & ~a7180;
assign a7186 = l806 & ~l534;
assign a7188 = l820 & l534;
assign a7190 = ~a7188 & ~a7186;
assign a7192 = ~a7190 & ~l532;
assign a7194 = a7118 & l834;
assign a7196 = ~a7194 & ~a7192;
assign a7198 = ~a7196 & a7108;
assign a7200 = a7198 & ~a7106;
assign a7202 = l738 & ~l534;
assign a7204 = l752 & l534;
assign a7206 = ~a7204 & ~a7202;
assign a7208 = ~a7206 & ~l532;
assign a7210 = a7118 & l766;
assign a7212 = ~a7210 & ~a7208;
assign a7214 = ~a7212 & a7106;
assign a7216 = ~a7214 & ~a7200;
assign a7218 = ~a7216 & ~a7102;
assign a7220 = l670 & ~l534;
assign a7222 = l684 & l534;
assign a7224 = ~a7222 & ~a7220;
assign a7226 = ~a7224 & ~l532;
assign a7228 = a7118 & l698;
assign a7230 = ~a7228 & ~a7226;
assign a7232 = ~a7230 & a7102;
assign a7234 = ~a7232 & ~a7218;
assign a7236 = ~a7234 & ~a7098;
assign a7238 = l602 & ~l534;
assign a7240 = l616 & l534;
assign a7242 = ~a7240 & ~a7238;
assign a7244 = ~a7242 & ~l532;
assign a7246 = a7118 & l630;
assign a7248 = ~a7246 & ~a7244;
assign a7250 = ~a7248 & a7098;
assign a7252 = ~a7250 & ~a7236;
assign a7254 = a7252 & ~l694;
assign a7256 = ~a7252 & l694;
assign a7258 = ~a7256 & ~a7254;
assign a7260 = a7258 & a7184;
assign a7262 = ~a7260 & ~a7094;
assign a7264 = a6004 & ~l536;
assign a7266 = l540 & ~l538;
assign a7268 = a7266 & ~l536;
assign a7270 = ~l540 & l538;
assign a7272 = a7270 & ~l536;
assign a7274 = l540 & l538;
assign a7276 = a7274 & ~l536;
assign a7278 = a6004 & l536;
assign a7280 = ~l804 & ~l544;
assign a7282 = ~l818 & l544;
assign a7284 = ~a7282 & ~a7280;
assign a7286 = ~a7284 & ~l542;
assign a7288 = ~l544 & l542;
assign a7290 = a7288 & ~l832;
assign a7292 = ~a7290 & ~a7286;
assign a7294 = ~a7292 & a7278;
assign a7296 = a7294 & ~a7276;
assign a7298 = ~l736 & ~l544;
assign a7300 = ~l750 & l544;
assign a7302 = ~a7300 & ~a7298;
assign a7304 = ~a7302 & ~l542;
assign a7306 = a7288 & ~l764;
assign a7308 = ~a7306 & ~a7304;
assign a7310 = ~a7308 & a7276;
assign a7312 = ~a7310 & ~a7296;
assign a7314 = ~a7312 & ~a7272;
assign a7316 = ~l668 & ~l544;
assign a7318 = ~l682 & l544;
assign a7320 = ~a7318 & ~a7316;
assign a7322 = ~a7320 & ~l542;
assign a7324 = a7288 & ~l696;
assign a7326 = ~a7324 & ~a7322;
assign a7328 = ~a7326 & a7272;
assign a7330 = ~a7328 & ~a7314;
assign a7332 = ~a7330 & ~a7268;
assign a7334 = ~l600 & ~l544;
assign a7336 = ~l614 & l544;
assign a7338 = ~a7336 & ~a7334;
assign a7340 = ~a7338 & ~l542;
assign a7342 = a7288 & ~l628;
assign a7344 = ~a7342 & ~a7340;
assign a7346 = ~a7344 & a7268;
assign a7348 = ~a7346 & ~a7332;
assign a7350 = a7348 & ~l732;
assign a7352 = ~a7348 & l732;
assign a7354 = ~a7352 & ~a7350;
assign a7356 = l806 & ~l544;
assign a7358 = l820 & l544;
assign a7360 = ~a7358 & ~a7356;
assign a7362 = ~a7360 & ~l542;
assign a7364 = a7288 & l834;
assign a7366 = ~a7364 & ~a7362;
assign a7368 = ~a7366 & a7278;
assign a7370 = a7368 & ~a7276;
assign a7372 = l738 & ~l544;
assign a7374 = l752 & l544;
assign a7376 = ~a7374 & ~a7372;
assign a7378 = ~a7376 & ~l542;
assign a7380 = a7288 & l766;
assign a7382 = ~a7380 & ~a7378;
assign a7384 = ~a7382 & a7276;
assign a7386 = ~a7384 & ~a7370;
assign a7388 = ~a7386 & ~a7272;
assign a7390 = l670 & ~l544;
assign a7392 = l684 & l544;
assign a7394 = ~a7392 & ~a7390;
assign a7396 = ~a7394 & ~l542;
assign a7398 = a7288 & l698;
assign a7400 = ~a7398 & ~a7396;
assign a7402 = ~a7400 & a7272;
assign a7404 = ~a7402 & ~a7388;
assign a7406 = ~a7404 & ~a7268;
assign a7408 = l602 & ~l544;
assign a7410 = l616 & l544;
assign a7412 = ~a7410 & ~a7408;
assign a7414 = ~a7412 & ~l542;
assign a7416 = a7288 & l630;
assign a7418 = ~a7416 & ~a7414;
assign a7420 = ~a7418 & a7268;
assign a7422 = ~a7420 & ~a7406;
assign a7424 = a7422 & ~l734;
assign a7426 = ~a7422 & l734;
assign a7428 = ~a7426 & ~a7424;
assign a7430 = a7428 & a7354;
assign a7432 = ~a7430 & ~a7264;
assign a7434 = a6010 & ~l546;
assign a7436 = l550 & ~l548;
assign a7438 = a7436 & ~l546;
assign a7440 = ~l550 & l548;
assign a7442 = a7440 & ~l546;
assign a7444 = l550 & l548;
assign a7446 = a7444 & ~l546;
assign a7448 = a6010 & l546;
assign a7450 = ~l804 & ~l554;
assign a7452 = ~l818 & l554;
assign a7454 = ~a7452 & ~a7450;
assign a7456 = ~a7454 & ~l552;
assign a7458 = ~l554 & l552;
assign a7460 = a7458 & ~l832;
assign a7462 = ~a7460 & ~a7456;
assign a7464 = ~a7462 & a7448;
assign a7466 = a7464 & ~a7446;
assign a7468 = ~l736 & ~l554;
assign a7470 = ~l750 & l554;
assign a7472 = ~a7470 & ~a7468;
assign a7474 = ~a7472 & ~l552;
assign a7476 = a7458 & ~l764;
assign a7478 = ~a7476 & ~a7474;
assign a7480 = ~a7478 & a7446;
assign a7482 = ~a7480 & ~a7466;
assign a7484 = ~a7482 & ~a7442;
assign a7486 = ~l668 & ~l554;
assign a7488 = ~l682 & l554;
assign a7490 = ~a7488 & ~a7486;
assign a7492 = ~a7490 & ~l552;
assign a7494 = a7458 & ~l696;
assign a7496 = ~a7494 & ~a7492;
assign a7498 = ~a7496 & a7442;
assign a7500 = ~a7498 & ~a7484;
assign a7502 = ~a7500 & ~a7438;
assign a7504 = ~l600 & ~l554;
assign a7506 = ~l614 & l554;
assign a7508 = ~a7506 & ~a7504;
assign a7510 = ~a7508 & ~l552;
assign a7512 = a7458 & ~l628;
assign a7514 = ~a7512 & ~a7510;
assign a7516 = ~a7514 & a7438;
assign a7518 = ~a7516 & ~a7502;
assign a7520 = a7518 & ~l746;
assign a7522 = ~a7518 & l746;
assign a7524 = ~a7522 & ~a7520;
assign a7526 = l806 & ~l554;
assign a7528 = l820 & l554;
assign a7530 = ~a7528 & ~a7526;
assign a7532 = ~a7530 & ~l552;
assign a7534 = a7458 & l834;
assign a7536 = ~a7534 & ~a7532;
assign a7538 = ~a7536 & a7448;
assign a7540 = a7538 & ~a7446;
assign a7542 = l738 & ~l554;
assign a7544 = l752 & l554;
assign a7546 = ~a7544 & ~a7542;
assign a7548 = ~a7546 & ~l552;
assign a7550 = a7458 & l766;
assign a7552 = ~a7550 & ~a7548;
assign a7554 = ~a7552 & a7446;
assign a7556 = ~a7554 & ~a7540;
assign a7558 = ~a7556 & ~a7442;
assign a7560 = l670 & ~l554;
assign a7562 = l684 & l554;
assign a7564 = ~a7562 & ~a7560;
assign a7566 = ~a7564 & ~l552;
assign a7568 = a7458 & l698;
assign a7570 = ~a7568 & ~a7566;
assign a7572 = ~a7570 & a7442;
assign a7574 = ~a7572 & ~a7558;
assign a7576 = ~a7574 & ~a7438;
assign a7578 = l602 & ~l554;
assign a7580 = l616 & l554;
assign a7582 = ~a7580 & ~a7578;
assign a7584 = ~a7582 & ~l552;
assign a7586 = a7458 & l630;
assign a7588 = ~a7586 & ~a7584;
assign a7590 = ~a7588 & a7438;
assign a7592 = ~a7590 & ~a7576;
assign a7594 = a7592 & ~l748;
assign a7596 = ~a7592 & l748;
assign a7598 = ~a7596 & ~a7594;
assign a7600 = a7598 & a7524;
assign a7602 = ~a7600 & ~a7434;
assign a7604 = a6016 & ~l556;
assign a7606 = l560 & ~l558;
assign a7608 = a7606 & ~l556;
assign a7610 = ~l560 & l558;
assign a7612 = a7610 & ~l556;
assign a7614 = l560 & l558;
assign a7616 = a7614 & ~l556;
assign a7618 = a6016 & l556;
assign a7620 = ~l804 & ~l564;
assign a7622 = ~l818 & l564;
assign a7624 = ~a7622 & ~a7620;
assign a7626 = ~a7624 & ~l562;
assign a7628 = ~l564 & l562;
assign a7630 = a7628 & ~l832;
assign a7632 = ~a7630 & ~a7626;
assign a7634 = ~a7632 & a7618;
assign a7636 = a7634 & ~a7616;
assign a7638 = ~l736 & ~l564;
assign a7640 = ~l750 & l564;
assign a7642 = ~a7640 & ~a7638;
assign a7644 = ~a7642 & ~l562;
assign a7646 = a7628 & ~l764;
assign a7648 = ~a7646 & ~a7644;
assign a7650 = ~a7648 & a7616;
assign a7652 = ~a7650 & ~a7636;
assign a7654 = ~a7652 & ~a7612;
assign a7656 = ~l668 & ~l564;
assign a7658 = ~l682 & l564;
assign a7660 = ~a7658 & ~a7656;
assign a7662 = ~a7660 & ~l562;
assign a7664 = a7628 & ~l696;
assign a7666 = ~a7664 & ~a7662;
assign a7668 = ~a7666 & a7612;
assign a7670 = ~a7668 & ~a7654;
assign a7672 = ~a7670 & ~a7608;
assign a7674 = ~l600 & ~l564;
assign a7676 = ~l614 & l564;
assign a7678 = ~a7676 & ~a7674;
assign a7680 = ~a7678 & ~l562;
assign a7682 = a7628 & ~l628;
assign a7684 = ~a7682 & ~a7680;
assign a7686 = ~a7684 & a7608;
assign a7688 = ~a7686 & ~a7672;
assign a7690 = a7688 & ~l760;
assign a7692 = ~a7688 & l760;
assign a7694 = ~a7692 & ~a7690;
assign a7696 = l806 & ~l564;
assign a7698 = l820 & l564;
assign a7700 = ~a7698 & ~a7696;
assign a7702 = ~a7700 & ~l562;
assign a7704 = a7628 & l834;
assign a7706 = ~a7704 & ~a7702;
assign a7708 = ~a7706 & a7618;
assign a7710 = a7708 & ~a7616;
assign a7712 = l738 & ~l564;
assign a7714 = l752 & l564;
assign a7716 = ~a7714 & ~a7712;
assign a7718 = ~a7716 & ~l562;
assign a7720 = a7628 & l766;
assign a7722 = ~a7720 & ~a7718;
assign a7724 = ~a7722 & a7616;
assign a7726 = ~a7724 & ~a7710;
assign a7728 = ~a7726 & ~a7612;
assign a7730 = l670 & ~l564;
assign a7732 = l684 & l564;
assign a7734 = ~a7732 & ~a7730;
assign a7736 = ~a7734 & ~l562;
assign a7738 = a7628 & l698;
assign a7740 = ~a7738 & ~a7736;
assign a7742 = ~a7740 & a7612;
assign a7744 = ~a7742 & ~a7728;
assign a7746 = ~a7744 & ~a7608;
assign a7748 = l602 & ~l564;
assign a7750 = l616 & l564;
assign a7752 = ~a7750 & ~a7748;
assign a7754 = ~a7752 & ~l562;
assign a7756 = a7628 & l630;
assign a7758 = ~a7756 & ~a7754;
assign a7760 = ~a7758 & a7608;
assign a7762 = ~a7760 & ~a7746;
assign a7764 = a7762 & ~l762;
assign a7766 = ~a7762 & l762;
assign a7768 = ~a7766 & ~a7764;
assign a7770 = a7768 & a7694;
assign a7772 = ~a7770 & ~a7604;
assign a7774 = a6022 & ~l566;
assign a7776 = l570 & ~l568;
assign a7778 = a7776 & ~l566;
assign a7780 = ~l570 & l568;
assign a7782 = a7780 & ~l566;
assign a7784 = l570 & l568;
assign a7786 = a7784 & ~l566;
assign a7788 = a6022 & l566;
assign a7790 = ~l804 & ~l574;
assign a7792 = ~l818 & l574;
assign a7794 = ~a7792 & ~a7790;
assign a7796 = ~a7794 & ~l572;
assign a7798 = ~l574 & l572;
assign a7800 = a7798 & ~l832;
assign a7802 = ~a7800 & ~a7796;
assign a7804 = ~a7802 & a7788;
assign a7806 = a7804 & ~a7786;
assign a7808 = ~l736 & ~l574;
assign a7810 = ~l750 & l574;
assign a7812 = ~a7810 & ~a7808;
assign a7814 = ~a7812 & ~l572;
assign a7816 = a7798 & ~l764;
assign a7818 = ~a7816 & ~a7814;
assign a7820 = ~a7818 & a7786;
assign a7822 = ~a7820 & ~a7806;
assign a7824 = ~a7822 & ~a7782;
assign a7826 = ~l668 & ~l574;
assign a7828 = ~l682 & l574;
assign a7830 = ~a7828 & ~a7826;
assign a7832 = ~a7830 & ~l572;
assign a7834 = a7798 & ~l696;
assign a7836 = ~a7834 & ~a7832;
assign a7838 = ~a7836 & a7782;
assign a7840 = ~a7838 & ~a7824;
assign a7842 = ~a7840 & ~a7778;
assign a7844 = ~l600 & ~l574;
assign a7846 = ~l614 & l574;
assign a7848 = ~a7846 & ~a7844;
assign a7850 = ~a7848 & ~l572;
assign a7852 = a7798 & ~l628;
assign a7854 = ~a7852 & ~a7850;
assign a7856 = ~a7854 & a7778;
assign a7858 = ~a7856 & ~a7842;
assign a7860 = a7858 & ~l800;
assign a7862 = ~a7858 & l800;
assign a7864 = ~a7862 & ~a7860;
assign a7866 = l806 & ~l574;
assign a7868 = l820 & l574;
assign a7870 = ~a7868 & ~a7866;
assign a7872 = ~a7870 & ~l572;
assign a7874 = a7798 & l834;
assign a7876 = ~a7874 & ~a7872;
assign a7878 = ~a7876 & a7788;
assign a7880 = a7878 & ~a7786;
assign a7882 = l738 & ~l574;
assign a7884 = l752 & l574;
assign a7886 = ~a7884 & ~a7882;
assign a7888 = ~a7886 & ~l572;
assign a7890 = a7798 & l766;
assign a7892 = ~a7890 & ~a7888;
assign a7894 = ~a7892 & a7786;
assign a7896 = ~a7894 & ~a7880;
assign a7898 = ~a7896 & ~a7782;
assign a7900 = l670 & ~l574;
assign a7902 = l684 & l574;
assign a7904 = ~a7902 & ~a7900;
assign a7906 = ~a7904 & ~l572;
assign a7908 = a7798 & l698;
assign a7910 = ~a7908 & ~a7906;
assign a7912 = ~a7910 & a7782;
assign a7914 = ~a7912 & ~a7898;
assign a7916 = ~a7914 & ~a7778;
assign a7918 = l602 & ~l574;
assign a7920 = l616 & l574;
assign a7922 = ~a7920 & ~a7918;
assign a7924 = ~a7922 & ~l572;
assign a7926 = a7798 & l630;
assign a7928 = ~a7926 & ~a7924;
assign a7930 = ~a7928 & a7778;
assign a7932 = ~a7930 & ~a7916;
assign a7934 = a7932 & ~l802;
assign a7936 = ~a7932 & l802;
assign a7938 = ~a7936 & ~a7934;
assign a7940 = a7938 & a7864;
assign a7942 = ~a7940 & ~a7774;
assign a7944 = a6028 & ~l576;
assign a7946 = l580 & ~l578;
assign a7948 = a7946 & ~l576;
assign a7950 = ~l580 & l578;
assign a7952 = a7950 & ~l576;
assign a7954 = l580 & l578;
assign a7956 = a7954 & ~l576;
assign a7958 = a6028 & l576;
assign a7960 = ~l804 & ~l584;
assign a7962 = ~l818 & l584;
assign a7964 = ~a7962 & ~a7960;
assign a7966 = ~a7964 & ~l582;
assign a7968 = ~l584 & l582;
assign a7970 = a7968 & ~l832;
assign a7972 = ~a7970 & ~a7966;
assign a7974 = ~a7972 & a7958;
assign a7976 = a7974 & ~a7956;
assign a7978 = ~l736 & ~l584;
assign a7980 = ~l750 & l584;
assign a7982 = ~a7980 & ~a7978;
assign a7984 = ~a7982 & ~l582;
assign a7986 = a7968 & ~l764;
assign a7988 = ~a7986 & ~a7984;
assign a7990 = ~a7988 & a7956;
assign a7992 = ~a7990 & ~a7976;
assign a7994 = ~a7992 & ~a7952;
assign a7996 = ~l668 & ~l584;
assign a7998 = ~l682 & l584;
assign a8000 = ~a7998 & ~a7996;
assign a8002 = ~a8000 & ~l582;
assign a8004 = a7968 & ~l696;
assign a8006 = ~a8004 & ~a8002;
assign a8008 = ~a8006 & a7952;
assign a8010 = ~a8008 & ~a7994;
assign a8012 = ~a8010 & ~a7948;
assign a8014 = ~l600 & ~l584;
assign a8016 = ~l614 & l584;
assign a8018 = ~a8016 & ~a8014;
assign a8020 = ~a8018 & ~l582;
assign a8022 = a7968 & ~l628;
assign a8024 = ~a8022 & ~a8020;
assign a8026 = ~a8024 & a7948;
assign a8028 = ~a8026 & ~a8012;
assign a8030 = a8028 & ~l814;
assign a8032 = ~a8028 & l814;
assign a8034 = ~a8032 & ~a8030;
assign a8036 = l806 & ~l584;
assign a8038 = l820 & l584;
assign a8040 = ~a8038 & ~a8036;
assign a8042 = ~a8040 & ~l582;
assign a8044 = a7968 & l834;
assign a8046 = ~a8044 & ~a8042;
assign a8048 = ~a8046 & a7958;
assign a8050 = a8048 & ~a7956;
assign a8052 = l738 & ~l584;
assign a8054 = l752 & l584;
assign a8056 = ~a8054 & ~a8052;
assign a8058 = ~a8056 & ~l582;
assign a8060 = a7968 & l766;
assign a8062 = ~a8060 & ~a8058;
assign a8064 = ~a8062 & a7956;
assign a8066 = ~a8064 & ~a8050;
assign a8068 = ~a8066 & ~a7952;
assign a8070 = l670 & ~l584;
assign a8072 = l684 & l584;
assign a8074 = ~a8072 & ~a8070;
assign a8076 = ~a8074 & ~l582;
assign a8078 = a7968 & l698;
assign a8080 = ~a8078 & ~a8076;
assign a8082 = ~a8080 & a7952;
assign a8084 = ~a8082 & ~a8068;
assign a8086 = ~a8084 & ~a7948;
assign a8088 = l602 & ~l584;
assign a8090 = l616 & l584;
assign a8092 = ~a8090 & ~a8088;
assign a8094 = ~a8092 & ~l582;
assign a8096 = a7968 & l630;
assign a8098 = ~a8096 & ~a8094;
assign a8100 = ~a8098 & a7948;
assign a8102 = ~a8100 & ~a8086;
assign a8104 = a8102 & ~l816;
assign a8106 = ~a8102 & l816;
assign a8108 = ~a8106 & ~a8104;
assign a8110 = a8108 & a8034;
assign a8112 = ~a8110 & ~a7944;
assign a8114 = a6034 & ~l586;
assign a8116 = l590 & ~l588;
assign a8118 = a8116 & ~l586;
assign a8120 = ~l590 & l588;
assign a8122 = a8120 & ~l586;
assign a8124 = l590 & l588;
assign a8126 = a8124 & ~l586;
assign a8128 = a6034 & l586;
assign a8130 = ~l804 & ~l594;
assign a8132 = ~l818 & l594;
assign a8134 = ~a8132 & ~a8130;
assign a8136 = ~a8134 & ~l592;
assign a8138 = ~l594 & l592;
assign a8140 = a8138 & ~l832;
assign a8142 = ~a8140 & ~a8136;
assign a8144 = ~a8142 & a8128;
assign a8146 = a8144 & ~a8126;
assign a8148 = ~l736 & ~l594;
assign a8150 = ~l750 & l594;
assign a8152 = ~a8150 & ~a8148;
assign a8154 = ~a8152 & ~l592;
assign a8156 = a8138 & ~l764;
assign a8158 = ~a8156 & ~a8154;
assign a8160 = ~a8158 & a8126;
assign a8162 = ~a8160 & ~a8146;
assign a8164 = ~a8162 & ~a8122;
assign a8166 = ~l668 & ~l594;
assign a8168 = ~l682 & l594;
assign a8170 = ~a8168 & ~a8166;
assign a8172 = ~a8170 & ~l592;
assign a8174 = a8138 & ~l696;
assign a8176 = ~a8174 & ~a8172;
assign a8178 = ~a8176 & a8122;
assign a8180 = ~a8178 & ~a8164;
assign a8182 = ~a8180 & ~a8118;
assign a8184 = ~l600 & ~l594;
assign a8186 = ~l614 & l594;
assign a8188 = ~a8186 & ~a8184;
assign a8190 = ~a8188 & ~l592;
assign a8192 = a8138 & ~l628;
assign a8194 = ~a8192 & ~a8190;
assign a8196 = ~a8194 & a8118;
assign a8198 = ~a8196 & ~a8182;
assign a8200 = a8198 & ~l828;
assign a8202 = ~a8198 & l828;
assign a8204 = ~a8202 & ~a8200;
assign a8206 = l806 & ~l594;
assign a8208 = l820 & l594;
assign a8210 = ~a8208 & ~a8206;
assign a8212 = ~a8210 & ~l592;
assign a8214 = a8138 & l834;
assign a8216 = ~a8214 & ~a8212;
assign a8218 = ~a8216 & a8128;
assign a8220 = a8218 & ~a8126;
assign a8222 = l738 & ~l594;
assign a8224 = l752 & l594;
assign a8226 = ~a8224 & ~a8222;
assign a8228 = ~a8226 & ~l592;
assign a8230 = a8138 & l766;
assign a8232 = ~a8230 & ~a8228;
assign a8234 = ~a8232 & a8126;
assign a8236 = ~a8234 & ~a8220;
assign a8238 = ~a8236 & ~a8122;
assign a8240 = l670 & ~l594;
assign a8242 = l684 & l594;
assign a8244 = ~a8242 & ~a8240;
assign a8246 = ~a8244 & ~l592;
assign a8248 = a8138 & l698;
assign a8250 = ~a8248 & ~a8246;
assign a8252 = ~a8250 & a8122;
assign a8254 = ~a8252 & ~a8238;
assign a8256 = ~a8254 & ~a8118;
assign a8258 = l602 & ~l594;
assign a8260 = l616 & l594;
assign a8262 = ~a8260 & ~a8258;
assign a8264 = ~a8262 & ~l592;
assign a8266 = a8138 & l630;
assign a8268 = ~a8266 & ~a8264;
assign a8270 = ~a8268 & a8118;
assign a8272 = ~a8270 & ~a8256;
assign a8274 = a8272 & ~l830;
assign a8276 = ~a8272 & l830;
assign a8278 = ~a8276 & ~a8274;
assign a8280 = a8278 & a8204;
assign a8282 = ~a8280 & ~a8114;
assign a8284 = ~l574 & ~l572;
assign a8286 = a8284 & a7778;
assign a8288 = ~a8286 & ~l484;
assign a8290 = ~l584 & ~l582;
assign a8292 = a8290 & a7948;
assign a8294 = ~a8292 & l484;
assign a8296 = ~a8294 & ~a8288;
assign a8298 = ~a8296 & ~l482;
assign a8300 = ~l594 & ~l592;
assign a8302 = a8300 & a8118;
assign a8304 = ~a8302 & a6268;
assign a8306 = ~a8304 & ~a8298;
assign a8308 = ~a8306 & a6258;
assign a8310 = a8308 & ~a6256;
assign a8312 = ~l544 & ~l542;
assign a8314 = a8312 & a7268;
assign a8316 = ~a8314 & ~l484;
assign a8318 = ~l554 & ~l552;
assign a8320 = a8318 & a7438;
assign a8322 = ~a8320 & l484;
assign a8324 = ~a8322 & ~a8316;
assign a8326 = ~a8324 & ~l482;
assign a8328 = ~l564 & ~l562;
assign a8330 = a8328 & a7608;
assign a8332 = ~a8330 & a6268;
assign a8334 = ~a8332 & ~a8326;
assign a8336 = ~a8334 & a6256;
assign a8338 = ~a8336 & ~a8310;
assign a8340 = ~a8338 & ~a6252;
assign a8342 = ~l514 & ~l512;
assign a8344 = a8342 & a6758;
assign a8346 = ~a8344 & ~l484;
assign a8348 = ~l524 & ~l522;
assign a8350 = a8348 & a6928;
assign a8352 = ~a8350 & l484;
assign a8354 = ~a8352 & ~a8346;
assign a8356 = ~a8354 & ~l482;
assign a8358 = ~l534 & ~l532;
assign a8360 = a8358 & a7098;
assign a8362 = ~a8360 & a6268;
assign a8364 = ~a8362 & ~a8356;
assign a8366 = ~a8364 & a6252;
assign a8368 = ~a8366 & ~a8340;
assign a8370 = ~a8368 & ~a6248;
assign a8372 = ~l484 & ~l482;
assign a8374 = a8372 & a6248;
assign a8376 = ~a8374 & ~l484;
assign a8378 = ~l494 & ~l492;
assign a8380 = a8378 & a6418;
assign a8382 = ~a8380 & l484;
assign a8384 = ~a8382 & ~a8376;
assign a8386 = ~a8384 & ~l482;
assign a8388 = ~l504 & ~l502;
assign a8390 = a8388 & a6588;
assign a8392 = ~a8390 & a6268;
assign a8394 = ~a8392 & ~a8386;
assign a8396 = ~a8394 & a6248;
assign a8398 = ~a8396 & ~a8370;
assign a8400 = l574 & ~l572;
assign a8402 = a8400 & a7778;
assign a8404 = ~a8402 & ~l494;
assign a8406 = l584 & ~l582;
assign a8408 = a8406 & a7948;
assign a8410 = ~a8408 & l494;
assign a8412 = ~a8410 & ~a8404;
assign a8414 = ~a8412 & ~l492;
assign a8416 = l594 & ~l592;
assign a8418 = a8416 & a8118;
assign a8420 = ~a8418 & a6438;
assign a8422 = ~a8420 & ~a8414;
assign a8424 = ~a8422 & a6428;
assign a8426 = a8424 & ~a6426;
assign a8428 = l544 & ~l542;
assign a8430 = a8428 & a7268;
assign a8432 = ~a8430 & ~l494;
assign a8434 = l554 & ~l552;
assign a8436 = a8434 & a7438;
assign a8438 = ~a8436 & l494;
assign a8440 = ~a8438 & ~a8432;
assign a8442 = ~a8440 & ~l492;
assign a8444 = l564 & ~l562;
assign a8446 = a8444 & a7608;
assign a8448 = ~a8446 & a6438;
assign a8450 = ~a8448 & ~a8442;
assign a8452 = ~a8450 & a6426;
assign a8454 = ~a8452 & ~a8426;
assign a8456 = ~a8454 & ~a6422;
assign a8458 = l514 & ~l512;
assign a8460 = a8458 & a6758;
assign a8462 = ~a8460 & ~l494;
assign a8464 = l524 & ~l522;
assign a8466 = a8464 & a6928;
assign a8468 = ~a8466 & l494;
assign a8470 = ~a8468 & ~a8462;
assign a8472 = ~a8470 & ~l492;
assign a8474 = l534 & ~l532;
assign a8476 = a8474 & a7098;
assign a8478 = ~a8476 & a6438;
assign a8480 = ~a8478 & ~a8472;
assign a8482 = ~a8480 & a6422;
assign a8484 = ~a8482 & ~a8456;
assign a8486 = ~a8484 & ~a6418;
assign a8488 = l484 & ~l482;
assign a8490 = a8488 & a6248;
assign a8492 = ~a8490 & ~l494;
assign a8494 = l494 & ~l492;
assign a8496 = a8494 & a6418;
assign a8498 = ~a8496 & l494;
assign a8500 = ~a8498 & ~a8492;
assign a8502 = ~a8500 & ~l492;
assign a8504 = l504 & ~l502;
assign a8506 = a8504 & a6588;
assign a8508 = ~a8506 & a6438;
assign a8510 = ~a8508 & ~a8502;
assign a8512 = ~a8510 & a6418;
assign a8514 = ~a8512 & ~a8486;
assign a8516 = a7798 & a7778;
assign a8518 = ~a8516 & ~l504;
assign a8520 = a7968 & a7948;
assign a8522 = ~a8520 & l504;
assign a8524 = ~a8522 & ~a8518;
assign a8526 = ~a8524 & ~l502;
assign a8528 = a8138 & a8118;
assign a8530 = ~a8528 & a6608;
assign a8532 = ~a8530 & ~a8526;
assign a8534 = ~a8532 & a6598;
assign a8536 = a8534 & ~a6596;
assign a8538 = a7288 & a7268;
assign a8540 = ~a8538 & ~l504;
assign a8542 = a7458 & a7438;
assign a8544 = ~a8542 & l504;
assign a8546 = ~a8544 & ~a8540;
assign a8548 = ~a8546 & ~l502;
assign a8550 = a7628 & a7608;
assign a8552 = ~a8550 & a6608;
assign a8554 = ~a8552 & ~a8548;
assign a8556 = ~a8554 & a6596;
assign a8558 = ~a8556 & ~a8536;
assign a8560 = ~a8558 & ~a6592;
assign a8562 = a6778 & a6758;
assign a8564 = ~a8562 & ~l504;
assign a8566 = a6948 & a6928;
assign a8568 = ~a8566 & l504;
assign a8570 = ~a8568 & ~a8564;
assign a8572 = ~a8570 & ~l502;
assign a8574 = a7118 & a7098;
assign a8576 = ~a8574 & a6608;
assign a8578 = ~a8576 & ~a8572;
assign a8580 = ~a8578 & a6592;
assign a8582 = ~a8580 & ~a8560;
assign a8584 = ~a8582 & ~a6588;
assign a8586 = a6268 & a6248;
assign a8588 = ~a8586 & ~l504;
assign a8590 = a6438 & a6418;
assign a8592 = ~a8590 & l504;
assign a8594 = ~a8592 & ~a8588;
assign a8596 = ~a8594 & ~l502;
assign a8598 = a6608 & ~a6588;
assign a8600 = ~a8598 & ~a8596;
assign a8602 = ~a8600 & a6588;
assign a8604 = ~a8602 & ~a8584;
assign a8606 = a8284 & a7782;
assign a8608 = ~a8606 & ~l514;
assign a8610 = a8290 & a7952;
assign a8612 = ~a8610 & l514;
assign a8614 = ~a8612 & ~a8608;
assign a8616 = ~a8614 & ~l512;
assign a8618 = a8300 & a8122;
assign a8620 = ~a8618 & a6778;
assign a8622 = ~a8620 & ~a8616;
assign a8624 = ~a8622 & a6768;
assign a8626 = a8624 & ~a6766;
assign a8628 = a8312 & a7272;
assign a8630 = ~a8628 & ~l514;
assign a8632 = a8318 & a7442;
assign a8634 = ~a8632 & l514;
assign a8636 = ~a8634 & ~a8630;
assign a8638 = ~a8636 & ~l512;
assign a8640 = a8328 & a7612;
assign a8642 = ~a8640 & a6778;
assign a8644 = ~a8642 & ~a8638;
assign a8646 = ~a8644 & a6766;
assign a8648 = ~a8646 & ~a8626;
assign a8650 = ~a8648 & ~a6762;
assign a8652 = a8342 & a6762;
assign a8654 = ~a8652 & ~l514;
assign a8656 = a8348 & a6932;
assign a8658 = ~a8656 & l514;
assign a8660 = ~a8658 & ~a8654;
assign a8662 = ~a8660 & ~l512;
assign a8664 = a8358 & a7102;
assign a8666 = ~a8664 & a6778;
assign a8668 = ~a8666 & ~a8662;
assign a8670 = ~a8668 & a6762;
assign a8672 = ~a8670 & ~a8650;
assign a8674 = ~a8672 & ~a6758;
assign a8676 = a8372 & a6252;
assign a8678 = ~a8676 & ~l514;
assign a8680 = a8378 & a6422;
assign a8682 = ~a8680 & l514;
assign a8684 = ~a8682 & ~a8678;
assign a8686 = ~a8684 & ~l512;
assign a8688 = a8388 & a6592;
assign a8690 = ~a8688 & a6778;
assign a8692 = ~a8690 & ~a8686;
assign a8694 = ~a8692 & a6758;
assign a8696 = ~a8694 & ~a8674;
assign a8698 = a8400 & a7782;
assign a8700 = ~a8698 & ~l524;
assign a8702 = a8406 & a7952;
assign a8704 = ~a8702 & l524;
assign a8706 = ~a8704 & ~a8700;
assign a8708 = ~a8706 & ~l522;
assign a8710 = a8416 & a8122;
assign a8712 = ~a8710 & a6948;
assign a8714 = ~a8712 & ~a8708;
assign a8716 = ~a8714 & a6938;
assign a8718 = a8716 & ~a6936;
assign a8720 = a8428 & a7272;
assign a8722 = ~a8720 & ~l524;
assign a8724 = a8434 & a7442;
assign a8726 = ~a8724 & l524;
assign a8728 = ~a8726 & ~a8722;
assign a8730 = ~a8728 & ~l522;
assign a8732 = a8444 & a7612;
assign a8734 = ~a8732 & a6948;
assign a8736 = ~a8734 & ~a8730;
assign a8738 = ~a8736 & a6936;
assign a8740 = ~a8738 & ~a8718;
assign a8742 = ~a8740 & ~a6932;
assign a8744 = a8458 & a6762;
assign a8746 = ~a8744 & ~l524;
assign a8748 = a8464 & a6932;
assign a8750 = ~a8748 & l524;
assign a8752 = ~a8750 & ~a8746;
assign a8754 = ~a8752 & ~l522;
assign a8756 = a8474 & a7102;
assign a8758 = ~a8756 & a6948;
assign a8760 = ~a8758 & ~a8754;
assign a8762 = ~a8760 & a6932;
assign a8764 = ~a8762 & ~a8742;
assign a8766 = ~a8764 & ~a6928;
assign a8768 = a8488 & a6252;
assign a8770 = ~a8768 & ~l524;
assign a8772 = a8494 & a6422;
assign a8774 = ~a8772 & l524;
assign a8776 = ~a8774 & ~a8770;
assign a8778 = ~a8776 & ~l522;
assign a8780 = a8504 & a6592;
assign a8782 = ~a8780 & a6948;
assign a8784 = ~a8782 & ~a8778;
assign a8786 = ~a8784 & a6928;
assign a8788 = ~a8786 & ~a8766;
assign a8790 = a7798 & a7782;
assign a8792 = ~a8790 & ~l534;
assign a8794 = a7968 & a7952;
assign a8796 = ~a8794 & l534;
assign a8798 = ~a8796 & ~a8792;
assign a8800 = ~a8798 & ~l532;
assign a8802 = a8138 & a8122;
assign a8804 = ~a8802 & a7118;
assign a8806 = ~a8804 & ~a8800;
assign a8808 = ~a8806 & a7108;
assign a8810 = a8808 & ~a7106;
assign a8812 = a7288 & a7272;
assign a8814 = ~a8812 & ~l534;
assign a8816 = a7458 & a7442;
assign a8818 = ~a8816 & l534;
assign a8820 = ~a8818 & ~a8814;
assign a8822 = ~a8820 & ~l532;
assign a8824 = a7628 & a7612;
assign a8826 = ~a8824 & a7118;
assign a8828 = ~a8826 & ~a8822;
assign a8830 = ~a8828 & a7106;
assign a8832 = ~a8830 & ~a8810;
assign a8834 = ~a8832 & ~a7102;
assign a8836 = a6778 & a6762;
assign a8838 = ~a8836 & ~l534;
assign a8840 = a6948 & a6932;
assign a8842 = ~a8840 & l534;
assign a8844 = ~a8842 & ~a8838;
assign a8846 = ~a8844 & ~l532;
assign a8848 = a7118 & ~a7102;
assign a8850 = ~a8848 & ~a8846;
assign a8852 = ~a8850 & a7102;
assign a8854 = ~a8852 & ~a8834;
assign a8856 = ~a8854 & ~a7098;
assign a8858 = a6268 & a6252;
assign a8860 = ~a8858 & ~l534;
assign a8862 = a6438 & a6422;
assign a8864 = ~a8862 & l534;
assign a8866 = ~a8864 & ~a8860;
assign a8868 = ~a8866 & ~l532;
assign a8870 = a6608 & a6592;
assign a8872 = ~a8870 & a7118;
assign a8874 = ~a8872 & ~a8868;
assign a8876 = ~a8874 & a7098;
assign a8878 = ~a8876 & ~a8856;
assign a8880 = a8284 & a7786;
assign a8882 = ~a8880 & ~l544;
assign a8884 = a8290 & a7956;
assign a8886 = ~a8884 & l544;
assign a8888 = ~a8886 & ~a8882;
assign a8890 = ~a8888 & ~l542;
assign a8892 = a8300 & a8126;
assign a8894 = ~a8892 & a7288;
assign a8896 = ~a8894 & ~a8890;
assign a8898 = ~a8896 & a7278;
assign a8900 = a8898 & ~a7276;
assign a8902 = a8312 & a7276;
assign a8904 = ~a8902 & ~l544;
assign a8906 = a8318 & a7446;
assign a8908 = ~a8906 & l544;
assign a8910 = ~a8908 & ~a8904;
assign a8912 = ~a8910 & ~l542;
assign a8914 = a8328 & a7616;
assign a8916 = ~a8914 & a7288;
assign a8918 = ~a8916 & ~a8912;
assign a8920 = ~a8918 & a7276;
assign a8922 = ~a8920 & ~a8900;
assign a8924 = ~a8922 & ~a7272;
assign a8926 = a8342 & a6766;
assign a8928 = ~a8926 & ~l544;
assign a8930 = a8348 & a6936;
assign a8932 = ~a8930 & l544;
assign a8934 = ~a8932 & ~a8928;
assign a8936 = ~a8934 & ~l542;
assign a8938 = a8358 & a7106;
assign a8940 = ~a8938 & a7288;
assign a8942 = ~a8940 & ~a8936;
assign a8944 = ~a8942 & a7272;
assign a8946 = ~a8944 & ~a8924;
assign a8948 = ~a8946 & ~a7268;
assign a8950 = a8372 & a6256;
assign a8952 = ~a8950 & ~l544;
assign a8954 = a8378 & a6426;
assign a8956 = ~a8954 & l544;
assign a8958 = ~a8956 & ~a8952;
assign a8960 = ~a8958 & ~l542;
assign a8962 = a8388 & a6596;
assign a8964 = ~a8962 & a7288;
assign a8966 = ~a8964 & ~a8960;
assign a8968 = ~a8966 & a7268;
assign a8970 = ~a8968 & ~a8948;
assign a8972 = a8400 & a7786;
assign a8974 = ~a8972 & ~l554;
assign a8976 = a8406 & a7956;
assign a8978 = ~a8976 & l554;
assign a8980 = ~a8978 & ~a8974;
assign a8982 = ~a8980 & ~l552;
assign a8984 = a8416 & a8126;
assign a8986 = ~a8984 & a7458;
assign a8988 = ~a8986 & ~a8982;
assign a8990 = ~a8988 & a7448;
assign a8992 = a8990 & ~a7446;
assign a8994 = a8428 & a7276;
assign a8996 = ~a8994 & ~l554;
assign a8998 = a8434 & a7446;
assign a9000 = ~a8998 & l554;
assign a9002 = ~a9000 & ~a8996;
assign a9004 = ~a9002 & ~l552;
assign a9006 = a8444 & a7616;
assign a9008 = ~a9006 & a7458;
assign a9010 = ~a9008 & ~a9004;
assign a9012 = ~a9010 & a7446;
assign a9014 = ~a9012 & ~a8992;
assign a9016 = ~a9014 & ~a7442;
assign a9018 = a8458 & a6766;
assign a9020 = ~a9018 & ~l554;
assign a9022 = a8464 & a6936;
assign a9024 = ~a9022 & l554;
assign a9026 = ~a9024 & ~a9020;
assign a9028 = ~a9026 & ~l552;
assign a9030 = a8474 & a7106;
assign a9032 = ~a9030 & a7458;
assign a9034 = ~a9032 & ~a9028;
assign a9036 = ~a9034 & a7442;
assign a9038 = ~a9036 & ~a9016;
assign a9040 = ~a9038 & ~a7438;
assign a9042 = a8488 & a6256;
assign a9044 = ~a9042 & ~l554;
assign a9046 = a8494 & a6426;
assign a9048 = ~a9046 & l554;
assign a9050 = ~a9048 & ~a9044;
assign a9052 = ~a9050 & ~l552;
assign a9054 = a8504 & a6596;
assign a9056 = ~a9054 & a7458;
assign a9058 = ~a9056 & ~a9052;
assign a9060 = ~a9058 & a7438;
assign a9062 = ~a9060 & ~a9040;
assign a9064 = a7798 & a7786;
assign a9066 = ~a9064 & ~l564;
assign a9068 = a7968 & a7956;
assign a9070 = ~a9068 & l564;
assign a9072 = ~a9070 & ~a9066;
assign a9074 = ~a9072 & ~l562;
assign a9076 = a8138 & a8126;
assign a9078 = ~a9076 & a7628;
assign a9080 = ~a9078 & ~a9074;
assign a9082 = ~a9080 & a7618;
assign a9084 = a9082 & ~a7616;
assign a9086 = a7288 & a7276;
assign a9088 = ~a9086 & ~l564;
assign a9090 = a7458 & a7446;
assign a9092 = ~a9090 & l564;
assign a9094 = ~a9092 & ~a9088;
assign a9096 = ~a9094 & ~l562;
assign a9098 = a7628 & ~a7616;
assign a9100 = ~a9098 & ~a9096;
assign a9102 = ~a9100 & a7616;
assign a9104 = ~a9102 & ~a9084;
assign a9106 = ~a9104 & ~a7612;
assign a9108 = a6778 & a6766;
assign a9110 = ~a9108 & ~l564;
assign a9112 = a6948 & a6936;
assign a9114 = ~a9112 & l564;
assign a9116 = ~a9114 & ~a9110;
assign a9118 = ~a9116 & ~l562;
assign a9120 = a7118 & a7106;
assign a9122 = ~a9120 & a7628;
assign a9124 = ~a9122 & ~a9118;
assign a9126 = ~a9124 & a7612;
assign a9128 = ~a9126 & ~a9106;
assign a9130 = ~a9128 & ~a7608;
assign a9132 = a6268 & a6256;
assign a9134 = ~a9132 & ~l564;
assign a9136 = a6438 & a6426;
assign a9138 = ~a9136 & l564;
assign a9140 = ~a9138 & ~a9134;
assign a9142 = ~a9140 & ~l562;
assign a9144 = a6608 & a6596;
assign a9146 = ~a9144 & a7628;
assign a9148 = ~a9146 & ~a9142;
assign a9150 = ~a9148 & a7608;
assign a9152 = ~a9150 & ~a9130;
assign a9154 = a8284 & a7788;
assign a9156 = ~a9154 & ~l574;
assign a9158 = a8290 & a7958;
assign a9160 = ~a9158 & l574;
assign a9162 = ~a9160 & ~a9156;
assign a9164 = ~a9162 & ~l572;
assign a9166 = a8300 & a8128;
assign a9168 = ~a9166 & a7798;
assign a9170 = ~a9168 & ~a9164;
assign a9172 = ~a9170 & a7788;
assign a9174 = a9172 & ~a7786;
assign a9176 = a8312 & a7278;
assign a9178 = ~a9176 & ~l574;
assign a9180 = a8318 & a7448;
assign a9182 = ~a9180 & l574;
assign a9184 = ~a9182 & ~a9178;
assign a9186 = ~a9184 & ~l572;
assign a9188 = a8328 & a7618;
assign a9190 = ~a9188 & a7798;
assign a9192 = ~a9190 & ~a9186;
assign a9194 = ~a9192 & a7786;
assign a9196 = ~a9194 & ~a9174;
assign a9198 = ~a9196 & ~a7782;
assign a9200 = a8342 & a6768;
assign a9202 = ~a9200 & ~l574;
assign a9204 = a8348 & a6938;
assign a9206 = ~a9204 & l574;
assign a9208 = ~a9206 & ~a9202;
assign a9210 = ~a9208 & ~l572;
assign a9212 = a8358 & a7108;
assign a9214 = ~a9212 & a7798;
assign a9216 = ~a9214 & ~a9210;
assign a9218 = ~a9216 & a7782;
assign a9220 = ~a9218 & ~a9198;
assign a9222 = ~a9220 & ~a7778;
assign a9224 = a8372 & a6258;
assign a9226 = ~a9224 & ~l574;
assign a9228 = a8378 & a6428;
assign a9230 = ~a9228 & l574;
assign a9232 = ~a9230 & ~a9226;
assign a9234 = ~a9232 & ~l572;
assign a9236 = a8388 & a6598;
assign a9238 = ~a9236 & a7798;
assign a9240 = ~a9238 & ~a9234;
assign a9242 = ~a9240 & a7778;
assign a9244 = ~a9242 & ~a9222;
assign a9246 = a8400 & a7788;
assign a9248 = ~a9246 & ~l584;
assign a9250 = a8406 & a7958;
assign a9252 = ~a9250 & l584;
assign a9254 = ~a9252 & ~a9248;
assign a9256 = ~a9254 & ~l582;
assign a9258 = a8416 & a8128;
assign a9260 = ~a9258 & a7968;
assign a9262 = ~a9260 & ~a9256;
assign a9264 = ~a9262 & a7958;
assign a9266 = a9264 & ~a7956;
assign a9268 = a8428 & a7278;
assign a9270 = ~a9268 & ~l584;
assign a9272 = a8434 & a7448;
assign a9274 = ~a9272 & l584;
assign a9276 = ~a9274 & ~a9270;
assign a9278 = ~a9276 & ~l582;
assign a9280 = a8444 & a7618;
assign a9282 = ~a9280 & a7968;
assign a9284 = ~a9282 & ~a9278;
assign a9286 = ~a9284 & a7956;
assign a9288 = ~a9286 & ~a9266;
assign a9290 = ~a9288 & ~a7952;
assign a9292 = a8458 & a6768;
assign a9294 = ~a9292 & ~l584;
assign a9296 = a8464 & a6938;
assign a9298 = ~a9296 & l584;
assign a9300 = ~a9298 & ~a9294;
assign a9302 = ~a9300 & ~l582;
assign a9304 = a8474 & a7108;
assign a9306 = ~a9304 & a7968;
assign a9308 = ~a9306 & ~a9302;
assign a9310 = ~a9308 & a7952;
assign a9312 = ~a9310 & ~a9290;
assign a9314 = ~a9312 & ~a7948;
assign a9316 = a8488 & a6258;
assign a9318 = ~a9316 & ~l584;
assign a9320 = a8494 & a6428;
assign a9322 = ~a9320 & l584;
assign a9324 = ~a9322 & ~a9318;
assign a9326 = ~a9324 & ~l582;
assign a9328 = a8504 & a6598;
assign a9330 = ~a9328 & a7968;
assign a9332 = ~a9330 & ~a9326;
assign a9334 = ~a9332 & a7948;
assign a9336 = ~a9334 & ~a9314;
assign a9338 = a7798 & a7788;
assign a9340 = ~a9338 & ~l594;
assign a9342 = a7968 & a7958;
assign a9344 = ~a9342 & l594;
assign a9346 = ~a9344 & ~a9340;
assign a9348 = ~a9346 & ~l592;
assign a9350 = a8138 & ~a8128;
assign a9352 = ~a9350 & ~a9348;
assign a9354 = ~a9352 & a8128;
assign a9356 = a9354 & ~a8126;
assign a9358 = a7288 & a7278;
assign a9360 = ~a9358 & ~l594;
assign a9362 = a7458 & a7448;
assign a9364 = ~a9362 & l594;
assign a9366 = ~a9364 & ~a9360;
assign a9368 = ~a9366 & ~l592;
assign a9370 = a7628 & a7618;
assign a9372 = ~a9370 & a8138;
assign a9374 = ~a9372 & ~a9368;
assign a9376 = ~a9374 & a8126;
assign a9378 = ~a9376 & ~a9356;
assign a9380 = ~a9378 & ~a8122;
assign a9382 = a6778 & a6768;
assign a9384 = ~a9382 & ~l594;
assign a9386 = a6948 & a6938;
assign a9388 = ~a9386 & l594;
assign a9390 = ~a9388 & ~a9384;
assign a9392 = ~a9390 & ~l592;
assign a9394 = a7118 & a7108;
assign a9396 = ~a9394 & a8138;
assign a9398 = ~a9396 & ~a9392;
assign a9400 = ~a9398 & a8122;
assign a9402 = ~a9400 & ~a9380;
assign a9404 = ~a9402 & ~a8118;
assign a9406 = a6268 & a6258;
assign a9408 = ~a9406 & ~l594;
assign a9410 = a6438 & a6428;
assign a9412 = ~a9410 & l594;
assign a9414 = ~a9412 & ~a9408;
assign a9416 = ~a9414 & ~l592;
assign a9418 = a6608 & a6598;
assign a9420 = ~a9418 & a8138;
assign a9422 = ~a9420 & ~a9416;
assign a9424 = ~a9422 & a8118;
assign a9426 = ~a9424 & ~a9404;
assign a9428 = ~a8342 & a6758;
assign a9430 = ~a8348 & a6928;
assign a9432 = ~a9430 & ~a9428;
assign a9434 = ~a8358 & a7098;
assign a9436 = ~a9434 & a9432;
assign a9438 = ~a8312 & a7268;
assign a9440 = ~a6936 & ~a6766;
assign a9442 = a9440 & ~a7106;
assign a9444 = ~a6938 & ~a6768;
assign a9446 = a9444 & ~a7108;
assign a9448 = ~a7956 & ~a7786;
assign a9450 = a9448 & ~a8126;
assign a9452 = ~a9450 & ~a9446;
assign a9454 = ~a9452 & a9442;
assign a9456 = ~a9454 & a9438;
assign a9458 = ~a8318 & a7438;
assign a9460 = a9458 & ~a9454;
assign a9462 = ~a8328 & a7608;
assign a9464 = a9462 & ~a9454;
assign a9466 = ~a8284 & a7778;
assign a9468 = ~a7448 & ~a7278;
assign a9470 = a9468 & ~a7618;
assign a9472 = ~a9470 & ~a9442;
assign a9474 = ~a9472 & a9446;
assign a9476 = ~a9474 & a9466;
assign a9478 = ~a8290 & a7948;
assign a9480 = a9478 & ~a9474;
assign a9482 = ~a8300 & a8118;
assign a9484 = a9482 & ~a9474;
assign a9486 = ~a9484 & ~a9480;
assign a9488 = a9486 & ~a9476;
assign a9490 = a9488 & ~a9464;
assign a9492 = a9490 & ~a9460;
assign a9494 = a9492 & ~a9456;
assign a9496 = a9494 & a9436;
assign a9498 = ~a9496 & a6252;
assign a9500 = ~a8458 & a6758;
assign a9502 = ~a8464 & a6928;
assign a9504 = ~a9502 & ~a9500;
assign a9506 = ~a8474 & a7098;
assign a9508 = ~a9506 & a9504;
assign a9510 = ~a8428 & a7268;
assign a9512 = a9510 & ~a9454;
assign a9514 = ~a8434 & a7438;
assign a9516 = a9514 & ~a9454;
assign a9518 = ~a8444 & a7608;
assign a9520 = a9518 & ~a9454;
assign a9522 = ~a8400 & a7778;
assign a9524 = a9522 & ~a9474;
assign a9526 = ~a8406 & a7948;
assign a9528 = a9526 & ~a9474;
assign a9530 = ~a8416 & a8118;
assign a9532 = a9530 & ~a9474;
assign a9534 = ~a9532 & ~a9528;
assign a9536 = a9534 & ~a9524;
assign a9538 = a9536 & ~a9520;
assign a9540 = a9538 & ~a9516;
assign a9542 = a9540 & ~a9512;
assign a9544 = a9542 & a9508;
assign a9546 = ~a9544 & a6422;
assign a9548 = ~a6778 & a6758;
assign a9550 = ~a6948 & a6928;
assign a9552 = ~a9550 & ~a9548;
assign a9554 = ~a7118 & a7098;
assign a9556 = ~a9554 & a9552;
assign a9558 = ~a7288 & a7268;
assign a9560 = a9558 & ~a9454;
assign a9562 = ~a7458 & a7438;
assign a9564 = a9562 & ~a9454;
assign a9566 = ~a7628 & a7608;
assign a9568 = a9566 & ~a9454;
assign a9570 = ~a7798 & a7778;
assign a9572 = a9570 & ~a9474;
assign a9574 = ~a7968 & a7948;
assign a9576 = a9574 & ~a9474;
assign a9578 = ~a8138 & a8118;
assign a9580 = a9578 & ~a9474;
assign a9582 = ~a9580 & ~a9576;
assign a9584 = a9582 & ~a9572;
assign a9586 = a9584 & ~a9568;
assign a9588 = a9586 & ~a9564;
assign a9590 = a9588 & ~a9560;
assign a9592 = a9590 & a9556;
assign a9594 = ~a9592 & a6592;
assign a9596 = ~a7442 & ~a7272;
assign a9598 = a9596 & ~a7612;
assign a9600 = ~a7952 & ~a7782;
assign a9602 = a9600 & ~a8122;
assign a9604 = ~a9602 & ~a9470;
assign a9606 = ~a9604 & a9598;
assign a9608 = ~a9606 & ~a9436;
assign a9610 = ~a9598 & ~a9446;
assign a9612 = ~a9610 & a9470;
assign a9614 = ~a9612 & a9466;
assign a9616 = ~a9612 & a9478;
assign a9618 = ~a9612 & a9482;
assign a9620 = ~a9618 & ~a9616;
assign a9622 = a9620 & ~a9614;
assign a9624 = a9622 & ~a9608;
assign a9626 = a9624 & ~a9438;
assign a9628 = a9626 & ~a9458;
assign a9630 = a9628 & ~a9462;
assign a9632 = ~a9630 & a6256;
assign a9634 = ~a9606 & ~a9508;
assign a9636 = ~a9612 & a9522;
assign a9638 = ~a9612 & a9526;
assign a9640 = ~a9612 & a9530;
assign a9642 = ~a9640 & ~a9638;
assign a9644 = a9642 & ~a9636;
assign a9646 = a9644 & ~a9634;
assign a9648 = a9646 & ~a9510;
assign a9650 = a9648 & ~a9514;
assign a9652 = a9650 & ~a9518;
assign a9654 = ~a9652 & a6426;
assign a9656 = ~a9606 & ~a9556;
assign a9658 = ~a9612 & a9570;
assign a9660 = ~a9612 & a9574;
assign a9662 = ~a9612 & a9578;
assign a9664 = ~a9662 & ~a9660;
assign a9666 = a9664 & ~a9658;
assign a9668 = a9666 & ~a9656;
assign a9670 = a9668 & ~a9558;
assign a9672 = a9670 & ~a9562;
assign a9674 = a9672 & ~a9566;
assign a9676 = ~a9674 & a6596;
assign a9678 = ~a9598 & ~a9450;
assign a9680 = ~a9678 & a9602;
assign a9682 = ~a9680 & ~a9436;
assign a9684 = ~a9602 & ~a9442;
assign a9686 = ~a9684 & a9450;
assign a9688 = ~a9686 & a9438;
assign a9690 = ~a9686 & a9458;
assign a9692 = ~a9686 & a9462;
assign a9694 = ~a9692 & ~a9690;
assign a9696 = a9694 & ~a9688;
assign a9698 = a9696 & ~a9682;
assign a9700 = a9698 & ~a9466;
assign a9702 = a9700 & ~a9478;
assign a9704 = a9702 & ~a9482;
assign a9706 = ~a9704 & a6258;
assign a9708 = ~a9680 & ~a9508;
assign a9710 = ~a9686 & a9510;
assign a9712 = ~a9686 & a9514;
assign a9714 = ~a9686 & a9518;
assign a9716 = ~a9714 & ~a9712;
assign a9718 = a9716 & ~a9710;
assign a9720 = a9718 & ~a9708;
assign a9722 = a9720 & ~a9522;
assign a9724 = a9722 & ~a9526;
assign a9726 = a9724 & ~a9530;
assign a9728 = ~a9726 & a6428;
assign a9730 = ~a9680 & ~a9556;
assign a9732 = ~a9686 & a9558;
assign a9734 = ~a9686 & a9562;
assign a9736 = ~a9686 & a9566;
assign a9738 = ~a9736 & ~a9734;
assign a9740 = a9738 & ~a9732;
assign a9742 = a9740 & ~a9730;
assign a9744 = a9742 & ~a9570;
assign a9746 = a9744 & ~a9574;
assign a9748 = a9746 & ~a9578;
assign a9750 = ~a9748 & a6598;
assign a9752 = ~a8372 & a6252;
assign a9754 = ~a8378 & a6422;
assign a9756 = ~a9754 & ~a9752;
assign a9758 = ~a8388 & a6592;
assign a9760 = ~a9758 & a9756;
assign a9762 = ~a8312 & a7272;
assign a9764 = ~a6426 & ~a6256;
assign a9766 = a9764 & ~a6596;
assign a9768 = ~a6428 & ~a6258;
assign a9770 = a9768 & ~a6598;
assign a9772 = ~a9770 & ~a9450;
assign a9774 = ~a9772 & a9766;
assign a9776 = ~a9774 & a9762;
assign a9778 = ~a8318 & a7442;
assign a9780 = a9778 & ~a9774;
assign a9782 = ~a8328 & a7612;
assign a9784 = a9782 & ~a9774;
assign a9786 = ~a8284 & a7782;
assign a9788 = ~a9766 & ~a9470;
assign a9790 = ~a9788 & a9770;
assign a9792 = ~a9790 & a9786;
assign a9794 = ~a8290 & a7952;
assign a9796 = a9794 & ~a9790;
assign a9798 = ~a8300 & a8122;
assign a9800 = a9798 & ~a9790;
assign a9802 = ~a9800 & ~a9796;
assign a9804 = a9802 & ~a9792;
assign a9806 = a9804 & ~a9784;
assign a9808 = a9806 & ~a9780;
assign a9810 = a9808 & ~a9776;
assign a9812 = a9810 & a9760;
assign a9814 = ~a9812 & a6758;
assign a9816 = ~a8488 & a6252;
assign a9818 = ~a8494 & a6422;
assign a9820 = ~a9818 & ~a9816;
assign a9822 = ~a8504 & a6592;
assign a9824 = ~a9822 & a9820;
assign a9826 = ~a8428 & a7272;
assign a9828 = a9826 & ~a9774;
assign a9830 = ~a8434 & a7442;
assign a9832 = a9830 & ~a9774;
assign a9834 = ~a8444 & a7612;
assign a9836 = a9834 & ~a9774;
assign a9838 = ~a8400 & a7782;
assign a9840 = a9838 & ~a9790;
assign a9842 = ~a8406 & a7952;
assign a9844 = a9842 & ~a9790;
assign a9846 = ~a8416 & a8122;
assign a9848 = a9846 & ~a9790;
assign a9850 = ~a9848 & ~a9844;
assign a9852 = a9850 & ~a9840;
assign a9854 = a9852 & ~a9836;
assign a9856 = a9854 & ~a9832;
assign a9858 = a9856 & ~a9828;
assign a9860 = a9858 & a9824;
assign a9862 = ~a9860 & a6928;
assign a9864 = ~a6268 & a6252;
assign a9866 = ~a6438 & a6422;
assign a9868 = ~a9866 & ~a9864;
assign a9870 = ~a6608 & a6592;
assign a9872 = ~a9870 & a9868;
assign a9874 = ~a7288 & a7272;
assign a9876 = a9874 & ~a9774;
assign a9878 = ~a7458 & a7442;
assign a9880 = a9878 & ~a9774;
assign a9882 = ~a7628 & a7612;
assign a9884 = a9882 & ~a9774;
assign a9886 = ~a7798 & a7782;
assign a9888 = a9886 & ~a9790;
assign a9890 = ~a7968 & a7952;
assign a9892 = a9890 & ~a9790;
assign a9894 = ~a8138 & a8122;
assign a9896 = a9894 & ~a9790;
assign a9898 = ~a9896 & ~a9892;
assign a9900 = a9898 & ~a9888;
assign a9902 = a9900 & ~a9884;
assign a9904 = a9902 & ~a9880;
assign a9906 = a9904 & ~a9876;
assign a9908 = a9906 & a9872;
assign a9910 = ~a9908 & a7098;
assign a9912 = ~a7438 & ~a7268;
assign a9914 = a9912 & ~a7608;
assign a9916 = ~a7948 & ~a7778;
assign a9918 = a9916 & ~a8118;
assign a9920 = ~a9918 & ~a9470;
assign a9922 = ~a9920 & a9914;
assign a9924 = ~a9922 & ~a9760;
assign a9926 = ~a9914 & ~a9770;
assign a9928 = ~a9926 & a9470;
assign a9930 = ~a9928 & a9786;
assign a9932 = ~a9928 & a9794;
assign a9934 = ~a9928 & a9798;
assign a9936 = ~a9934 & ~a9932;
assign a9938 = a9936 & ~a9930;
assign a9940 = a9938 & ~a9924;
assign a9942 = a9940 & ~a9762;
assign a9944 = a9942 & ~a9778;
assign a9946 = a9944 & ~a9782;
assign a9948 = ~a9946 & a6766;
assign a9950 = ~a9922 & ~a9824;
assign a9952 = ~a9928 & a9838;
assign a9954 = ~a9928 & a9842;
assign a9956 = ~a9928 & a9846;
assign a9958 = ~a9956 & ~a9954;
assign a9960 = a9958 & ~a9952;
assign a9962 = a9960 & ~a9950;
assign a9964 = a9962 & ~a9826;
assign a9966 = a9964 & ~a9830;
assign a9968 = a9966 & ~a9834;
assign a9970 = ~a9968 & a6936;
assign a9972 = ~a9922 & ~a9872;
assign a9974 = ~a9928 & a9886;
assign a9976 = ~a9928 & a9890;
assign a9978 = ~a9928 & a9894;
assign a9980 = ~a9978 & ~a9976;
assign a9982 = a9980 & ~a9974;
assign a9984 = a9982 & ~a9972;
assign a9986 = a9984 & ~a9874;
assign a9988 = a9986 & ~a9878;
assign a9990 = a9988 & ~a9882;
assign a9992 = ~a9990 & a7106;
assign a9994 = ~a9914 & ~a9450;
assign a9996 = ~a9994 & a9918;
assign a9998 = ~a9996 & ~a9760;
assign a10000 = ~a9918 & ~a9766;
assign a10002 = ~a10000 & a9450;
assign a10004 = ~a10002 & a9762;
assign a10006 = ~a10002 & a9778;
assign a10008 = ~a10002 & a9782;
assign a10010 = ~a10008 & ~a10006;
assign a10012 = a10010 & ~a10004;
assign a10014 = a10012 & ~a9998;
assign a10016 = a10014 & ~a9786;
assign a10018 = a10016 & ~a9794;
assign a10020 = a10018 & ~a9798;
assign a10022 = ~a10020 & a6768;
assign a10024 = ~a9996 & ~a9824;
assign a10026 = ~a10002 & a9826;
assign a10028 = ~a10002 & a9830;
assign a10030 = ~a10002 & a9834;
assign a10032 = ~a10030 & ~a10028;
assign a10034 = a10032 & ~a10026;
assign a10036 = a10034 & ~a10024;
assign a10038 = a10036 & ~a9838;
assign a10040 = a10038 & ~a9842;
assign a10042 = a10040 & ~a9846;
assign a10044 = ~a10042 & a6938;
assign a10046 = ~a9996 & ~a9872;
assign a10048 = ~a10002 & a9874;
assign a10050 = ~a10002 & a9878;
assign a10052 = ~a10002 & a9882;
assign a10054 = ~a10052 & ~a10050;
assign a10056 = a10054 & ~a10048;
assign a10058 = a10056 & ~a10046;
assign a10060 = a10058 & ~a9886;
assign a10062 = a10060 & ~a9890;
assign a10064 = a10062 & ~a9894;
assign a10066 = ~a10064 & a7108;
assign a10068 = ~a8372 & a6256;
assign a10070 = ~a8378 & a6426;
assign a10072 = ~a10070 & ~a10068;
assign a10074 = ~a8388 & a6596;
assign a10076 = ~a10074 & a10072;
assign a10078 = ~a8342 & a6766;
assign a10080 = ~a6422 & ~a6252;
assign a10082 = a10080 & ~a6592;
assign a10084 = ~a9770 & ~a9602;
assign a10086 = ~a10084 & a10082;
assign a10088 = ~a10086 & a10078;
assign a10090 = ~a8348 & a6936;
assign a10092 = a10090 & ~a10086;
assign a10094 = ~a8358 & a7106;
assign a10096 = a10094 & ~a10086;
assign a10098 = ~a8284 & a7786;
assign a10100 = ~a10082 & ~a9446;
assign a10102 = ~a10100 & a9770;
assign a10104 = ~a10102 & a10098;
assign a10106 = ~a8290 & a7956;
assign a10108 = a10106 & ~a10102;
assign a10110 = ~a8300 & a8126;
assign a10112 = a10110 & ~a10102;
assign a10114 = ~a10112 & ~a10108;
assign a10116 = a10114 & ~a10104;
assign a10118 = a10116 & ~a10096;
assign a10120 = a10118 & ~a10092;
assign a10122 = a10120 & ~a10088;
assign a10124 = a10122 & a10076;
assign a10126 = ~a10124 & a7268;
assign a10128 = ~a8488 & a6256;
assign a10130 = ~a8494 & a6426;
assign a10132 = ~a10130 & ~a10128;
assign a10134 = ~a8504 & a6596;
assign a10136 = ~a10134 & a10132;
assign a10138 = ~a8458 & a6766;
assign a10140 = a10138 & ~a10086;
assign a10142 = ~a8464 & a6936;
assign a10144 = a10142 & ~a10086;
assign a10146 = ~a8474 & a7106;
assign a10148 = a10146 & ~a10086;
assign a10150 = ~a8400 & a7786;
assign a10152 = a10150 & ~a10102;
assign a10154 = ~a8406 & a7956;
assign a10156 = a10154 & ~a10102;
assign a10158 = ~a8416 & a8126;
assign a10160 = a10158 & ~a10102;
assign a10162 = ~a10160 & ~a10156;
assign a10164 = a10162 & ~a10152;
assign a10166 = a10164 & ~a10148;
assign a10168 = a10166 & ~a10144;
assign a10170 = a10168 & ~a10140;
assign a10172 = a10170 & a10136;
assign a10174 = ~a10172 & a7438;
assign a10176 = ~a6268 & a6256;
assign a10178 = ~a6438 & a6426;
assign a10180 = ~a10178 & ~a10176;
assign a10182 = ~a6608 & a6596;
assign a10184 = ~a10182 & a10180;
assign a10186 = ~a6778 & a6766;
assign a10188 = a10186 & ~a10086;
assign a10190 = ~a6948 & a6936;
assign a10192 = a10190 & ~a10086;
assign a10194 = ~a7118 & a7106;
assign a10196 = a10194 & ~a10086;
assign a10198 = ~a7798 & a7786;
assign a10200 = a10198 & ~a10102;
assign a10202 = ~a7968 & a7956;
assign a10204 = a10202 & ~a10102;
assign a10206 = ~a8138 & a8126;
assign a10208 = a10206 & ~a10102;
assign a10210 = ~a10208 & ~a10204;
assign a10212 = a10210 & ~a10200;
assign a10214 = a10212 & ~a10196;
assign a10216 = a10214 & ~a10192;
assign a10218 = a10216 & ~a10188;
assign a10220 = a10218 & a10184;
assign a10222 = ~a10220 & a7608;
assign a10224 = ~a6928 & ~a6758;
assign a10226 = a10224 & ~a7098;
assign a10228 = ~a9918 & ~a9446;
assign a10230 = ~a10228 & a10226;
assign a10232 = ~a10230 & ~a10076;
assign a10234 = ~a10226 & ~a9770;
assign a10236 = ~a10234 & a9446;
assign a10238 = ~a10236 & a10098;
assign a10240 = ~a10236 & a10106;
assign a10242 = ~a10236 & a10110;
assign a10244 = ~a10242 & ~a10240;
assign a10246 = a10244 & ~a10238;
assign a10248 = a10246 & ~a10232;
assign a10250 = a10248 & ~a10078;
assign a10252 = a10250 & ~a10090;
assign a10254 = a10252 & ~a10094;
assign a10256 = ~a10254 & a7272;
assign a10258 = ~a10230 & ~a10136;
assign a10260 = ~a10236 & a10150;
assign a10262 = ~a10236 & a10154;
assign a10264 = ~a10236 & a10158;
assign a10266 = ~a10264 & ~a10262;
assign a10268 = a10266 & ~a10260;
assign a10270 = a10268 & ~a10258;
assign a10272 = a10270 & ~a10138;
assign a10274 = a10272 & ~a10142;
assign a10276 = a10274 & ~a10146;
assign a10278 = ~a10276 & a7442;
assign a10280 = ~a10230 & ~a10184;
assign a10282 = ~a10236 & a10198;
assign a10284 = ~a10236 & a10202;
assign a10286 = ~a10236 & a10206;
assign a10288 = ~a10286 & ~a10284;
assign a10290 = a10288 & ~a10282;
assign a10292 = a10290 & ~a10280;
assign a10294 = a10292 & ~a10186;
assign a10296 = a10294 & ~a10190;
assign a10298 = a10296 & ~a10194;
assign a10300 = ~a10298 & a7612;
assign a10302 = ~a10226 & ~a9602;
assign a10304 = ~a10302 & a9918;
assign a10306 = ~a10304 & ~a10076;
assign a10308 = ~a10082 & ~a9918;
assign a10310 = ~a10308 & a9602;
assign a10312 = ~a10310 & a10078;
assign a10314 = ~a10310 & a10090;
assign a10316 = ~a10310 & a10094;
assign a10318 = ~a10316 & ~a10314;
assign a10320 = a10318 & ~a10312;
assign a10322 = a10320 & ~a10306;
assign a10324 = a10322 & ~a10098;
assign a10326 = a10324 & ~a10106;
assign a10328 = a10326 & ~a10110;
assign a10330 = ~a10328 & a7278;
assign a10332 = ~a10304 & ~a10136;
assign a10334 = ~a10310 & a10138;
assign a10336 = ~a10310 & a10142;
assign a10338 = ~a10310 & a10146;
assign a10340 = ~a10338 & ~a10336;
assign a10342 = a10340 & ~a10334;
assign a10344 = a10342 & ~a10332;
assign a10346 = a10344 & ~a10150;
assign a10348 = a10346 & ~a10154;
assign a10350 = a10348 & ~a10158;
assign a10352 = ~a10350 & a7448;
assign a10354 = ~a10304 & ~a10184;
assign a10356 = ~a10310 & a10186;
assign a10358 = ~a10310 & a10190;
assign a10360 = ~a10310 & a10194;
assign a10362 = ~a10360 & ~a10358;
assign a10364 = a10362 & ~a10356;
assign a10366 = a10364 & ~a10354;
assign a10368 = a10366 & ~a10198;
assign a10370 = a10368 & ~a10202;
assign a10372 = a10370 & ~a10206;
assign a10374 = ~a10372 & a7618;
assign a10376 = ~a8372 & a6258;
assign a10378 = ~a8378 & a6428;
assign a10380 = ~a10378 & ~a10376;
assign a10382 = ~a8388 & a6598;
assign a10384 = ~a10382 & a10380;
assign a10386 = ~a8342 & a6768;
assign a10388 = ~a9766 & ~a9598;
assign a10390 = ~a10388 & a10082;
assign a10392 = ~a10390 & a10386;
assign a10394 = ~a8348 & a6938;
assign a10396 = a10394 & ~a10390;
assign a10398 = ~a8358 & a7108;
assign a10400 = a10398 & ~a10390;
assign a10402 = ~a8312 & a7278;
assign a10404 = ~a10082 & ~a9442;
assign a10406 = ~a10404 & a9766;
assign a10408 = ~a10406 & a10402;
assign a10410 = ~a8318 & a7448;
assign a10412 = a10410 & ~a10406;
assign a10414 = ~a8328 & a7618;
assign a10416 = a10414 & ~a10406;
assign a10418 = ~a10416 & ~a10412;
assign a10420 = a10418 & ~a10408;
assign a10422 = a10420 & ~a10400;
assign a10424 = a10422 & ~a10396;
assign a10426 = a10424 & ~a10392;
assign a10428 = a10426 & a10384;
assign a10430 = ~a10428 & a7778;
assign a10432 = ~a8488 & a6258;
assign a10434 = ~a8494 & a6428;
assign a10436 = ~a10434 & ~a10432;
assign a10438 = ~a8504 & a6598;
assign a10440 = ~a10438 & a10436;
assign a10442 = ~a8458 & a6768;
assign a10444 = a10442 & ~a10390;
assign a10446 = ~a8464 & a6938;
assign a10448 = a10446 & ~a10390;
assign a10450 = ~a8474 & a7108;
assign a10452 = a10450 & ~a10390;
assign a10454 = ~a8428 & a7278;
assign a10456 = a10454 & ~a10406;
assign a10458 = ~a8434 & a7448;
assign a10460 = a10458 & ~a10406;
assign a10462 = ~a8444 & a7618;
assign a10464 = a10462 & ~a10406;
assign a10466 = ~a10464 & ~a10460;
assign a10468 = a10466 & ~a10456;
assign a10470 = a10468 & ~a10452;
assign a10472 = a10470 & ~a10448;
assign a10474 = a10472 & ~a10444;
assign a10476 = a10474 & a10440;
assign a10478 = ~a10476 & a7948;
assign a10480 = ~a6268 & a6258;
assign a10482 = ~a6438 & a6428;
assign a10484 = ~a10482 & ~a10480;
assign a10486 = ~a6608 & a6598;
assign a10488 = ~a10486 & a10484;
assign a10490 = ~a6778 & a6768;
assign a10492 = a10490 & ~a10390;
assign a10494 = ~a6948 & a6938;
assign a10496 = a10494 & ~a10390;
assign a10498 = ~a7118 & a7108;
assign a10500 = a10498 & ~a10390;
assign a10502 = ~a7288 & a7278;
assign a10504 = a10502 & ~a10406;
assign a10506 = ~a7458 & a7448;
assign a10508 = a10506 & ~a10406;
assign a10510 = ~a7628 & a7618;
assign a10512 = a10510 & ~a10406;
assign a10514 = ~a10512 & ~a10508;
assign a10516 = a10514 & ~a10504;
assign a10518 = a10516 & ~a10500;
assign a10520 = a10518 & ~a10496;
assign a10522 = a10520 & ~a10492;
assign a10524 = a10522 & a10488;
assign a10526 = ~a10524 & a8118;
assign a10528 = ~a9914 & ~a9442;
assign a10530 = ~a10528 & a10226;
assign a10532 = ~a10530 & ~a10384;
assign a10534 = ~a10226 & ~a9766;
assign a10536 = ~a10534 & a9442;
assign a10538 = ~a10536 & a10402;
assign a10540 = ~a10536 & a10410;
assign a10542 = ~a10536 & a10414;
assign a10544 = ~a10542 & ~a10540;
assign a10546 = a10544 & ~a10538;
assign a10548 = a10546 & ~a10532;
assign a10550 = a10548 & ~a10386;
assign a10552 = a10550 & ~a10394;
assign a10554 = a10552 & ~a10398;
assign a10556 = ~a10554 & a7782;
assign a10558 = ~a10530 & ~a10440;
assign a10560 = ~a10536 & a10454;
assign a10562 = ~a10536 & a10458;
assign a10564 = ~a10536 & a10462;
assign a10566 = ~a10564 & ~a10562;
assign a10568 = a10566 & ~a10560;
assign a10570 = a10568 & ~a10558;
assign a10572 = a10570 & ~a10442;
assign a10574 = a10572 & ~a10446;
assign a10576 = a10574 & ~a10450;
assign a10578 = ~a10576 & a7952;
assign a10580 = ~a10530 & ~a10488;
assign a10582 = ~a10536 & a10502;
assign a10584 = ~a10536 & a10506;
assign a10586 = ~a10536 & a10510;
assign a10588 = ~a10586 & ~a10584;
assign a10590 = a10588 & ~a10582;
assign a10592 = a10590 & ~a10580;
assign a10594 = a10592 & ~a10490;
assign a10596 = a10594 & ~a10494;
assign a10598 = a10596 & ~a10498;
assign a10600 = ~a10598 & a8122;
assign a10602 = ~a10226 & ~a9598;
assign a10604 = ~a10602 & a9914;
assign a10606 = ~a10604 & ~a10384;
assign a10608 = ~a10082 & ~a9914;
assign a10610 = ~a10608 & a9598;
assign a10612 = ~a10610 & a10386;
assign a10614 = ~a10610 & a10394;
assign a10616 = ~a10610 & a10398;
assign a10618 = ~a10616 & ~a10614;
assign a10620 = a10618 & ~a10612;
assign a10622 = a10620 & ~a10606;
assign a10624 = a10622 & ~a10402;
assign a10626 = a10624 & ~a10410;
assign a10628 = a10626 & ~a10414;
assign a10630 = ~a10628 & a7786;
assign a10632 = ~a10604 & ~a10440;
assign a10634 = ~a10610 & a10442;
assign a10636 = ~a10610 & a10446;
assign a10638 = ~a10610 & a10450;
assign a10640 = ~a10638 & ~a10636;
assign a10642 = a10640 & ~a10634;
assign a10644 = a10642 & ~a10632;
assign a10646 = a10644 & ~a10454;
assign a10648 = a10646 & ~a10458;
assign a10650 = a10648 & ~a10462;
assign a10652 = ~a10650 & a7956;
assign a10654 = ~a10604 & ~a10488;
assign a10656 = ~a10610 & a10490;
assign a10658 = ~a10610 & a10494;
assign a10660 = ~a10610 & a10498;
assign a10662 = ~a10660 & ~a10658;
assign a10664 = a10662 & ~a10656;
assign a10666 = a10664 & ~a10654;
assign a10668 = a10666 & ~a10502;
assign a10670 = a10668 & ~a10506;
assign a10672 = a10670 & ~a10510;
assign a10674 = ~a10672 & a8126;
assign a10676 = ~a9766 & a9604;
assign a10678 = ~a9770 & a9678;
assign a10680 = ~a10678 & ~a10676;
assign a10682 = a10680 & ~a10388;
assign a10684 = a10682 & ~a10084;
assign a10686 = a10684 & a10082;
assign a10688 = ~a10226 & a9772;
assign a10690 = a10000 & ~a9446;
assign a10692 = ~a10690 & ~a10688;
assign a10694 = a10692 & ~a10534;
assign a10696 = a10694 & ~a9452;
assign a10698 = a10696 & a9442;
assign a10700 = a10100 & ~a9914;
assign a10702 = a10234 & ~a9598;
assign a10704 = ~a10702 & ~a10700;
assign a10706 = a10704 & ~a9926;
assign a10708 = a10706 & ~a9610;
assign a10710 = a10708 & a9470;
assign a10712 = a6244 & l604;
assign a10714 = ~a6244 & ~l604;
assign a10716 = ~a10714 & ~a10712;
assign a10718 = a6414 & l618;
assign a10720 = ~a6414 & ~l618;
assign a10722 = ~a10720 & ~a10718;
assign a10724 = a6584 & l632;
assign a10726 = ~a6584 & ~l632;
assign a10728 = ~a10726 & ~a10724;
assign a10730 = a6754 & l672;
assign a10732 = ~a6754 & ~l672;
assign a10734 = ~a10732 & ~a10730;
assign a10736 = a6924 & l686;
assign a10738 = ~a6924 & ~l686;
assign a10740 = ~a10738 & ~a10736;
assign a10742 = a7094 & l700;
assign a10744 = ~a7094 & ~l700;
assign a10746 = ~a10744 & ~a10742;
assign a10748 = a7264 & l740;
assign a10750 = ~a7264 & ~l740;
assign a10752 = ~a10750 & ~a10748;
assign a10754 = a7434 & l754;
assign a10756 = ~a7434 & ~l754;
assign a10758 = ~a10756 & ~a10754;
assign a10760 = a7604 & l768;
assign a10762 = ~a7604 & ~l768;
assign a10764 = ~a10762 & ~a10760;
assign a10766 = a7774 & l808;
assign a10768 = ~a7774 & ~l808;
assign a10770 = ~a10768 & ~a10766;
assign a10772 = a7944 & l822;
assign a10774 = ~a7944 & ~l822;
assign a10776 = ~a10774 & ~a10772;
assign a10778 = a8114 & l836;
assign a10780 = ~a8114 & ~l836;
assign a10782 = ~a10780 & ~a10778;
assign a10784 = ~l878 & ~l602;
assign a10786 = l878 & l602;
assign a10788 = ~a10786 & ~a10784;
assign a10790 = ~l876 & l600;
assign a10792 = l876 & ~l600;
assign a10794 = ~a10792 & ~a10790;
assign a10796 = ~l882 & ~l608;
assign a10798 = l882 & l608;
assign a10800 = ~a10798 & ~a10796;
assign a10802 = ~l880 & l606;
assign a10804 = l880 & ~l606;
assign a10806 = ~a10804 & ~a10802;
assign a10808 = ~l886 & ~l616;
assign a10810 = l886 & l616;
assign a10812 = ~a10810 & ~a10808;
assign a10814 = ~l884 & l614;
assign a10816 = l884 & ~l614;
assign a10818 = ~a10816 & ~a10814;
assign a10820 = ~l890 & ~l622;
assign a10822 = l890 & l622;
assign a10824 = ~a10822 & ~a10820;
assign a10826 = ~l888 & l620;
assign a10828 = l888 & ~l620;
assign a10830 = ~a10828 & ~a10826;
assign a10832 = ~l894 & ~l630;
assign a10834 = l894 & l630;
assign a10836 = ~a10834 & ~a10832;
assign a10838 = ~l892 & l628;
assign a10840 = l892 & ~l628;
assign a10842 = ~a10840 & ~a10838;
assign a10844 = ~l898 & ~l636;
assign a10846 = l898 & l636;
assign a10848 = ~a10846 & ~a10844;
assign a10850 = ~l896 & l634;
assign a10852 = l896 & ~l634;
assign a10854 = ~a10852 & ~a10850;
assign a10856 = ~l904 & ~l642;
assign a10858 = l904 & l642;
assign a10860 = ~a10858 & ~a10856;
assign a10862 = ~l902 & l640;
assign a10864 = l902 & ~l640;
assign a10866 = ~a10864 & ~a10862;
assign a10868 = ~l900 & l638;
assign a10870 = l900 & ~l638;
assign a10872 = ~a10870 & ~a10868;
assign a10874 = ~l906 & l644;
assign a10876 = l906 & ~l644;
assign a10878 = ~a10876 & ~a10874;
assign a10880 = ~l910 & l648;
assign a10882 = l910 & ~l648;
assign a10884 = ~a10882 & ~a10880;
assign a10886 = ~l908 & l646;
assign a10888 = l908 & ~l646;
assign a10890 = ~a10888 & ~a10886;
assign a10892 = ~l912 & l652;
assign a10894 = l912 & ~l652;
assign a10896 = ~a10894 & ~a10892;
assign a10898 = ~l914 & l654;
assign a10900 = l914 & ~l654;
assign a10902 = ~a10900 & ~a10898;
assign a10904 = ~l922 & l662;
assign a10906 = l922 & ~l662;
assign a10908 = ~a10906 & ~a10904;
assign a10910 = ~l920 & l660;
assign a10912 = l920 & ~l660;
assign a10914 = ~a10912 & ~a10910;
assign a10916 = ~l918 & l658;
assign a10918 = l918 & ~l658;
assign a10920 = ~a10918 & ~a10916;
assign a10922 = ~l916 & l656;
assign a10924 = l916 & ~l656;
assign a10926 = ~a10924 & ~a10922;
assign a10928 = ~l926 & ~l670;
assign a10930 = l926 & l670;
assign a10932 = ~a10930 & ~a10928;
assign a10934 = ~l924 & l668;
assign a10936 = l924 & ~l668;
assign a10938 = ~a10936 & ~a10934;
assign a10940 = ~l930 & ~l676;
assign a10942 = l930 & l676;
assign a10944 = ~a10942 & ~a10940;
assign a10946 = ~l928 & l674;
assign a10948 = l928 & ~l674;
assign a10950 = ~a10948 & ~a10946;
assign a10952 = ~l934 & ~l684;
assign a10954 = l934 & l684;
assign a10956 = ~a10954 & ~a10952;
assign a10958 = ~l932 & l682;
assign a10960 = l932 & ~l682;
assign a10962 = ~a10960 & ~a10958;
assign a10964 = ~l938 & ~l690;
assign a10966 = l938 & l690;
assign a10968 = ~a10966 & ~a10964;
assign a10970 = ~l936 & l688;
assign a10972 = l936 & ~l688;
assign a10974 = ~a10972 & ~a10970;
assign a10976 = ~l942 & ~l698;
assign a10978 = l942 & l698;
assign a10980 = ~a10978 & ~a10976;
assign a10982 = ~l940 & l696;
assign a10984 = l940 & ~l696;
assign a10986 = ~a10984 & ~a10982;
assign a10988 = ~l946 & ~l704;
assign a10990 = l946 & l704;
assign a10992 = ~a10990 & ~a10988;
assign a10994 = ~l944 & l702;
assign a10996 = l944 & ~l702;
assign a10998 = ~a10996 & ~a10994;
assign a11000 = ~l952 & ~l710;
assign a11002 = l952 & l710;
assign a11004 = ~a11002 & ~a11000;
assign a11006 = ~l950 & l708;
assign a11008 = l950 & ~l708;
assign a11010 = ~a11008 & ~a11006;
assign a11012 = ~l948 & l706;
assign a11014 = l948 & ~l706;
assign a11016 = ~a11014 & ~a11012;
assign a11018 = ~l954 & l712;
assign a11020 = l954 & ~l712;
assign a11022 = ~a11020 & ~a11018;
assign a11024 = ~l958 & l716;
assign a11026 = l958 & ~l716;
assign a11028 = ~a11026 & ~a11024;
assign a11030 = ~l956 & l714;
assign a11032 = l956 & ~l714;
assign a11034 = ~a11032 & ~a11030;
assign a11036 = ~l960 & l720;
assign a11038 = l960 & ~l720;
assign a11040 = ~a11038 & ~a11036;
assign a11042 = ~l962 & l722;
assign a11044 = l962 & ~l722;
assign a11046 = ~a11044 & ~a11042;
assign a11048 = ~l970 & l730;
assign a11050 = l970 & ~l730;
assign a11052 = ~a11050 & ~a11048;
assign a11054 = ~l968 & l728;
assign a11056 = l968 & ~l728;
assign a11058 = ~a11056 & ~a11054;
assign a11060 = ~l966 & l726;
assign a11062 = l966 & ~l726;
assign a11064 = ~a11062 & ~a11060;
assign a11066 = ~l964 & l724;
assign a11068 = l964 & ~l724;
assign a11070 = ~a11068 & ~a11066;
assign a11072 = ~l974 & ~l738;
assign a11074 = l974 & l738;
assign a11076 = ~a11074 & ~a11072;
assign a11078 = ~l972 & l736;
assign a11080 = l972 & ~l736;
assign a11082 = ~a11080 & ~a11078;
assign a11084 = ~l978 & ~l744;
assign a11086 = l978 & l744;
assign a11088 = ~a11086 & ~a11084;
assign a11090 = ~l976 & l742;
assign a11092 = l976 & ~l742;
assign a11094 = ~a11092 & ~a11090;
assign a11096 = ~l982 & ~l752;
assign a11098 = l982 & l752;
assign a11100 = ~a11098 & ~a11096;
assign a11102 = ~l980 & l750;
assign a11104 = l980 & ~l750;
assign a11106 = ~a11104 & ~a11102;
assign a11108 = ~l986 & ~l758;
assign a11110 = l986 & l758;
assign a11112 = ~a11110 & ~a11108;
assign a11114 = ~l984 & l756;
assign a11116 = l984 & ~l756;
assign a11118 = ~a11116 & ~a11114;
assign a11120 = ~l990 & ~l766;
assign a11122 = l990 & l766;
assign a11124 = ~a11122 & ~a11120;
assign a11126 = ~l988 & l764;
assign a11128 = l988 & ~l764;
assign a11130 = ~a11128 & ~a11126;
assign a11132 = ~l994 & ~l772;
assign a11134 = l994 & l772;
assign a11136 = ~a11134 & ~a11132;
assign a11138 = ~l992 & l770;
assign a11140 = l992 & ~l770;
assign a11142 = ~a11140 & ~a11138;
assign a11144 = ~l1000 & ~l778;
assign a11146 = l1000 & l778;
assign a11148 = ~a11146 & ~a11144;
assign a11150 = ~l998 & l776;
assign a11152 = l998 & ~l776;
assign a11154 = ~a11152 & ~a11150;
assign a11156 = ~l996 & l774;
assign a11158 = l996 & ~l774;
assign a11160 = ~a11158 & ~a11156;
assign a11162 = ~l1002 & l780;
assign a11164 = l1002 & ~l780;
assign a11166 = ~a11164 & ~a11162;
assign a11168 = ~l1006 & l784;
assign a11170 = l1006 & ~l784;
assign a11172 = ~a11170 & ~a11168;
assign a11174 = ~l1004 & l782;
assign a11176 = l1004 & ~l782;
assign a11178 = ~a11176 & ~a11174;
assign a11180 = ~l1008 & l788;
assign a11182 = l1008 & ~l788;
assign a11184 = ~a11182 & ~a11180;
assign a11186 = ~l1010 & l790;
assign a11188 = l1010 & ~l790;
assign a11190 = ~a11188 & ~a11186;
assign a11192 = ~l1018 & l798;
assign a11194 = l1018 & ~l798;
assign a11196 = ~a11194 & ~a11192;
assign a11198 = ~l1016 & l796;
assign a11200 = l1016 & ~l796;
assign a11202 = ~a11200 & ~a11198;
assign a11204 = ~l1014 & l794;
assign a11206 = l1014 & ~l794;
assign a11208 = ~a11206 & ~a11204;
assign a11210 = ~l1012 & l792;
assign a11212 = l1012 & ~l792;
assign a11214 = ~a11212 & ~a11210;
assign a11216 = ~l1022 & ~l806;
assign a11218 = l1022 & l806;
assign a11220 = ~a11218 & ~a11216;
assign a11222 = ~l1020 & l804;
assign a11224 = l1020 & ~l804;
assign a11226 = ~a11224 & ~a11222;
assign a11228 = ~l1026 & ~l812;
assign a11230 = l1026 & l812;
assign a11232 = ~a11230 & ~a11228;
assign a11234 = ~l1024 & l810;
assign a11236 = l1024 & ~l810;
assign a11238 = ~a11236 & ~a11234;
assign a11240 = ~l1030 & ~l820;
assign a11242 = l1030 & l820;
assign a11244 = ~a11242 & ~a11240;
assign a11246 = ~l1028 & l818;
assign a11248 = l1028 & ~l818;
assign a11250 = ~a11248 & ~a11246;
assign a11252 = ~l1034 & ~l826;
assign a11254 = l1034 & l826;
assign a11256 = ~a11254 & ~a11252;
assign a11258 = ~l1032 & l824;
assign a11260 = l1032 & ~l824;
assign a11262 = ~a11260 & ~a11258;
assign a11264 = ~l1038 & ~l834;
assign a11266 = l1038 & l834;
assign a11268 = ~a11266 & ~a11264;
assign a11270 = ~l1036 & l832;
assign a11272 = l1036 & ~l832;
assign a11274 = ~a11272 & ~a11270;
assign a11276 = ~l1042 & ~l840;
assign a11278 = l1042 & l840;
assign a11280 = ~a11278 & ~a11276;
assign a11282 = ~l1040 & l838;
assign a11284 = l1040 & ~l838;
assign a11286 = ~a11284 & ~a11282;
assign a11288 = ~l1046 & l844;
assign a11290 = l1046 & ~l844;
assign a11292 = ~a11290 & ~a11288;
assign a11294 = ~l1044 & l842;
assign a11296 = l1044 & ~l842;
assign a11298 = ~a11296 & ~a11294;
assign a11300 = ~l1050 & l848;
assign a11302 = l1050 & ~l848;
assign a11304 = ~a11302 & ~a11300;
assign a11306 = ~l1054 & l852;
assign a11308 = l1054 & ~l852;
assign a11310 = ~a11308 & ~a11306;
assign a11312 = ~l1052 & l850;
assign a11314 = l1052 & ~l850;
assign a11316 = ~a11314 & ~a11312;
assign a11318 = ~l1056 & l856;
assign a11320 = l1056 & ~l856;
assign a11322 = ~a11320 & ~a11318;
assign a11324 = ~l1058 & l858;
assign a11326 = l1058 & ~l858;
assign a11328 = ~a11326 & ~a11324;
assign a11330 = ~l1066 & l866;
assign a11332 = l1066 & ~l866;
assign a11334 = ~a11332 & ~a11330;
assign a11336 = ~l1064 & l864;
assign a11338 = l1064 & ~l864;
assign a11340 = ~a11338 & ~a11336;
assign a11342 = ~l1062 & l862;
assign a11344 = l1062 & ~l862;
assign a11346 = ~a11344 & ~a11342;
assign a11348 = ~l1060 & l860;
assign a11350 = l1060 & ~l860;
assign a11352 = ~a11350 & ~a11348;
assign a11354 = ~l1068 & l868;
assign a11356 = l1068 & ~l868;
assign a11358 = ~a11356 & ~a11354;
assign a11360 = l1070 & ~l870;
assign a11362 = ~l1070 & l870;
assign a11364 = ~a11362 & ~a11360;
assign a11366 = l1072 & ~l872;
assign a11368 = ~l1072 & l872;
assign a11370 = ~a11368 & ~a11366;
assign a11372 = l1074 & ~l874;
assign a11374 = ~l1074 & l874;
assign a11376 = ~a11374 & ~a11372;
assign a11378 = a11376 & a11370;
assign a11380 = a11378 & a11364;
assign a11382 = a11380 & a11358;
assign a11384 = a11382 & a11352;
assign a11386 = a11384 & a11346;
assign a11388 = a11386 & a11340;
assign a11390 = a11388 & a11334;
assign a11392 = a11390 & a11328;
assign a11394 = a11392 & a11322;
assign a11396 = a11394 & a11316;
assign a11398 = a11396 & a11310;
assign a11400 = a11398 & a11304;
assign a11402 = a11400 & a11298;
assign a11404 = a11402 & a11292;
assign a11406 = ~l1048 & ~l846;
assign a11408 = l1048 & l846;
assign a11410 = ~a11408 & ~a11406;
assign a11412 = a11410 & a11404;
assign a11414 = a11412 & a11286;
assign a11416 = a11414 & a11280;
assign a11418 = a11416 & a11274;
assign a11420 = a11418 & a11268;
assign a11422 = a11420 & a11262;
assign a11424 = a11422 & a11256;
assign a11426 = a11424 & a11250;
assign a11428 = a11426 & a11244;
assign a11430 = a11428 & a11238;
assign a11432 = a11430 & a11232;
assign a11434 = a11432 & a11226;
assign a11436 = a11434 & a11220;
assign a11438 = a11436 & a11214;
assign a11440 = a11438 & a11208;
assign a11442 = a11440 & a11202;
assign a11444 = a11442 & a11196;
assign a11446 = a11444 & a11190;
assign a11448 = a11446 & a11184;
assign a11450 = a11448 & a11178;
assign a11452 = a11450 & a11172;
assign a11454 = a11452 & a11166;
assign a11456 = a11454 & a11160;
assign a11458 = a11456 & a11154;
assign a11460 = a11458 & a11148;
assign a11462 = a11460 & a11142;
assign a11464 = a11462 & a11136;
assign a11466 = a11464 & a11130;
assign a11468 = a11466 & a11124;
assign a11470 = a11468 & a11118;
assign a11472 = a11470 & a11112;
assign a11474 = a11472 & a11106;
assign a11476 = a11474 & a11100;
assign a11478 = a11476 & a11094;
assign a11480 = a11478 & a11088;
assign a11482 = a11480 & a11082;
assign a11484 = a11482 & a11076;
assign a11486 = a11484 & a11070;
assign a11488 = a11486 & a11064;
assign a11490 = a11488 & a11058;
assign a11492 = a11490 & a11052;
assign a11494 = a11492 & a11046;
assign a11496 = a11494 & a11040;
assign a11498 = a11496 & a11034;
assign a11500 = a11498 & a11028;
assign a11502 = a11500 & a11022;
assign a11504 = a11502 & a11016;
assign a11506 = a11504 & a11010;
assign a11508 = a11506 & a11004;
assign a11510 = a11508 & a10998;
assign a11512 = a11510 & a10992;
assign a11514 = a11512 & a10986;
assign a11516 = a11514 & a10980;
assign a11518 = a11516 & a10974;
assign a11520 = a11518 & a10968;
assign a11522 = a11520 & a10962;
assign a11524 = a11522 & a10956;
assign a11526 = a11524 & a10950;
assign a11528 = a11526 & a10944;
assign a11530 = a11528 & a10938;
assign a11532 = a11530 & a10932;
assign a11534 = a11532 & a10926;
assign a11536 = a11534 & a10920;
assign a11538 = a11536 & a10914;
assign a11540 = a11538 & a10908;
assign a11542 = a11540 & a10902;
assign a11544 = a11542 & a10896;
assign a11546 = a11544 & a10890;
assign a11548 = a11546 & a10884;
assign a11550 = a11548 & a10878;
assign a11552 = a11550 & a10872;
assign a11554 = a11552 & a10866;
assign a11556 = a11554 & a10860;
assign a11558 = a11556 & a10854;
assign a11560 = a11558 & a10848;
assign a11562 = a11560 & a10842;
assign a11564 = a11562 & a10836;
assign a11566 = a11564 & a10830;
assign a11568 = a11566 & a10824;
assign a11570 = a11568 & a10818;
assign a11572 = a11570 & a10812;
assign a11574 = a11572 & a10806;
assign a11576 = a11574 & a10800;
assign a11578 = a11576 & a10794;
assign a11580 = a11578 & a10788;
assign a11582 = a11580 & l1084;
assign a11584 = a11582 & l1076;
assign a11586 = a11584 & l1078;
assign a11588 = a11586 & l1080;
assign a11590 = ~a11588 & i466;
assign a11592 = ~a11590 & a10782;
assign a11594 = a11592 & a10776;
assign a11596 = a11594 & a10770;
assign a11598 = a11596 & a10764;
assign a11600 = a11598 & a10758;
assign a11602 = a11600 & a10752;
assign a11604 = a11602 & a10746;
assign a11606 = a11604 & a10740;
assign a11608 = a11606 & a10734;
assign a11610 = a11608 & a10728;
assign a11612 = a11610 & a10722;
assign a11614 = a11612 & a10716;
assign a11616 = a11614 & ~a10710;
assign a11618 = a11616 & ~a10698;
assign a11620 = a11618 & ~a10686;
assign a11622 = a11620 & ~a10674;
assign a11624 = a11622 & ~a10652;
assign a11626 = a11624 & ~a10630;
assign a11628 = a11626 & ~a10600;
assign a11630 = a11628 & ~a10578;
assign a11632 = a11630 & ~a10556;
assign a11634 = a11632 & ~a10526;
assign a11636 = a11634 & ~a10478;
assign a11638 = a11636 & ~a10430;
assign a11640 = a11638 & ~a10374;
assign a11642 = a11640 & ~a10352;
assign a11644 = a11642 & ~a10330;
assign a11646 = a11644 & ~a10300;
assign a11648 = a11646 & ~a10278;
assign a11650 = a11648 & ~a10256;
assign a11652 = a11650 & ~a10222;
assign a11654 = a11652 & ~a10174;
assign a11656 = a11654 & ~a10126;
assign a11658 = a11656 & ~a10066;
assign a11660 = a11658 & ~a10044;
assign a11662 = a11660 & ~a10022;
assign a11664 = a11662 & ~a9992;
assign a11666 = a11664 & ~a9970;
assign a11668 = a11666 & ~a9948;
assign a11670 = a11668 & ~a9910;
assign a11672 = a11670 & ~a9862;
assign a11674 = a11672 & ~a9814;
assign a11676 = a11674 & ~a9750;
assign a11678 = a11676 & ~a9728;
assign a11680 = a11678 & ~a9706;
assign a11682 = a11680 & ~a9676;
assign a11684 = a11682 & ~a9654;
assign a11686 = a11684 & ~a9632;
assign a11688 = a11686 & ~a9594;
assign a11690 = a11688 & ~a9546;
assign a11692 = a11690 & ~a9498;
assign a11694 = a11692 & a9426;
assign a11696 = a11694 & ~a8128;
assign a11698 = a11696 & a9336;
assign a11700 = a11698 & ~a7958;
assign a11702 = a11700 & a9244;
assign a11704 = a11702 & ~a7788;
assign a11706 = a11704 & a9152;
assign a11708 = a11706 & ~a7616;
assign a11710 = a11708 & a9062;
assign a11712 = a11710 & ~a7446;
assign a11714 = a11712 & a8970;
assign a11716 = a11714 & ~a7276;
assign a11718 = a11716 & a8878;
assign a11720 = a11718 & ~a7102;
assign a11722 = a11720 & a8788;
assign a11724 = a11722 & ~a6932;
assign a11726 = a11724 & a8696;
assign a11728 = a11726 & ~a6762;
assign a11730 = a11728 & a8604;
assign a11732 = a11730 & ~a6588;
assign a11734 = a11732 & a8514;
assign a11736 = a11734 & ~a6418;
assign a11738 = a11736 & a8398;
assign a11740 = a11738 & ~a6248;
assign a11742 = a11740 & ~a8282;
assign a11744 = a11742 & ~a8112;
assign a11746 = a11744 & ~a7942;
assign a11748 = a11746 & ~a7772;
assign a11750 = a11748 & ~a7602;
assign a11752 = a11750 & ~a7432;
assign a11754 = a11752 & ~a7262;
assign a11756 = a11754 & ~a7092;
assign a11758 = a11756 & ~a6922;
assign a11760 = a11758 & ~a6752;
assign a11762 = a11760 & ~a6582;
assign a11764 = a11762 & ~a6412;
assign a11766 = a11764 & ~a6242;
assign a11768 = a11766 & ~a6174;
assign a11770 = a11768 & ~a6170;
assign a11772 = a11770 & ~a6168;
assign a11774 = a11772 & ~a6164;
assign a11776 = a11774 & ~a6162;
assign a11778 = a11776 & ~a6160;
assign a11780 = a11778 & ~a6158;
assign a11782 = a11780 & ~a6154;
assign a11784 = a11782 & ~a6152;
assign a11786 = a11784 & ~a6148;
assign a11788 = a11786 & ~a6146;
assign a11790 = a11788 & ~a6144;
assign a11792 = a11790 & ~a6142;
assign a11794 = a11792 & ~a6138;
assign a11796 = a11794 & ~a6136;
assign a11798 = a11796 & ~a6132;
assign a11800 = a11798 & ~a6130;
assign a11802 = a11800 & ~a6128;
assign a11804 = a11802 & ~a6126;
assign a11806 = a11804 & ~a6122;
assign a11808 = a11806 & ~a6120;
assign a11810 = a11808 & ~a6116;
assign a11812 = a11810 & ~a6114;
assign a11814 = a11812 & ~a6112;
assign a11816 = a11814 & ~a6110;
assign a11818 = a11816 & ~a6108;
assign a11820 = a11818 & ~a6106;
assign a11822 = a11820 & ~a6104;
assign a11824 = a11822 & ~a6102;
assign a11826 = a11824 & ~a6100;
assign a11828 = a11826 & ~a6098;
assign a11830 = a11828 & ~a6096;
assign a11832 = a11830 & ~a6094;
assign a11834 = a11832 & ~a6092;
assign a11836 = a11834 & ~a6090;
assign a11838 = a11836 & ~a6088;
assign a11840 = a11838 & ~a6086;
assign a11842 = a11840 & ~a6084;
assign a11844 = a11842 & ~a6082;
assign a11846 = a11844 & ~a6080;
assign a11848 = a11846 & ~a6078;
assign a11850 = a11848 & ~a6076;
assign a11852 = a11850 & ~a6074;
assign a11854 = a11852 & ~a6072;
assign a11856 = a11854 & ~a6070;
assign a11858 = a11856 & ~a6068;
assign a11860 = a11858 & ~a6066;
assign a11862 = a11860 & ~a6064;
assign a11864 = a11862 & ~a6062;
assign a11866 = a11864 & ~a6060;
assign a11868 = a11866 & ~a6058;
assign a11870 = a11868 & ~a6056;
assign a11872 = a11870 & ~a6054;
assign a11874 = a11872 & ~a6052;
assign a11876 = a11874 & ~a6050;
assign a11878 = a11876 & ~a6048;
assign a11880 = a11878 & ~a6046;
assign a11882 = a11880 & ~a6044;
assign a11884 = a11882 & ~a6042;
assign a11886 = a11884 & ~a6040;
assign a11888 = a11886 & ~a6038;
assign a11890 = a11888 & ~a6036;
assign a11892 = a11890 & ~a6032;
assign a11894 = a11892 & ~a6030;
assign a11896 = a11894 & ~a6026;
assign a11898 = a11896 & ~a6024;
assign a11900 = a11898 & ~a6020;
assign a11902 = a11900 & ~a6018;
assign a11904 = a11902 & ~a6014;
assign a11906 = a11904 & ~a6012;
assign a11908 = a11906 & ~a6008;
assign a11910 = a11908 & ~a6006;
assign a11912 = a11910 & ~a6002;
assign a11914 = a11912 & ~a6000;
assign a11916 = a11914 & ~a5996;
assign a11918 = a11916 & ~a5994;
assign a11920 = a11918 & ~a5990;
assign a11922 = a11920 & ~a5988;
assign a11924 = a11922 & ~a5984;
assign a11926 = a11924 & ~a5982;
assign a11928 = a11926 & ~a5978;
assign a11930 = a11928 & ~a5976;
assign a11932 = a11930 & ~a5972;
assign a11934 = a11932 & ~a5970;
assign a11936 = a11934 & l1094;
assign a11938 = a11936 & a5966;
assign a11942 = a11936 & i466;
assign p0 = a11942;

assert property (~p0);

endmodule
