module ms177 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26;

output p0;

wire a394,a410,a418,a430,a440,a456,a506,a518,a526,a530,na536,na572,a576,a584,a590,
a594,a602,a610,a622,z0,z1,a630,c1,a650,a652,na648,a656,a664,a670,a674,
a682,a700,a708,na714,a730,a744,a754,na760,na778,na786,na794,na802,na810,nl188,a822,
a834,na840,nl126,na860,na880,a886,na892,na898,a928,na934,na944,na952,na960,na968,na990,
na998,na1006,na1014,na1022,na1030,na1038,na1046,na1054,na1062,na1068,na1074,na1080,na1086,na1094,na1104,
na1108,a1112,z2,nl194,na1118,na1128,na1134,a1142,z3,a1150,na1158,na1170,na1178,na1186,a1192,
a1200,a1210,a1254,na1258,z4,a1268,a1292,a1320,na356,na1322,c0,z5,z6,z7,z8,
a570,a1328,a1336,na1342,a1350,na1356,z9,a1362,a1368,na1376,na1388,na1396,na1404,z10,na1410,
z11,a1444,a1454,a1464,na1470,a1474,na1480,a1504,a1530,a1538,z12,na1544,na1546,a634,na466,
z13,na1552,na1558,a1560,a1562,z14,na1576,na1584,na1592,na1600,na1608,a348,a350,a352,a354,
a356,a358,a360,a362,a364,a366,a368,a370,a372,a374,a376,a378,a380,a382,a384,
a386,a388,a390,a392,a396,a398,a400,a402,a404,a406,a408,a412,a414,a416,a420,
a422,a424,a426,a428,a432,a434,a436,a438,a442,a444,a446,a448,a450,a452,a454,
a458,a460,a462,a464,a466,a468,a470,a472,a474,a476,a478,a480,a482,a484,a486,
a488,a490,a492,a494,a496,a498,a500,a502,a504,a508,a510,a512,a514,a516,a520,
a522,a524,a528,a532,a534,a536,a538,a540,a542,a544,a546,a548,a550,a552,a554,
a556,a558,a560,a562,a564,a566,a568,a572,a574,a578,a580,a582,a586,a588,a592,
a596,a598,a600,a604,a606,a608,a612,a614,a616,a618,a620,a624,a626,a628,a632,
a636,a638,a640,a642,a644,a646,a648,a654,a658,a660,a662,a666,a668,a672,a676,
a678,a680,a684,a686,a688,a690,a692,a694,a696,a698,a702,a704,a706,a710,a712,
a714,a716,a718,a720,a722,a724,a726,a728,a732,a734,a736,a738,a740,a742,a746,
a748,a750,a752,a756,a758,a760,a762,a764,a766,a768,a770,a772,a774,a776,a778,
a780,a782,a784,a786,a788,a790,a792,a794,a796,a798,a800,a802,a804,a806,a808,
a810,a812,a814,a816,a818,a820,a824,a826,a828,a830,a832,a836,a838,a840,a842,
a844,a846,a848,a850,a852,a854,a856,a858,a860,a862,a864,a866,a868,a870,a872,
a874,a876,a878,a880,a882,a884,a888,a890,a892,a894,a896,a898,a900,a902,a904,
a906,a908,a910,a912,a914,a916,a918,a920,a922,a924,a926,a930,a932,a934,a936,
a938,a940,a942,a944,a946,a948,a950,a952,a954,a956,a958,a960,a962,a964,a966,
a968,a970,a972,a974,a976,a978,a980,a982,a984,a986,a988,a990,a992,a994,a996,
a998,a1000,a1002,a1004,a1006,a1008,a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,
a1028,a1030,a1032,a1034,a1036,a1038,a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,
a1058,a1060,a1062,a1064,a1066,a1068,a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,
a1088,a1090,a1092,a1094,a1096,a1098,a1100,a1102,a1104,a1106,a1108,a1110,a1114,a1116,a1118,
a1120,a1122,a1124,a1126,a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1144,a1146,a1148,a1152,
a1154,a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,a1178,a1180,a1182,
a1184,a1186,a1188,a1190,a1194,a1196,a1198,a1202,a1204,a1206,a1208,a1212,a1214,a1216,a1218,
a1220,a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,a1248,
a1250,a1252,a1256,a1258,a1260,a1262,a1264,a1266,a1270,a1272,a1274,a1276,a1278,a1280,a1282,
a1284,a1286,a1288,a1290,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,a1310,a1312,a1314,
a1316,a1318,a1322,a1324,a1326,a1330,a1332,a1334,a1338,a1340,a1342,a1344,a1346,a1348,a1352,
a1354,a1356,a1358,a1360,a1364,a1366,a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,
a1388,a1390,a1392,a1394,a1396,a1398,a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,
a1418,a1420,a1422,a1424,a1426,a1428,a1430,a1432,a1434,a1436,a1438,a1440,a1442,a1446,a1448,
a1450,a1452,a1456,a1458,a1460,a1462,a1466,a1468,a1470,a1472,a1476,a1478,a1480,a1482,a1484,
a1486,a1488,a1490,a1492,a1494,a1496,a1498,a1500,a1502,a1506,a1508,a1510,a1512,a1514,a1516,
a1518,a1520,a1522,a1524,a1526,a1528,a1532,a1534,a1536,a1540,a1542,a1544,a1546,a1548,a1550,
a1552,a1554,a1556,a1558,a1564,a1566,a1568,a1570,a1572,a1574,a1576,a1578,a1580,a1582,a1584,
a1586,a1588,a1590,a1592,a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,a1610,a1612,a1614,
a1616,a1618,a1620,p0;

reg l28,l30,l32,l34,l36,l38,l40,l42,l44,l46,l48,l50,l52,l54,l56,
l58,l60,l62,l64,l66,l68,l70,l72,l74,l76,l78,l80,l82,l84,l86,
l88,l90,l92,l94,l96,l98,l100,l102,l104,l106,l108,l110,l112,l114,l116,
l118,l120,l122,l124,l126,l128,l130,l132,l134,l136,l138,l140,l142,l144,l146,
l148,l150,l152,l154,l156,l158,l160,l162,l164,l166,l168,l170,l172,l174,l176,
l178,l180,l182,l184,l186,l188,l190,l192,l194,l196,l198,l200,l202,l204,l206,
l208,l210,l212,l214,l216,l218,l220,l222,l224,l226,l228,l230,l232,l234,l236,
l238,l240,l242,l244,l246,l248,l250,l252,l254,l256,l258,l260,l262,l264,l266,
l268,l270,l272,l274,l276,l278,l280,l282,l284,l286,l288,l290,l292,l294,l296,
l298,l300,l302,l304,l306,l308,l310,l312,l314,l316,l318,l320,l322,l324,l326,
l328,l330,l332,l334,l336,l338,l340,l342,l344,l346;

initial
begin
   l28 = 0;
   l30 = 0;
   l32 = 0;
   l34 = 0;
   l36 = 0;
   l38 = 0;
   l40 = 0;
   l42 = 0;
   l44 = 0;
   l46 = 0;
   l48 = 0;
   l50 = 0;
   l52 = 0;
   l54 = 0;
   l56 = 0;
   l58 = 0;
   l60 = 0;
   l62 = 0;
   l64 = 0;
   l66 = 0;
   l68 = 0;
   l70 = 0;
   l72 = 0;
   l74 = 0;
   l76 = 0;
   l78 = 0;
   l80 = 0;
   l82 = 0;
   l84 = 0;
   l86 = 0;
   l88 = 0;
   l90 = 0;
   l92 = 0;
   l94 = 0;
   l96 = 0;
   l98 = 0;
   l100 = 0;
   l102 = 0;
   l104 = 0;
   l106 = 0;
   l108 = 0;
   l110 = 0;
   l112 = 0;
   l114 = 0;
   l116 = 0;
   l118 = 0;
   l120 = 0;
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
end

always @(posedge a394)
   l28 <= a394;

always @(posedge a410)
   l30 <= a410;

always @(posedge a418)
   l32 <= a418;

always @(posedge a430)
   l34 <= a430;

always @(posedge a440)
   l36 <= a440;

always @(posedge a456)
   l38 <= a456;

always @(posedge l66)
   l40 <= l66;

always @(posedge a506)
   l42 <= a506;

always @(posedge a518)
   l44 <= a518;

always @(posedge a526)
   l46 <= a526;

always @(posedge l96)
   l48 <= l96;

always @(posedge a530)
   l50 <= a530;

always @(posedge na536)
   l52 <= na536;

always @(posedge na572)
   l54 <= na572;

always @(posedge a576)
   l56 <= a576;

always @(posedge a584)
   l58 <= a584;

always @(posedge a590)
   l60 <= a590;

always @(posedge a594)
   l62 <= a594;

always @(posedge a602)
   l64 <= a602;

always @(posedge a610)
   l66 <= a610;

always @(posedge a622)
   l68 <= a622;

always @(posedge z0)
   l70 <= z0;

always @(posedge z1)
   l72 <= z1;

always @(posedge a630)
   l74 <= a630;

always @(posedge c1)
   l76 <= c1;

always @(posedge a650)
   l78 <= a650;

always @(posedge a652)
   l80 <= a652;

always @(posedge na648)
   l82 <= na648;

always @(posedge a656)
   l84 <= a656;

always @(posedge a664)
   l86 <= a664;

always @(posedge a670)
   l88 <= a670;

always @(posedge a674)
   l90 <= a674;

always @(posedge a682)
   l92 <= a682;

always @(posedge a700)
   l94 <= a700;

always @(posedge a708)
   l96 <= a708;

always @(posedge na714)
   l98 <= na714;

always @(posedge a730)
   l100 <= a730;

always @(posedge a744)
   l102 <= a744;

always @(posedge a754)
   l104 <= a754;

always @(posedge l196)
   l106 <= l196;

always @(posedge na760)
   l108 <= na760;

always @(posedge na778)
   l110 <= na778;

always @(posedge na786)
   l112 <= na786;

always @(posedge na794)
   l114 <= na794;

always @(posedge na802)
   l116 <= na802;

always @(posedge na810)
   l118 <= na810;

always @(posedge nl188)
   l120 <= nl188;

always @(posedge a822)
   l122 <= a822;

always @(posedge a834)
   l124 <= a834;

always @(posedge na840)
   l126 <= na840;

always @(posedge nl126)
   l128 <= nl126;

always @(posedge na860)
   l130 <= na860;

always @(posedge na880)
   l132 <= na880;

always @(posedge a886)
   l134 <= a886;

always @(posedge na892)
   l136 <= na892;

always @(posedge na898)
   l138 <= na898;

always @(posedge a928)
   l140 <= a928;

always @(posedge na934)
   l142 <= na934;

always @(posedge na944)
   l144 <= na944;

always @(posedge na952)
   l146 <= na952;

always @(posedge na960)
   l148 <= na960;

always @(posedge na968)
   l150 <= na968;

always @(posedge na990)
   l152 <= na990;

always @(posedge na998)
   l154 <= na998;

always @(posedge na1006)
   l156 <= na1006;

always @(posedge na1014)
   l158 <= na1014;

always @(posedge na1022)
   l160 <= na1022;

always @(posedge na1030)
   l162 <= na1030;

always @(posedge na1038)
   l164 <= na1038;

always @(posedge na1046)
   l166 <= na1046;

always @(posedge na1054)
   l168 <= na1054;

always @(posedge na1062)
   l170 <= na1062;

always @(posedge na1068)
   l172 <= na1068;

always @(posedge na1074)
   l174 <= na1074;

always @(posedge na1080)
   l176 <= na1080;

always @(posedge na1086)
   l178 <= na1086;

always @(posedge na1094)
   l180 <= na1094;

always @(posedge na1104)
   l182 <= na1104;

always @(posedge na1108)
   l184 <= na1108;

always @(posedge a1112)
   l186 <= a1112;

always @(posedge l190)
   l188 <= l190;

always @(posedge l192)
   l190 <= l192;

always @(posedge z2)
   l192 <= z2;

always @(posedge nl194)
   l194 <= nl194;

always @(posedge na1118)
   l196 <= na1118;

always @(posedge na1128)
   l198 <= na1128;

always @(posedge na1134)
   l200 <= na1134;

always @(posedge a1142)
   l202 <= a1142;

always @(posedge z3)
   l204 <= z3;

always @(posedge a1150)
   l206 <= a1150;

always @(posedge na1158)
   l208 <= na1158;

always @(posedge na1170)
   l210 <= na1170;

always @(posedge na1178)
   l212 <= na1178;

always @(posedge na1186)
   l214 <= na1186;

always @(posedge a1192)
   l216 <= a1192;

always @(posedge a1200)
   l218 <= a1200;

always @(posedge l222)
   l220 <= l222;

always @(posedge l224)
   l222 <= l224;

always @(posedge a1210)
   l224 <= a1210;

always @(posedge a1254)
   l226 <= a1254;

always @(posedge na1258)
   l228 <= na1258;

always @(posedge l232)
   l230 <= l232;

always @(posedge z4)
   l232 <= z4;

always @(posedge a1268)
   l234 <= a1268;

always @(posedge a1292)
   l236 <= a1292;

always @(posedge a1320)
   l238 <= a1320;

always @(posedge na356)
   l240 <= na356;

always @(posedge l252)
   l242 <= l252;

always @(posedge na1322)
   l244 <= na1322;

always @(posedge c0)
   l246 <= c0;

always @(posedge z5)
   l248 <= z5;

always @(posedge z6)
   l250 <= z6;

always @(posedge z7)
   l252 <= z7;

always @(posedge z8)
   l254 <= z8;

always @(posedge a570)
   l256 <= a570;

always @(posedge l286)
   l258 <= l286;

always @(posedge a1328)
   l260 <= a1328;

always @(posedge a1336)
   l262 <= a1336;

always @(posedge na1342)
   l264 <= na1342;

always @(posedge a1350)
   l266 <= a1350;

always @(posedge na1356)
   l268 <= na1356;

always @(posedge z9)
   l270 <= z9;

always @(posedge a1362)
   l272 <= a1362;

always @(posedge a1368)
   l274 <= a1368;

always @(posedge na1376)
   l276 <= na1376;

always @(posedge na1388)
   l278 <= na1388;

always @(posedge na1396)
   l280 <= na1396;

always @(posedge na1404)
   l282 <= na1404;

always @(posedge z10)
   l284 <= z10;

always @(posedge na1410)
   l286 <= na1410;

always @(posedge l290)
   l288 <= l290;

always @(posedge z11)
   l290 <= z11;

always @(posedge a1444)
   l292 <= a1444;

always @(posedge a1454)
   l294 <= a1454;

always @(posedge a1464)
   l296 <= a1464;

always @(posedge na1470)
   l298 <= na1470;

always @(posedge a1474)
   l300 <= a1474;

always @(posedge na1480)
   l302 <= na1480;

always @(posedge a1504)
   l304 <= a1504;

always @(posedge a1530)
   l306 <= a1530;

always @(posedge a1538)
   l308 <= a1538;

always @(posedge z12)
   l310 <= z12;

always @(posedge na1544)
   l312 <= na1544;

always @(posedge na1546)
   l314 <= na1546;

always @(posedge a634)
   l316 <= a634;

always @(posedge i22)
   l318 <= i22;

always @(posedge na466)
   l320 <= na466;

always @(posedge z13)
   l322 <= z13;

always @(posedge na1552)
   l324 <= na1552;

always @(posedge i26)
   l326 <= i26;

always @(posedge na1558)
   l328 <= na1558;

always @(posedge i24)
   l330 <= i24;

always @(posedge a1560)
   l332 <= a1560;

always @(posedge a1562)
   l334 <= a1562;

always @(posedge z14)
   l336 <= z14;

always @(posedge na1576)
   l338 <= na1576;

always @(posedge na1584)
   l340 <= na1584;

always @(posedge na1592)
   l342 <= na1592;

always @(posedge na1600)
   l344 <= na1600;

always @(posedge na1608)
   l346 <= na1608;


assign a394 = ~a392 & a356;
assign a410 = ~a408 & ~a396;
assign a418 = ~a416 & ~a414;
assign a430 = ~a428 & ~a422;
assign a440 = ~a438 & ~a436;
assign a456 = ~a454 & ~a450;
assign a506 = ~a504 & a466;
assign a518 = ~a516 & ~a508;
assign a526 = a524 & a520;
assign a530 = ~a528 & l28;
assign na536 = ~a536;
assign na572 = ~a572;
assign a576 = ~a574 & a572;
assign a584 = ~a582 & a578;
assign a590 = ~a588 & a578;
assign a594 = ~a592 & a572;
assign a602 = a600 & a572;
assign a610 = ~a608 & ~l334;
assign a622 = ~a620 & ~a618;
assign z0 = l42;
assign z1 = l28;
assign a630 = ~a628 & ~l80;
assign c1 = 1;
assign a650 = ~a648 & ~l82;
assign a652 = ~l70 & ~l42;
assign na648 = ~a648;
assign a656 = ~a654 & a648;
assign a664 = ~a662 & a658;
assign a670 = ~a668 & a658;
assign a674 = ~a672 & a648;
assign a682 = a680 & a648;
assign a700 = ~a698 & l42;
assign a708 = a706 & l122;
assign na714 = ~a714;
assign a730 = ~a728 & ~a724;
assign a744 = ~a742 & ~a734;
assign a754 = ~a752 & ~a750;
assign na760 = ~a760;
assign na778 = ~a778;
assign na786 = ~a786;
assign na794 = ~a794;
assign na802 = ~a802;
assign na810 = ~a810;
assign nl188 = ~l188;
assign a822 = ~a820 & ~a708;
assign a834 = ~a832 & ~a830;
assign na840 = ~a840;
assign nl126 = ~l126;
assign na860 = ~a860;
assign na880 = ~a880;
assign a886 = ~a884 & ~a882;
assign na892 = ~a892;
assign na898 = ~a898;
assign a928 = ~a926 & l142;
assign na934 = ~a934;
assign na944 = ~a944;
assign na952 = ~a952;
assign na960 = ~a960;
assign na968 = ~a968;
assign na990 = ~a990;
assign na998 = ~a998;
assign na1006 = ~a1006;
assign na1014 = ~a1014;
assign na1022 = ~a1022;
assign na1030 = ~a1030;
assign na1038 = ~a1038;
assign na1046 = ~a1046;
assign na1054 = ~a1054;
assign na1062 = ~a1062;
assign na1068 = ~a1068;
assign na1074 = ~a1074;
assign na1080 = ~a1080;
assign na1086 = ~a1086;
assign na1094 = ~a1094;
assign na1104 = ~a1104;
assign na1108 = ~a1108;
assign a1112 = ~a1110 & ~l54;
assign z2 = l120;
assign nl194 = ~l194;
assign na1118 = ~a1118;
assign na1128 = ~a1128;
assign na1134 = ~a1134;
assign a1142 = a1140 & a1136;
assign z3 = l74;
assign a1150 = ~a1148 & ~a1142;
assign na1158 = ~a1158;
assign na1170 = ~a1170;
assign na1178 = ~a1178;
assign na1186 = ~a1186;
assign a1192 = ~a1190 & ~l318;
assign a1200 = a1198 & ~a1196;
assign a1210 = a1208 & ~a1204;
assign a1254 = ~a1252 & ~a1214;
assign na1258 = ~a1258;
assign z4 = l218;
assign a1268 = a1266 & ~a1260;
assign a1292 = a1290 & ~a1286;
assign a1320 = a1318 & ~a1314;
assign na356 = ~a356;
assign na1322 = ~a1322;
assign c0 = 0;
assign z5 = c0;
assign z6 = c0;
assign z7 = c0;
assign z8 = l40;
assign a570 = a566 & i6;
assign a1328 = ~a1326 & ~a1324;
assign a1336 = ~a1334 & a1330;
assign na1342 = ~a1342;
assign a1350 = ~a1348 & a1330;
assign na1356 = ~a1356;
assign z9 = l258;
assign a1362 = ~a1360 & ~a1358;
assign a1368 = ~a1366 & ~a526;
assign na1376 = ~a1376;
assign na1388 = ~a1388;
assign na1396 = ~a1396;
assign na1404 = ~a1404;
assign z10 = c0;
assign na1410 = ~a1410;
assign z11 = l76;
assign a1444 = ~a1442 & ~a1414;
assign a1454 = a1452 & ~a1446;
assign a1464 = ~a1462 & a1456;
assign na1470 = ~a1470;
assign a1474 = ~a1472 & a1456;
assign na1480 = ~a1480;
assign a1504 = a1502 & ~a1498;
assign a1530 = a1528 & ~a1524;
assign a1538 = ~a1536 & ~a1534;
assign z12 = l204;
assign na1544 = ~a1544;
assign na1546 = ~a1546;
assign a634 = a632 & i10;
assign na466 = ~a466;
assign z13 = l68;
assign na1552 = ~a1552;
assign na1558 = ~a1558;
assign a1560 = ~a572 & ~l54;
assign a1562 = ~l72 & ~l28;
assign z14 = l32;
assign na1576 = ~a1576;
assign na1584 = ~a1584;
assign na1592 = ~a1592;
assign na1600 = ~a1600;
assign na1608 = ~a1608;
assign a348 = ~l36 & ~l34;
assign a350 = l40 & ~l38;
assign a352 = ~a350 & ~a348;
assign a354 = l46 & l30;
assign a356 = ~a354 & ~a352;
assign a358 = l52 & l32;
assign a360 = ~l44 & l42;
assign a362 = ~a360 & ~l50;
assign a364 = a362 & a358;
assign a366 = l54 & ~l28;
assign a368 = a366 & ~l38;
assign a370 = ~a360 & l34;
assign a372 = ~a370 & ~a368;
assign a374 = a372 & ~a364;
assign a376 = l108 & ~l28;
assign a378 = ~l340 & ~l338;
assign a380 = l344 & ~l342;
assign a382 = l346 & l34;
assign a384 = a382 & a380;
assign a386 = a384 & a378;
assign a388 = ~a386 & ~a376;
assign a390 = a388 & a374;
assign a392 = a390 & ~l28;
assign a396 = ~a356 & l30;
assign a398 = l50 & l32;
assign a400 = a398 & l48;
assign a402 = l50 & l36;
assign a404 = a402 & ~a360;
assign a406 = ~a404 & ~a400;
assign a408 = a406 & ~l30;
assign a412 = a406 & a374;
assign a414 = ~a412 & l32;
assign a416 = a388 & ~l32;
assign a420 = a390 & a356;
assign a422 = ~a420 & l34;
assign a424 = a360 & l36;
assign a426 = a424 & ~a352;
assign a428 = ~a426 & ~l34;
assign a432 = a406 & a356;
assign a434 = a432 & ~a426;
assign a436 = ~a434 & l36;
assign a438 = a374 & ~l36;
assign a442 = ~l236 & ~l234;
assign a444 = ~l238 & ~l228;
assign a446 = a444 & ~l28;
assign a448 = a446 & ~l240;
assign a450 = a448 & a442;
assign a452 = ~l38 & ~l30;
assign a454 = a452 & ~l108;
assign a458 = l202 & l44;
assign a460 = ~l104 & ~l102;
assign a462 = l204 & ~l100;
assign a464 = ~a462 & ~a460;
assign a466 = ~a464 & ~a458;
assign a468 = ~l30 & l28;
assign a470 = l98 & l68;
assign a472 = a470 & ~a468;
assign a474 = ~a472 & ~l96;
assign a476 = ~a474 & ~l94;
assign a478 = l82 & ~l42;
assign a480 = a478 & ~l100;
assign a482 = ~a468 & l102;
assign a484 = ~a482 & ~a480;
assign a486 = a484 & ~a476;
assign a488 = l108 & ~l42;
assign a490 = ~l110 & l102;
assign a492 = l114 & ~l112;
assign a494 = l118 & ~l116;
assign a496 = a494 & a492;
assign a498 = a496 & a490;
assign a500 = ~a498 & ~a488;
assign a502 = a500 & a486;
assign a504 = a502 & ~l42;
assign a508 = ~a466 & l44;
assign a510 = ~a468 & l104;
assign a512 = ~a510 & ~l96;
assign a514 = ~a512 & l94;
assign a516 = ~a514 & ~l44;
assign a520 = l276 & l274;
assign a522 = ~l280 & l278;
assign a524 = a522 & l282;
assign a528 = ~l108 & ~l50;
assign a532 = l336 & ~l120;
assign a534 = l120 & l52;
assign a536 = ~a534 & ~a532;
assign a538 = l64 & l62;
assign a540 = a538 & ~l60;
assign a542 = a540 & ~l58;
assign a544 = a542 & l56;
assign a546 = a544 & i2;
assign a548 = l70 & ~l42;
assign a550 = ~a548 & ~l68;
assign a552 = l72 & ~l28;
assign a554 = ~a552 & ~l32;
assign a556 = ~a554 & ~a550;
assign a558 = l74 & l66;
assign a560 = a558 & i4;
assign a562 = a560 & a556;
assign a564 = ~a562 & l76;
assign a566 = a564 & ~l66;
assign a568 = a566 & a546;
assign a572 = ~a570 & ~a568;
assign a574 = ~a542 & ~l56;
assign a578 = a572 & ~a544;
assign a580 = ~a540 & l58;
assign a582 = ~a580 & ~a542;
assign a586 = ~a538 & l60;
assign a588 = ~a586 & ~a540;
assign a592 = ~a544 & l62;
assign a596 = ~a544 & a538;
assign a598 = ~a592 & ~l64;
assign a600 = ~a598 & ~a596;
assign a604 = l28 & i14;
assign a606 = ~l332 & ~l66;
assign a608 = a606 & ~a604;
assign a612 = a470 & l106;
assign a614 = ~a612 & ~a514;
assign a616 = a614 & a486;
assign a618 = ~a616 & l68;
assign a620 = a500 & ~l68;
assign a624 = l42 & i8;
assign a626 = ~l78 & ~l74;
assign a628 = a626 & ~a624;
assign a632 = a564 & ~l74;
assign a636 = l92 & l90;
assign a638 = a636 & ~l88;
assign a640 = a638 & ~l86;
assign a642 = a640 & l84;
assign a644 = a642 & i12;
assign a646 = a644 & a632;
assign a648 = ~a646 & ~a634;
assign a654 = ~a640 & ~l84;
assign a658 = a648 & ~a642;
assign a660 = ~a638 & l86;
assign a662 = ~a660 & ~a640;
assign a666 = ~a636 & l88;
assign a668 = ~a666 & ~a638;
assign a672 = ~a642 & l90;
assign a676 = ~a642 & a636;
assign a678 = ~a672 & ~l92;
assign a680 = ~a678 & ~a676;
assign a684 = l326 & l324;
assign a686 = l330 & l328;
assign a688 = ~a686 & ~a684;
assign a690 = l186 & l180;
assign a692 = ~a690 & l308;
assign a694 = a692 & ~a688;
assign a696 = ~l108 & ~l94;
assign a698 = a696 & ~a694;
assign a702 = ~l112 & l110;
assign a704 = a494 & ~l114;
assign a706 = a704 & a702;
assign a710 = l322 & ~l120;
assign a712 = l120 & l98;
assign a714 = ~a712 & ~a710;
assign a716 = ~l304 & ~l216;
assign a718 = a716 & ~l306;
assign a720 = ~l294 & ~l42;
assign a722 = a720 & ~l320;
assign a724 = a722 & a718;
assign a726 = ~l108 & ~l100;
assign a728 = a726 & ~l44;
assign a732 = a502 & a466;
assign a734 = ~a732 & l102;
assign a736 = ~l200 & l104;
assign a738 = a736 & a468;
assign a740 = a738 & ~a464;
assign a742 = ~a740 & ~l102;
assign a746 = ~a740 & a466;
assign a748 = a746 & ~a514;
assign a750 = ~a748 & l104;
assign a752 = a486 & ~l104;
assign a756 = a562 & ~l194;
assign a758 = l194 & l108;
assign a760 = ~a758 & ~a756;
assign a762 = ~l124 & ~l122;
assign a764 = ~l126 & l102;
assign a766 = ~a764 & a762;
assign a768 = ~l114 & l112;
assign a770 = ~a768 & ~a492;
assign a772 = a770 & ~a766;
assign a774 = ~a772 & ~l120;
assign a776 = l120 & l110;
assign a778 = ~a776 & ~a774;
assign a780 = ~a766 & ~l118;
assign a782 = ~a780 & ~l120;
assign a784 = l120 & l112;
assign a786 = ~a784 & ~a782;
assign a788 = ~a766 & ~l110;
assign a790 = ~a788 & ~l120;
assign a792 = l120 & l114;
assign a794 = ~a792 & ~a790;
assign a796 = ~a766 & ~l114;
assign a798 = ~a796 & ~l120;
assign a800 = l120 & l116;
assign a802 = ~a800 & ~a798;
assign a804 = ~a766 & ~l116;
assign a806 = ~a804 & ~l120;
assign a808 = l120 & l118;
assign a810 = ~a808 & ~a806;
assign a812 = ~l132 & ~l130;
assign a814 = a812 & l124;
assign a816 = l136 & l134;
assign a818 = ~a816 & ~a814;
assign a820 = a818 & ~l122;
assign a824 = ~a812 & l124;
assign a826 = a824 & a706;
assign a828 = ~a826 & a818;
assign a830 = ~a828 & l124;
assign a832 = ~a612 & ~l124;
assign a836 = l128 & ~l120;
assign a838 = l126 & l120;
assign a840 = ~a838 & ~a836;
assign a842 = ~l178 & ~l176;
assign a844 = ~l182 & ~l180;
assign a846 = ~a844 & ~l120;
assign a848 = a846 & ~a842;
assign a850 = l182 & ~l180;
assign a852 = l178 & ~l176;
assign a854 = ~a852 & ~a850;
assign a856 = a854 & a848;
assign a858 = l130 & l120;
assign a860 = ~a858 & ~a856;
assign a862 = ~l180 & ~l132;
assign a864 = a862 & ~l176;
assign a866 = ~l178 & l176;
assign a868 = ~l182 & l180;
assign a870 = ~a868 & ~a866;
assign a872 = a870 & ~a864;
assign a874 = ~a872 & a854;
assign a876 = ~a874 & a848;
assign a878 = l132 & l120;
assign a880 = ~a878 & ~a876;
assign a882 = ~a818 & l134;
assign a884 = ~a826 & ~l134;
assign a888 = l138 & ~l120;
assign a890 = l136 & l120;
assign a892 = ~a890 & ~a888;
assign a894 = l140 & ~l120;
assign a896 = l138 & l120;
assign a898 = ~a896 & ~a894;
assign a900 = l146 & ~l144;
assign a902 = l150 & l148;
assign a904 = l154 & l152;
assign a906 = a904 & a902;
assign a908 = a906 & a900;
assign a910 = l158 & l156;
assign a912 = l162 & l160;
assign a914 = a912 & a910;
assign a916 = l166 & l164;
assign a918 = l170 & l168;
assign a920 = a918 & a916;
assign a922 = a920 & a914;
assign a924 = a922 & a908;
assign a926 = ~a924 & ~l140;
assign a930 = l174 & ~l120;
assign a932 = l142 & l120;
assign a934 = ~a932 & ~a930;
assign a936 = ~a924 & l142;
assign a938 = ~a936 & l144;
assign a940 = a936 & l164;
assign a942 = ~a940 & l172;
assign a944 = a942 & ~a938;
assign a946 = ~a936 & l146;
assign a948 = a936 & l148;
assign a950 = ~a948 & l172;
assign a952 = a950 & ~a946;
assign a954 = ~a936 & l148;
assign a956 = a936 & l150;
assign a958 = ~a956 & l172;
assign a960 = a958 & ~a954;
assign a962 = ~a936 & l150;
assign a964 = a936 & l154;
assign a966 = ~a964 & l172;
assign a968 = a966 & ~a962;
assign a970 = ~a936 & l152;
assign a972 = ~l146 & l144;
assign a974 = ~a972 & ~a900;
assign a976 = ~l150 & ~l148;
assign a978 = ~a976 & ~a902;
assign a980 = a978 & a974;
assign a982 = ~a978 & ~a974;
assign a984 = ~a982 & ~a980;
assign a986 = ~a984 & a936;
assign a988 = ~a986 & l172;
assign a990 = a988 & ~a970;
assign a992 = ~a936 & l154;
assign a994 = a936 & l152;
assign a996 = ~a994 & l172;
assign a998 = a996 & ~a992;
assign a1000 = ~a936 & l156;
assign a1002 = a936 & l146;
assign a1004 = ~a1002 & l172;
assign a1006 = a1004 & ~a1000;
assign a1008 = ~a936 & l158;
assign a1010 = a936 & l168;
assign a1012 = ~a1010 & l172;
assign a1014 = a1012 & ~a1008;
assign a1016 = ~a936 & l160;
assign a1018 = a936 & l156;
assign a1020 = ~a1018 & l172;
assign a1022 = a1020 & ~a1016;
assign a1024 = ~a936 & l162;
assign a1026 = a936 & l166;
assign a1028 = ~a1026 & l172;
assign a1030 = a1028 & ~a1024;
assign a1032 = ~a936 & l164;
assign a1034 = a936 & l158;
assign a1036 = ~a1034 & l172;
assign a1038 = a1036 & ~a1032;
assign a1040 = ~a936 & l166;
assign a1042 = a936 & l160;
assign a1044 = ~a1042 & l172;
assign a1046 = a1044 & ~a1040;
assign a1048 = ~a936 & l168;
assign a1050 = a936 & l170;
assign a1052 = ~a1050 & l172;
assign a1054 = a1052 & ~a1048;
assign a1056 = ~a936 & l170;
assign a1058 = a936 & l162;
assign a1060 = ~a1058 & l172;
assign a1062 = a1060 & ~a1056;
assign a1064 = l142 & ~l120;
assign a1066 = l172 & l120;
assign a1068 = ~a1066 & ~a1064;
assign a1070 = l134 & ~l120;
assign a1072 = l174 & l120;
assign a1074 = ~a1072 & ~a1070;
assign a1076 = l186 & ~l120;
assign a1078 = l176 & l120;
assign a1080 = ~a1078 & ~a1076;
assign a1082 = l184 & ~l120;
assign a1084 = l178 & l120;
assign a1086 = ~a1084 & ~a1082;
assign a1088 = l82 & i16;
assign a1090 = ~l180 & ~l108;
assign a1092 = ~a1090 & ~l82;
assign a1094 = ~a1092 & ~a1088;
assign a1096 = ~i18 & i16;
assign a1098 = ~a1096 & l82;
assign a1100 = l182 & ~l82;
assign a1102 = a1100 & ~l108;
assign a1104 = ~a1102 & ~a1098;
assign a1106 = l184 & ~l108;
assign a1108 = ~a1106 & ~l54;
assign a1110 = ~l186 & ~l108;
assign a1114 = l198 & ~l120;
assign a1116 = l196 & l120;
assign a1118 = ~a1116 & ~a1114;
assign a1120 = l94 & l68;
assign a1122 = ~a1120 & ~l200;
assign a1124 = ~a1122 & ~l194;
assign a1126 = l198 & l194;
assign a1128 = ~a1126 & ~a1124;
assign a1130 = a398 & ~l194;
assign a1132 = l200 & l194;
assign a1134 = ~a1132 & ~a1130;
assign a1136 = l208 & l206;
assign a1138 = ~l212 & l210;
assign a1140 = a1138 & l214;
assign a1144 = l220 & l218;
assign a1146 = a1144 & ~l216;
assign a1148 = ~a1146 & ~l206;
assign a1152 = ~l210 & l206;
assign a1154 = ~a1152 & ~l120;
assign a1156 = l208 & l120;
assign a1158 = ~a1156 & ~a1154;
assign a1160 = l212 & ~l210;
assign a1162 = ~a1138 & l206;
assign a1164 = a1162 & ~a1160;
assign a1166 = ~a1164 & ~l120;
assign a1168 = l210 & l120;
assign a1170 = ~a1168 & ~a1166;
assign a1172 = ~l214 & l206;
assign a1174 = ~a1172 & ~l120;
assign a1176 = l212 & l120;
assign a1178 = ~a1176 & ~a1174;
assign a1180 = ~l208 & l206;
assign a1182 = ~a1180 & ~l120;
assign a1184 = l214 & l120;
assign a1186 = ~a1184 & ~a1182;
assign a1188 = a724 & l100;
assign a1190 = ~a1188 & ~l216;
assign a1194 = l292 & l204;
assign a1196 = ~a1194 & ~l218;
assign a1198 = ~a1144 & ~l216;
assign a1202 = l226 & l40;
assign a1204 = ~a1202 & ~l224;
assign a1206 = l230 & l224;
assign a1208 = ~a1206 & ~l228;
assign a1212 = ~l228 & ~l40;
assign a1214 = ~a1212 & l226;
assign a1216 = ~l260 & l258;
assign a1218 = ~l264 & l262;
assign a1220 = l264 & ~l262;
assign a1222 = ~a1220 & ~a1218;
assign a1224 = a1222 & ~a1216;
assign a1226 = l268 & ~l266;
assign a1228 = ~l268 & l266;
assign a1230 = ~a1228 & ~l230;
assign a1232 = ~l272 & l270;
assign a1234 = ~a1232 & a1230;
assign a1236 = a1234 & ~a1226;
assign a1238 = a1236 & a1224;
assign a1240 = ~l236 & ~l38;
assign a1242 = a1240 & a444;
assign a1244 = a1242 & ~l242;
assign a1246 = a1244 & ~a1238;
assign a1248 = ~a1246 & ~l30;
assign a1250 = ~a1248 & ~l234;
assign a1252 = ~a1250 & ~l226;
assign a1256 = a450 & l38;
assign a1258 = ~a1256 & ~l228;
assign a1260 = a1248 & ~l234;
assign a1262 = ~l226 & ~l224;
assign a1264 = ~a1262 & l228;
assign a1266 = ~a1264 & ~l46;
assign a1270 = l244 & l226;
assign a1272 = ~l244 & ~l28;
assign a1274 = a1272 & a442;
assign a1276 = ~a1274 & ~a1270;
assign a1278 = ~a1276 & ~l40;
assign a1280 = a1240 & ~l252;
assign a1282 = a1280 & a444;
assign a1284 = a1282 & a1278;
assign a1286 = ~a1284 & ~l236;
assign a1288 = ~l252 & ~l40;
assign a1290 = a1288 & ~l256;
assign a1294 = l244 & ~l242;
assign a1296 = a1294 & a446;
assign a1298 = a1296 & a350;
assign a1300 = ~l250 & ~l248;
assign a1302 = a1300 & ~l246;
assign a1304 = ~a1302 & l244;
assign a1306 = ~a1304 & ~a1298;
assign a1308 = a446 & ~l234;
assign a1310 = a1308 & a1280;
assign a1312 = a1310 & ~a1306;
assign a1314 = ~a1312 & ~l238;
assign a1316 = l254 & ~l40;
assign a1318 = ~a1316 & ~l252;
assign a1322 = ~l244 & ~l108;
assign a1324 = l274 & ~l258;
assign a1326 = ~l274 & ~l260;
assign a1330 = a406 & ~a352;
assign a1332 = l284 & l36;
assign a1334 = ~a1332 & ~l262;
assign a1338 = l274 & l262;
assign a1340 = ~l274 & l264;
assign a1342 = ~a1340 & ~a1338;
assign a1344 = ~l186 & ~l184;
assign a1346 = ~a1344 & a1332;
assign a1348 = ~a1346 & ~l266;
assign a1352 = l274 & l266;
assign a1354 = ~l274 & l268;
assign a1356 = ~a1354 & ~a1352;
assign a1358 = l274 & ~l270;
assign a1360 = ~l274 & ~l272;
assign a1364 = a1206 & ~l228;
assign a1366 = ~a1364 & ~l274;
assign a1370 = ~l278 & l274;
assign a1372 = ~a1370 & ~l120;
assign a1374 = l276 & l120;
assign a1376 = ~a1374 & ~a1372;
assign a1378 = l280 & ~l278;
assign a1380 = ~a522 & l274;
assign a1382 = a1380 & ~a1378;
assign a1384 = ~a1382 & ~l120;
assign a1386 = l278 & l120;
assign a1388 = ~a1386 & ~a1384;
assign a1390 = ~l282 & l274;
assign a1392 = ~a1390 & ~l120;
assign a1394 = l280 & l120;
assign a1396 = ~a1394 & ~a1392;
assign a1398 = ~l276 & l274;
assign a1400 = ~a1398 & ~l120;
assign a1402 = l282 & l120;
assign a1404 = ~a1402 & ~a1400;
assign a1406 = l288 & ~l120;
assign a1408 = l286 & l120;
assign a1410 = ~a1408 & ~a1406;
assign a1412 = ~l216 & ~l204;
assign a1414 = ~a1412 & l292;
assign a1416 = l298 & ~l296;
assign a1418 = ~l298 & l296;
assign a1420 = ~a1418 & ~l220;
assign a1422 = ~l302 & l300;
assign a1424 = l302 & ~l300;
assign a1426 = ~a1424 & ~a1422;
assign a1428 = a1426 & a1420;
assign a1430 = a1428 & ~a1416;
assign a1432 = a718 & ~l100;
assign a1434 = a1432 & ~l242;
assign a1436 = a1434 & ~a1430;
assign a1438 = ~a1436 & ~l44;
assign a1440 = ~a1438 & ~l294;
assign a1442 = ~a1440 & ~l292;
assign a1446 = a1438 & ~l294;
assign a1448 = ~l292 & ~l218;
assign a1450 = ~a1448 & l216;
assign a1452 = ~a1450 & ~l202;
assign a1456 = ~a514 & ~a464;
assign a1458 = l284 & l104;
assign a1460 = a1458 & ~a844;
assign a1462 = ~a1460 & ~l296;
assign a1466 = l296 & l206;
assign a1468 = l298 & ~l206;
assign a1470 = ~a1468 & ~a1466;
assign a1472 = ~a1458 & ~l300;
assign a1476 = l300 & l206;
assign a1478 = l302 & ~l206;
assign a1480 = ~a1478 & ~a1476;
assign a1482 = a1432 & ~l252;
assign a1484 = ~l308 & ~l204;
assign a1486 = a1484 & ~l304;
assign a1488 = a1486 & a720;
assign a1490 = l308 & l292;
assign a1492 = a1490 & ~l204;
assign a1494 = ~a1492 & ~a1488;
assign a1496 = ~a1494 & a1482;
assign a1498 = ~a1496 & ~l304;
assign a1500 = ~l252 & ~l204;
assign a1502 = a1500 & ~l316;
assign a1506 = l308 & ~l216;
assign a1508 = a1506 & ~l306;
assign a1510 = a462 & ~l242;
assign a1512 = a1510 & ~l42;
assign a1514 = a1512 & a1508;
assign a1516 = ~a1302 & l308;
assign a1518 = ~a1516 & ~a1514;
assign a1520 = ~a1518 & a720;
assign a1522 = a1520 & a1482;
assign a1524 = ~a1522 & ~l306;
assign a1526 = l310 & ~l204;
assign a1528 = ~a1526 & ~l252;
assign a1532 = l312 & l308;
assign a1534 = a1532 & ~l314;
assign a1536 = ~l308 & ~l108;
assign a1540 = ~l120 & i20;
assign a1542 = l312 & l120;
assign a1544 = ~a1542 & ~a1540;
assign a1546 = ~l314 & ~l312;
assign a1548 = ~l194 & c0;
assign a1550 = l324 & l194;
assign a1552 = ~a1550 & ~a1548;
assign a1554 = ~l120 & c0;
assign a1556 = l328 & l120;
assign a1558 = ~a1556 & ~a1554;
assign a1564 = ~l344 & l342;
assign a1566 = ~l126 & l34;
assign a1568 = a1566 & ~a380;
assign a1570 = a1568 & ~a1564;
assign a1572 = ~a1570 & ~l120;
assign a1574 = l338 & l120;
assign a1576 = ~a1574 & ~a1572;
assign a1578 = a1566 & ~l344;
assign a1580 = ~a1578 & ~l120;
assign a1582 = l340 & l120;
assign a1584 = ~a1582 & ~a1580;
assign a1586 = a1566 & ~l346;
assign a1588 = ~a1586 & ~l120;
assign a1590 = l342 & l120;
assign a1592 = ~a1590 & ~a1588;
assign a1594 = a1566 & ~l338;
assign a1596 = ~a1594 & ~l120;
assign a1598 = l344 & l120;
assign a1600 = ~a1598 & ~a1596;
assign a1602 = a1566 & ~l340;
assign a1604 = ~a1602 & ~l120;
assign a1606 = l346 & l120;
assign a1608 = ~a1606 & ~a1604;
assign a1610 = a348 & ~l32;
assign a1612 = ~a1610 & ~a468;
assign a1614 = ~a348 & l32;
assign a1616 = l30 & ~l28;
assign a1618 = ~a1616 & ~a1614;
assign a1620 = a1618 & ~a1612;
assign p0 = ~a1620;

assert property (~p0);

endmodule
