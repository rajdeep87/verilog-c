module m6s17 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66;

output p0;

wire na526,na566,na614,na654,na674,na680,na704,a716,a726,na742,na758,a768,na778,na788,c1,
na1014,na1044,na1054,na1080,na1106,na1114,na1158,na1206,na1212,na1214,na1222,na1228,na1234,na1246,na1258,
na1270,na1272,a1502,na1510,na1516,na1522,na1532,na1542,na1552,na1558,na1564,na1570,a1612,a1620,a1626,
na1638,na1644,na1654,na1664,na1674,na1682,na1692,na1702,na1714,na1798,na1870,na1936,na2026,na2092,na2146,
na2194,na2266,na2308,na2314,na2320,na2328,na2336,na2344,na2352,na2360,na2366,na2374,na2382,na2390,na2398,
na2406,a2272,na2416,na2422,na2428,na2434,na2442,na2448,na2456,na2462,na2492,na2498,na2514,na2520,na2532,
na2538,na2546,na2552,na2560,na2566,na2574,na2580,na2588,na2594,na2600,na2606,na2612,na2620,na2626,na2634,
na2640,na2648,na2654,na2660,na2666,na2672,na2678,na2686,na2692,na2698,na2704,na2710,na2718,na2724,na2730,
na2736,na2742,na2750,na2756,na2762,na2768,na2774,na2782,na2788,na2794,na2802,na2808,na2816,na2822,na2828,
na2836,na2842,na2848,na2878,na2884,na2894,na2900,na2908,na2914,na2922,na2928,na2936,na2942,na2950,na2956,
na2964,na2970,na2976,na2982,na2990,na2996,na3004,na3010,na3018,na3024,na3032,na3038,na3044,na3052,na3058,
na3066,na3072,na3078,na3086,na3092,na3100,na3106,na3114,na3120,na3126,na3132,na3140,na3146,na3154,na3160,
na3168,na3174,na3184,na3194,na3204,a438,a440,a442,a444,a446,a448,a450,a452,a454,a456,
a458,a460,a462,a464,a466,a468,a470,a472,a474,a476,a478,a480,a482,a484,a486,
a488,a490,a492,a494,a496,a498,a500,a502,a504,a506,a508,a510,a512,a514,a516,
a518,a520,a522,a524,a526,a528,a530,a532,a534,a536,a538,a540,a542,a544,a546,
a548,a550,a552,a554,a556,a558,a560,a562,a564,a566,a568,a570,a572,a574,a576,
a578,a580,a582,a584,a586,a588,a590,a592,a594,a596,a598,a600,a602,a604,a606,
a608,a610,a612,a614,a616,a618,a620,a622,a624,a626,a628,a630,a632,a634,a636,
a638,a640,a642,a644,a646,a648,a650,a652,a654,a656,a658,a660,a662,a664,a666,
a668,a670,a672,a674,a676,a678,a680,a682,a684,a686,a688,a690,a692,a694,a696,
a698,a700,a702,a704,a706,a708,a710,a712,a714,a718,a720,a722,a724,a728,a730,
a732,a734,a736,a738,a740,a742,a744,a746,a748,a750,a752,a754,a756,a758,a760,
a762,a764,a766,a770,a772,a774,a776,a778,a780,a782,a784,a786,a788,a790,a792,
a794,a796,a798,a800,a802,a804,a806,a808,a810,a812,a814,a816,a818,a820,a822,
a824,a826,a828,a830,a832,a834,a836,a838,a840,a842,a844,a846,a848,a850,a852,
a854,a856,a858,a860,a862,a864,a866,a868,a870,a872,a874,a876,a878,a880,a882,
a884,a886,a888,a890,a892,a894,a896,a898,a900,a902,a904,a906,a908,a910,a912,
a914,a916,a918,a920,a922,a924,a926,a928,a930,a932,a934,a936,a938,a940,a942,
a944,a946,a948,a950,a952,a954,a956,a958,a960,a962,a964,a966,a968,a970,a972,
a974,a976,a978,a980,a982,a984,a986,a988,a990,a992,a994,a996,a998,a1000,a1002,
a1004,a1006,a1008,a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,
a1034,a1036,a1038,a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,a1062,
a1064,a1066,a1068,a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,a1092,
a1094,a1096,a1098,a1100,a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,
a1124,a1126,a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,
a1154,a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,a1178,a1180,a1182,
a1184,a1186,a1188,a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,a1208,a1210,a1212,
a1214,a1216,a1218,a1220,a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1242,
a1244,a1246,a1248,a1250,a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,a1268,a1270,a1272,
a1274,a1276,a1278,a1280,a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,
a1304,a1306,a1308,a1310,a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,
a1334,a1336,a1338,a1340,a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,
a1364,a1366,a1368,a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,a1388,a1390,a1392,
a1394,a1396,a1398,a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,
a1424,a1426,a1428,a1430,a1432,a1434,a1436,a1438,a1440,a1442,a1444,a1446,a1448,a1450,a1452,
a1454,a1456,a1458,a1460,a1462,a1464,a1466,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1482,
a1484,a1486,a1488,a1490,a1492,a1494,a1496,a1498,a1500,a1504,a1506,a1508,a1510,a1512,a1514,
a1516,a1518,a1520,a1522,a1524,a1526,a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,
a1546,a1548,a1550,a1552,a1554,a1556,a1558,a1560,a1562,a1564,a1566,a1568,a1570,a1572,a1574,
a1576,a1578,a1580,a1582,a1584,a1586,a1588,a1590,a1592,a1594,a1596,a1598,a1600,a1602,a1604,
a1606,a1608,a1610,a1614,a1616,a1618,a1622,a1624,a1628,a1630,a1632,a1634,a1636,a1638,a1640,
a1642,a1644,a1646,a1648,a1650,a1652,a1654,a1656,a1658,a1660,a1662,a1664,a1666,a1668,a1670,
a1672,a1674,a1676,a1678,a1680,a1682,a1684,a1686,a1688,a1690,a1692,a1694,a1696,a1698,a1700,
a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,
a1732,a1734,a1736,a1738,a1740,a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,a1758,a1760,
a1762,a1764,a1766,a1768,a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,a1790,
a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,
a1822,a1824,a1826,a1828,a1830,a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,a1848,a1850,
a1852,a1854,a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,
a1882,a1884,a1886,a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,a1910,
a1912,a1914,a1916,a1918,a1920,a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,a1938,a1940,
a1942,a1944,a1946,a1948,a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,
a1972,a1974,a1976,a1978,a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,a1998,a2000,
a2002,a2004,a2006,a2008,a2010,a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,a2030,
a2032,a2034,a2036,a2038,a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,a2058,a2060,
a2062,a2064,a2066,a2068,a2070,a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,a2090,
a2092,a2094,a2096,a2098,a2100,a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,a2120,
a2122,a2124,a2126,a2128,a2130,a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,
a2152,a2154,a2156,a2158,a2160,a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,a2178,a2180,
a2182,a2184,a2186,a2188,a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,a2208,a2210,
a2212,a2214,a2216,a2218,a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,a2238,a2240,
a2242,a2244,a2246,a2248,a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,a2268,a2270,
a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,a2298,a2300,a2302,
a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,a2328,a2330,a2332,
a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,a2358,a2360,a2362,
a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,a2388,a2390,a2392,
a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,a2420,a2422,
a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,a2448,a2450,a2452,
a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,a2478,a2480,a2482,
a2484,a2486,a2488,a2490,a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,a2508,a2510,a2512,
a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,a2540,a2542,
a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,a2572,
a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,a2602,
a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,a2630,a2632,
a2634,a2636,a2638,a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,a2662,
a2664,a2666,a2668,a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,a2692,
a2694,a2696,a2698,a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,a2718,a2720,a2722,
a2724,a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,a2752,
a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,a2782,
a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,a2810,a2812,
a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,a2840,a2842,
a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,a2870,a2872,
a2874,a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,a2900,a2902,
a2904,a2906,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2930,a2932,
a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,a2960,a2962,
a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,a2988,a2990,a2992,
a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,a3022,
a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,a3048,a3050,a3052,
a3054,a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,a3078,a3080,a3082,
a3084,a3086,a3088,a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,a3112,
a3114,a3116,a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,a3142,
a3144,a3146,a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,a3172,
a3174,a3176,a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3200,a3202,
a3204,p0;

reg l68,l70,l72,l74,l76,l78,l80,l82,l84,l86,l88,l90,l92,l94,l96,
l98,l100,l102,l104,l106,l108,l110,l112,l114,l116,l118,l120,l122,l124,l126,
l128,l130,l132,l134,l136,l138,l140,l142,l144,l146,l148,l150,l152,l154,l156,
l158,l160,l162,l164,l166,l168,l170,l172,l174,l176,l178,l180,l182,l184,l186,
l188,l190,l192,l194,l196,l198,l200,l202,l204,l206,l208,l210,l212,l214,l216,
l218,l220,l222,l224,l226,l228,l230,l232,l234,l236,l238,l240,l242,l244,l246,
l248,l250,l252,l254,l256,l258,l260,l262,l264,l266,l268,l270,l272,l274,l276,
l278,l280,l282,l284,l286,l288,l290,l292,l294,l296,l298,l300,l302,l304,l306,
l308,l310,l312,l314,l316,l318,l320,l322,l324,l326,l328,l330,l332,l334,l336,
l338,l340,l342,l344,l346,l348,l350,l352,l354,l356,l358,l360,l362,l364,l366,
l368,l370,l372,l374,l376,l378,l380,l382,l384,l386,l388,l390,l392,l394,l396,
l398,l400,l402,l404,l406,l408,l410,l412,l414,l416,l418,l420,l422,l424,l426,
l428,l430,l432,l434,l436;

initial
begin
   l68 = 0;
   l70 = 0;
   l72 = 0;
   l74 = 0;
   l76 = 0;
   l78 = 0;
   l80 = 0;
   l82 = 0;
   l84 = 0;
   l86 = 0;
   l88 = 0;
   l90 = 0;
   l92 = 0;
   l94 = 0;
   l96 = 0;
   l98 = 0;
   l100 = 0;
   l102 = 0;
   l104 = 0;
   l106 = 0;
   l108 = 0;
   l110 = 0;
   l112 = 0;
   l114 = 0;
   l116 = 0;
   l118 = 0;
   l120 = 0;
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
   l392 = 0;
   l394 = 0;
   l396 = 0;
   l398 = 0;
   l400 = 0;
   l402 = 0;
   l404 = 0;
   l406 = 0;
   l408 = 0;
   l410 = 0;
   l412 = 0;
   l414 = 0;
   l416 = 0;
   l418 = 0;
   l420 = 0;
   l422 = 0;
   l424 = 0;
   l426 = 0;
   l428 = 0;
   l430 = 0;
   l432 = 0;
   l434 = 0;
   l436 = 0;
end

always @(posedge na526)
   l68 <= na526;

always @(posedge na566)
   l70 <= na566;

always @(posedge na614)
   l72 <= na614;

always @(posedge na654)
   l74 <= na654;

always @(posedge na674)
   l76 <= na674;

always @(posedge na680)
   l78 <= na680;

always @(posedge na704)
   l80 <= na704;

always @(posedge a716)
   l82 <= a716;

always @(posedge a726)
   l84 <= a726;

always @(posedge na742)
   l86 <= na742;

always @(posedge na758)
   l88 <= na758;

always @(posedge a768)
   l90 <= a768;

always @(posedge na778)
   l92 <= na778;

always @(posedge na788)
   l94 <= na788;

always @(posedge c1)
   l96 <= c1;

always @(posedge na1014)
   l98 <= na1014;

always @(posedge na1044)
   l100 <= na1044;

always @(posedge na1054)
   l102 <= na1054;

always @(posedge na1080)
   l104 <= na1080;

always @(posedge na1106)
   l106 <= na1106;

always @(posedge na1114)
   l108 <= na1114;

always @(posedge na1158)
   l110 <= na1158;

always @(posedge na1206)
   l112 <= na1206;

always @(posedge na1212)
   l114 <= na1212;

always @(posedge na1214)
   l116 <= na1214;

always @(posedge na1222)
   l118 <= na1222;

always @(posedge na1228)
   l120 <= na1228;

always @(posedge na1234)
   l122 <= na1234;

always @(posedge na1246)
   l124 <= na1246;

always @(posedge na1258)
   l126 <= na1258;

always @(posedge na1270)
   l128 <= na1270;

always @(posedge na1272)
   l130 <= na1272;

always @(posedge a1502)
   l132 <= a1502;

always @(posedge na1510)
   l134 <= na1510;

always @(posedge na1516)
   l136 <= na1516;

always @(posedge na1522)
   l138 <= na1522;

always @(posedge na1532)
   l140 <= na1532;

always @(posedge na1542)
   l142 <= na1542;

always @(posedge na1552)
   l144 <= na1552;

always @(posedge na1558)
   l146 <= na1558;

always @(posedge na1564)
   l148 <= na1564;

always @(posedge na1570)
   l150 <= na1570;

always @(posedge a1612)
   l152 <= a1612;

always @(posedge a1620)
   l154 <= a1620;

always @(posedge a1626)
   l156 <= a1626;

always @(posedge na1638)
   l158 <= na1638;

always @(posedge na1644)
   l160 <= na1644;

always @(posedge na1654)
   l162 <= na1654;

always @(posedge na1664)
   l164 <= na1664;

always @(posedge na1674)
   l166 <= na1674;

always @(posedge na1682)
   l168 <= na1682;

always @(posedge na1692)
   l170 <= na1692;

always @(posedge na1702)
   l172 <= na1702;

always @(posedge na1714)
   l174 <= na1714;

always @(posedge na1798)
   l176 <= na1798;

always @(posedge na1870)
   l178 <= na1870;

always @(posedge na1936)
   l180 <= na1936;

always @(posedge na2026)
   l182 <= na2026;

always @(posedge na2092)
   l184 <= na2092;

always @(posedge na2146)
   l186 <= na2146;

always @(posedge na2194)
   l188 <= na2194;

always @(posedge na2266)
   l190 <= na2266;

always @(posedge na2308)
   l192 <= na2308;

always @(posedge na2314)
   l194 <= na2314;

always @(posedge na2320)
   l196 <= na2320;

always @(posedge na2328)
   l198 <= na2328;

always @(posedge na2336)
   l200 <= na2336;

always @(posedge na2344)
   l202 <= na2344;

always @(posedge na2352)
   l204 <= na2352;

always @(posedge na2360)
   l206 <= na2360;

always @(posedge na2366)
   l208 <= na2366;

always @(posedge na2374)
   l210 <= na2374;

always @(posedge na2382)
   l212 <= na2382;

always @(posedge na2390)
   l214 <= na2390;

always @(posedge na2398)
   l216 <= na2398;

always @(posedge na2406)
   l218 <= na2406;

always @(posedge a2272)
   l220 <= a2272;

always @(posedge na2416)
   l222 <= na2416;

always @(posedge na2422)
   l224 <= na2422;

always @(posedge na2428)
   l226 <= na2428;

always @(posedge na2434)
   l228 <= na2434;

always @(posedge na2442)
   l230 <= na2442;

always @(posedge na2448)
   l232 <= na2448;

always @(posedge na2456)
   l234 <= na2456;

always @(posedge na2462)
   l236 <= na2462;

always @(posedge na2492)
   l238 <= na2492;

always @(posedge na2498)
   l240 <= na2498;

always @(posedge na2514)
   l242 <= na2514;

always @(posedge na2520)
   l244 <= na2520;

always @(posedge na2532)
   l246 <= na2532;

always @(posedge na2538)
   l248 <= na2538;

always @(posedge na2546)
   l250 <= na2546;

always @(posedge na2552)
   l252 <= na2552;

always @(posedge na2560)
   l254 <= na2560;

always @(posedge na2566)
   l256 <= na2566;

always @(posedge na2574)
   l258 <= na2574;

always @(posedge na2580)
   l260 <= na2580;

always @(posedge na2588)
   l262 <= na2588;

always @(posedge na2594)
   l264 <= na2594;

always @(posedge na2600)
   l266 <= na2600;

always @(posedge na2606)
   l268 <= na2606;

always @(posedge na2612)
   l270 <= na2612;

always @(posedge na2620)
   l272 <= na2620;

always @(posedge na2626)
   l274 <= na2626;

always @(posedge na2634)
   l276 <= na2634;

always @(posedge na2640)
   l278 <= na2640;

always @(posedge na2648)
   l280 <= na2648;

always @(posedge na2654)
   l282 <= na2654;

always @(posedge na2660)
   l284 <= na2660;

always @(posedge na2666)
   l286 <= na2666;

always @(posedge na2672)
   l288 <= na2672;

always @(posedge na2678)
   l290 <= na2678;

always @(posedge na2686)
   l292 <= na2686;

always @(posedge na2692)
   l294 <= na2692;

always @(posedge na2698)
   l296 <= na2698;

always @(posedge na2704)
   l298 <= na2704;

always @(posedge na2710)
   l300 <= na2710;

always @(posedge na2718)
   l302 <= na2718;

always @(posedge na2724)
   l304 <= na2724;

always @(posedge na2730)
   l306 <= na2730;

always @(posedge na2736)
   l308 <= na2736;

always @(posedge na2742)
   l310 <= na2742;

always @(posedge na2750)
   l312 <= na2750;

always @(posedge na2756)
   l314 <= na2756;

always @(posedge na2762)
   l316 <= na2762;

always @(posedge na2768)
   l318 <= na2768;

always @(posedge na2774)
   l320 <= na2774;

always @(posedge na2782)
   l322 <= na2782;

always @(posedge na2788)
   l324 <= na2788;

always @(posedge na2794)
   l326 <= na2794;

always @(posedge na2802)
   l328 <= na2802;

always @(posedge na2808)
   l330 <= na2808;

always @(posedge na2816)
   l332 <= na2816;

always @(posedge na2822)
   l334 <= na2822;

always @(posedge na2828)
   l336 <= na2828;

always @(posedge na2836)
   l338 <= na2836;

always @(posedge na2842)
   l340 <= na2842;

always @(posedge na2848)
   l342 <= na2848;

always @(posedge na2878)
   l344 <= na2878;

always @(posedge na2884)
   l346 <= na2884;

always @(posedge na2894)
   l348 <= na2894;

always @(posedge na2900)
   l350 <= na2900;

always @(posedge na2908)
   l352 <= na2908;

always @(posedge na2914)
   l354 <= na2914;

always @(posedge na2922)
   l356 <= na2922;

always @(posedge na2928)
   l358 <= na2928;

always @(posedge na2936)
   l360 <= na2936;

always @(posedge na2942)
   l362 <= na2942;

always @(posedge na2950)
   l364 <= na2950;

always @(posedge na2956)
   l366 <= na2956;

always @(posedge na2964)
   l368 <= na2964;

always @(posedge na2970)
   l370 <= na2970;

always @(posedge na2976)
   l372 <= na2976;

always @(posedge na2982)
   l374 <= na2982;

always @(posedge na2990)
   l376 <= na2990;

always @(posedge na2996)
   l378 <= na2996;

always @(posedge na3004)
   l380 <= na3004;

always @(posedge na3010)
   l382 <= na3010;

always @(posedge na3018)
   l384 <= na3018;

always @(posedge na3024)
   l386 <= na3024;

always @(posedge na3032)
   l388 <= na3032;

always @(posedge na3038)
   l390 <= na3038;

always @(posedge na3044)
   l392 <= na3044;

always @(posedge na3052)
   l394 <= na3052;

always @(posedge na3058)
   l396 <= na3058;

always @(posedge na3066)
   l398 <= na3066;

always @(posedge na3072)
   l400 <= na3072;

always @(posedge na3078)
   l402 <= na3078;

always @(posedge na3086)
   l404 <= na3086;

always @(posedge na3092)
   l406 <= na3092;

always @(posedge na3100)
   l408 <= na3100;

always @(posedge na3106)
   l410 <= na3106;

always @(posedge na3114)
   l412 <= na3114;

always @(posedge na3120)
   l414 <= na3120;

always @(posedge na3126)
   l416 <= na3126;

always @(posedge na3132)
   l418 <= na3132;

always @(posedge na3140)
   l420 <= na3140;

always @(posedge na3146)
   l422 <= na3146;

always @(posedge na3154)
   l424 <= na3154;

always @(posedge na3160)
   l426 <= na3160;

always @(posedge na3168)
   l428 <= na3168;

always @(posedge na3174)
   l430 <= na3174;

always @(posedge na3184)
   l432 <= na3184;

always @(posedge na3194)
   l434 <= na3194;

always @(posedge na3204)
   l436 <= na3204;


assign na526 = ~a526;
assign na566 = ~a566;
assign na614 = ~a614;
assign na654 = ~a654;
assign na674 = ~a674;
assign na680 = ~a680;
assign na704 = ~a704;
assign a716 = ~a714 & ~a712;
assign a726 = ~a724 & ~a722;
assign na742 = ~a742;
assign na758 = ~a758;
assign a768 = a766 & ~a508;
assign na778 = ~a778;
assign na788 = ~a788;
assign c1 = 1;
assign na1014 = ~a1014;
assign na1044 = ~a1044;
assign na1054 = ~a1054;
assign na1080 = ~a1080;
assign na1106 = ~a1106;
assign na1114 = ~a1114;
assign na1158 = ~a1158;
assign na1206 = ~a1206;
assign na1212 = ~a1212;
assign na1214 = ~a1214;
assign na1222 = ~a1222;
assign na1228 = ~a1228;
assign na1234 = ~a1234;
assign na1246 = ~a1246;
assign na1258 = ~a1258;
assign na1270 = ~a1270;
assign na1272 = ~a1272;
assign a1502 = ~a1500 & ~a1442;
assign na1510 = ~a1510;
assign na1516 = ~a1516;
assign na1522 = ~a1522;
assign na1532 = ~a1532;
assign na1542 = ~a1542;
assign na1552 = ~a1552;
assign na1558 = ~a1558;
assign na1564 = ~a1564;
assign na1570 = ~a1570;
assign a1612 = ~a1610 & ~a1608;
assign a1620 = ~a1618 & ~a1616;
assign a1626 = ~a1624 & ~a1606;
assign na1638 = ~a1638;
assign na1644 = ~a1644;
assign na1654 = ~a1654;
assign na1664 = ~a1664;
assign na1674 = ~a1674;
assign na1682 = ~a1682;
assign na1692 = ~a1692;
assign na1702 = ~a1702;
assign na1714 = ~a1714;
assign na1798 = ~a1798;
assign na1870 = ~a1870;
assign na1936 = ~a1936;
assign na2026 = ~a2026;
assign na2092 = ~a2092;
assign na2146 = ~a2146;
assign na2194 = ~a2194;
assign na2266 = ~a2266;
assign na2308 = ~a2308;
assign na2314 = ~a2314;
assign na2320 = ~a2320;
assign na2328 = ~a2328;
assign na2336 = ~a2336;
assign na2344 = ~a2344;
assign na2352 = ~a2352;
assign na2360 = ~a2360;
assign na2366 = ~a2366;
assign na2374 = ~a2374;
assign na2382 = ~a2382;
assign na2390 = ~a2390;
assign na2398 = ~a2398;
assign na2406 = ~a2406;
assign a2272 = a2270 & i18;
assign na2416 = ~a2416;
assign na2422 = ~a2422;
assign na2428 = ~a2428;
assign na2434 = ~a2434;
assign na2442 = ~a2442;
assign na2448 = ~a2448;
assign na2456 = ~a2456;
assign na2462 = ~a2462;
assign na2492 = ~a2492;
assign na2498 = ~a2498;
assign na2514 = ~a2514;
assign na2520 = ~a2520;
assign na2532 = ~a2532;
assign na2538 = ~a2538;
assign na2546 = ~a2546;
assign na2552 = ~a2552;
assign na2560 = ~a2560;
assign na2566 = ~a2566;
assign na2574 = ~a2574;
assign na2580 = ~a2580;
assign na2588 = ~a2588;
assign na2594 = ~a2594;
assign na2600 = ~a2600;
assign na2606 = ~a2606;
assign na2612 = ~a2612;
assign na2620 = ~a2620;
assign na2626 = ~a2626;
assign na2634 = ~a2634;
assign na2640 = ~a2640;
assign na2648 = ~a2648;
assign na2654 = ~a2654;
assign na2660 = ~a2660;
assign na2666 = ~a2666;
assign na2672 = ~a2672;
assign na2678 = ~a2678;
assign na2686 = ~a2686;
assign na2692 = ~a2692;
assign na2698 = ~a2698;
assign na2704 = ~a2704;
assign na2710 = ~a2710;
assign na2718 = ~a2718;
assign na2724 = ~a2724;
assign na2730 = ~a2730;
assign na2736 = ~a2736;
assign na2742 = ~a2742;
assign na2750 = ~a2750;
assign na2756 = ~a2756;
assign na2762 = ~a2762;
assign na2768 = ~a2768;
assign na2774 = ~a2774;
assign na2782 = ~a2782;
assign na2788 = ~a2788;
assign na2794 = ~a2794;
assign na2802 = ~a2802;
assign na2808 = ~a2808;
assign na2816 = ~a2816;
assign na2822 = ~a2822;
assign na2828 = ~a2828;
assign na2836 = ~a2836;
assign na2842 = ~a2842;
assign na2848 = ~a2848;
assign na2878 = ~a2878;
assign na2884 = ~a2884;
assign na2894 = ~a2894;
assign na2900 = ~a2900;
assign na2908 = ~a2908;
assign na2914 = ~a2914;
assign na2922 = ~a2922;
assign na2928 = ~a2928;
assign na2936 = ~a2936;
assign na2942 = ~a2942;
assign na2950 = ~a2950;
assign na2956 = ~a2956;
assign na2964 = ~a2964;
assign na2970 = ~a2970;
assign na2976 = ~a2976;
assign na2982 = ~a2982;
assign na2990 = ~a2990;
assign na2996 = ~a2996;
assign na3004 = ~a3004;
assign na3010 = ~a3010;
assign na3018 = ~a3018;
assign na3024 = ~a3024;
assign na3032 = ~a3032;
assign na3038 = ~a3038;
assign na3044 = ~a3044;
assign na3052 = ~a3052;
assign na3058 = ~a3058;
assign na3066 = ~a3066;
assign na3072 = ~a3072;
assign na3078 = ~a3078;
assign na3086 = ~a3086;
assign na3092 = ~a3092;
assign na3100 = ~a3100;
assign na3106 = ~a3106;
assign na3114 = ~a3114;
assign na3120 = ~a3120;
assign na3126 = ~a3126;
assign na3132 = ~a3132;
assign na3140 = ~a3140;
assign na3146 = ~a3146;
assign na3154 = ~a3154;
assign na3160 = ~a3160;
assign na3168 = ~a3168;
assign na3174 = ~a3174;
assign na3184 = ~a3184;
assign na3194 = ~a3194;
assign na3204 = ~a3204;
assign a438 = l68 & i2;
assign a440 = l70 & i4;
assign a442 = ~a440 & ~a438;
assign a444 = l72 & i6;
assign a446 = l74 & i8;
assign a448 = ~a446 & ~a444;
assign a450 = a448 & a442;
assign a452 = ~l78 & ~l76;
assign a454 = a452 & ~a450;
assign a456 = ~l82 & ~l80;
assign a458 = ~l90 & ~l88;
assign a460 = ~l94 & ~l92;
assign a462 = a460 & a458;
assign a464 = a462 & ~l86;
assign a466 = a464 & ~l84;
assign a468 = a466 & a456;
assign a470 = a468 & a454;
assign a472 = l68 & ~i2;
assign a474 = l102 & l100;
assign a476 = a474 & ~l98;
assign a478 = l108 & l106;
assign a480 = a478 & ~l104;
assign a482 = ~a472 & ~l126;
assign a484 = a482 & ~a480;
assign a486 = a484 & a476;
assign a488 = a482 & a480;
assign a490 = ~a472 & l126;
assign a492 = ~a490 & ~a488;
assign a494 = a492 & ~a486;
assign a496 = a484 & ~a476;
assign a498 = l116 & l114;
assign a500 = a498 & ~l112;
assign a502 = ~a456 & l84;
assign a504 = l96 & i10;
assign a506 = a504 & a464;
assign a508 = a506 & ~a502;
assign a510 = ~i14 & i12;
assign a512 = a510 & a508;
assign a514 = l122 & l120;
assign a516 = a514 & ~l118;
assign a518 = ~a516 & ~a512;
assign a520 = a518 & ~a500;
assign a522 = ~a520 & a496;
assign a524 = ~a522 & a494;
assign a526 = a524 & ~a472;
assign a528 = l70 & ~i4;
assign a530 = a474 & l98;
assign a532 = a478 & l104;
assign a534 = ~a528 & ~l128;
assign a536 = a534 & ~a532;
assign a538 = a536 & a530;
assign a540 = a534 & a532;
assign a542 = ~a528 & l128;
assign a544 = ~a542 & ~a540;
assign a546 = a544 & ~a538;
assign a548 = a536 & ~a530;
assign a550 = a498 & l112;
assign a552 = i14 & i12;
assign a554 = a552 & a508;
assign a556 = a514 & l118;
assign a558 = ~a556 & ~a554;
assign a560 = a558 & ~a550;
assign a562 = ~a560 & a548;
assign a564 = ~a562 & a546;
assign a566 = a564 & ~a528;
assign a568 = l72 & ~i6;
assign a570 = l102 & ~l100;
assign a572 = a570 & ~l98;
assign a574 = l108 & ~l106;
assign a576 = a574 & ~l104;
assign a578 = ~a568 & ~l124;
assign a580 = a578 & ~a576;
assign a582 = a580 & a572;
assign a584 = a578 & a576;
assign a586 = ~a568 & l124;
assign a588 = ~a586 & ~a584;
assign a590 = a588 & ~a582;
assign a592 = a580 & ~a572;
assign a594 = l116 & ~l114;
assign a596 = a594 & ~l112;
assign a598 = l122 & ~l120;
assign a600 = a598 & ~l118;
assign a602 = ~i14 & ~i12;
assign a604 = a602 & a508;
assign a606 = ~a604 & ~a600;
assign a608 = a606 & ~a596;
assign a610 = ~a608 & a592;
assign a612 = ~a610 & a590;
assign a614 = a612 & ~a568;
assign a616 = l74 & ~i8;
assign a618 = a570 & l98;
assign a620 = a574 & l104;
assign a622 = ~a616 & ~l110;
assign a624 = a622 & ~a620;
assign a626 = a624 & a618;
assign a628 = a622 & a620;
assign a630 = ~a616 & l110;
assign a632 = ~a630 & ~a628;
assign a634 = a632 & ~a626;
assign a636 = a624 & ~a618;
assign a638 = a594 & l112;
assign a640 = i14 & ~i12;
assign a642 = a640 & a508;
assign a644 = a598 & l118;
assign a646 = ~a644 & ~a642;
assign a648 = a646 & ~a638;
assign a650 = ~a648 & a636;
assign a652 = ~a650 & a634;
assign a654 = a652 & ~a616;
assign a656 = ~a508 & ~a450;
assign a658 = l78 & l76;
assign a660 = ~a658 & ~a452;
assign a662 = ~a660 & a656;
assign a664 = a508 & a450;
assign a666 = a664 & a660;
assign a668 = ~a664 & ~a656;
assign a670 = a668 & l76;
assign a672 = ~a670 & ~a666;
assign a674 = a672 & ~a662;
assign a676 = a668 & l78;
assign a678 = ~a668 & ~l78;
assign a680 = ~a678 & ~a676;
assign a682 = a452 & ~l82;
assign a684 = a682 & ~l80;
assign a686 = ~a682 & l80;
assign a688 = ~a686 & ~a684;
assign a690 = ~a688 & a656;
assign a692 = a664 & a658;
assign a694 = a692 & l82;
assign a696 = a694 & l80;
assign a698 = ~a696 & ~a656;
assign a700 = ~a694 & ~l80;
assign a702 = ~a700 & a698;
assign a704 = ~a702 & ~a690;
assign a706 = a656 & ~a452;
assign a708 = ~a692 & ~a656;
assign a710 = ~a708 & ~a706;
assign a712 = a710 & l82;
assign a714 = ~a710 & ~l82;
assign a718 = ~a684 & a656;
assign a720 = ~a718 & ~a698;
assign a722 = a720 & l84;
assign a724 = ~a720 & ~l84;
assign a728 = ~a508 & a450;
assign a730 = a728 & l86;
assign a732 = a684 & ~l84;
assign a734 = a732 & ~l86;
assign a736 = ~a732 & l86;
assign a738 = ~a736 & ~a734;
assign a740 = ~a738 & a656;
assign a742 = ~a740 & ~a730;
assign a744 = a728 & l88;
assign a746 = a734 & ~l92;
assign a748 = a746 & ~l94;
assign a750 = a748 & ~l88;
assign a752 = ~a748 & l88;
assign a754 = ~a752 & ~a750;
assign a756 = ~a754 & a656;
assign a758 = ~a756 & ~a744;
assign a760 = a750 & ~a450;
assign a762 = a760 & l90;
assign a764 = ~a760 & ~l90;
assign a766 = ~a764 & ~a762;
assign a770 = a728 & l92;
assign a772 = ~a734 & l92;
assign a774 = ~a772 & ~a746;
assign a776 = ~a774 & a656;
assign a778 = ~a776 & ~a770;
assign a780 = a728 & l94;
assign a782 = ~a746 & l94;
assign a784 = ~a782 & ~a748;
assign a786 = ~a784 & a656;
assign a788 = ~a786 & ~a780;
assign a790 = ~a550 & a548;
assign a792 = a790 & a556;
assign a794 = ~a500 & a496;
assign a796 = a794 & a516;
assign a798 = ~a796 & ~a792;
assign a800 = ~a638 & a636;
assign a802 = a800 & a644;
assign a804 = ~a596 & a592;
assign a806 = a804 & a600;
assign a808 = ~a806 & ~a802;
assign a810 = a808 & a798;
assign a812 = a810 & a600;
assign a814 = a550 & a548;
assign a816 = a500 & a496;
assign a818 = ~a816 & ~a814;
assign a820 = a638 & a636;
assign a822 = a596 & a592;
assign a824 = ~a822 & ~a820;
assign a826 = a824 & a818;
assign a828 = a826 & a596;
assign a830 = ~a538 & ~a486;
assign a832 = ~a626 & ~a582;
assign a834 = a832 & a830;
assign a836 = a834 & a572;
assign a838 = ~a540 & ~a488;
assign a840 = ~a628 & ~a584;
assign a842 = a840 & a838;
assign a844 = a842 & a576;
assign a846 = ~a444 & l124;
assign a848 = ~a846 & ~a844;
assign a850 = a848 & ~a836;
assign a852 = a850 & ~a828;
assign a854 = a852 & a812;
assign a856 = ~a854 & a810;
assign a858 = a856 & a644;
assign a860 = a850 & a828;
assign a862 = ~a860 & a826;
assign a864 = a862 & a638;
assign a866 = a848 & a836;
assign a868 = ~a866 & a834;
assign a870 = a868 & a618;
assign a872 = ~a846 & a844;
assign a874 = ~a872 & a842;
assign a876 = a874 & a620;
assign a878 = ~a446 & l110;
assign a880 = ~a878 & ~a876;
assign a882 = a880 & ~a870;
assign a884 = a882 & ~a864;
assign a886 = a884 & a858;
assign a888 = ~a886 & a856;
assign a890 = a888 & a516;
assign a892 = a882 & a864;
assign a894 = ~a892 & a862;
assign a896 = a894 & a500;
assign a898 = a880 & a870;
assign a900 = ~a898 & a868;
assign a902 = a900 & a476;
assign a904 = ~a878 & a876;
assign a906 = ~a904 & a874;
assign a908 = a906 & a480;
assign a910 = ~a438 & l126;
assign a912 = ~a910 & ~a908;
assign a914 = a912 & ~a902;
assign a916 = a914 & ~a896;
assign a918 = a916 & a890;
assign a920 = ~a918 & a888;
assign a922 = a920 & a556;
assign a924 = a914 & a896;
assign a926 = ~a924 & a894;
assign a928 = a926 & a550;
assign a930 = a912 & a902;
assign a932 = ~a930 & a900;
assign a934 = a932 & a530;
assign a936 = ~a910 & a908;
assign a938 = ~a936 & a906;
assign a940 = a938 & a532;
assign a942 = ~a440 & l128;
assign a944 = ~a942 & ~a940;
assign a946 = a944 & ~a934;
assign a948 = a946 & ~a928;
assign a950 = a948 & a922;
assign a952 = ~a950 & a920;
assign a954 = a952 & l122;
assign a956 = a946 & a928;
assign a958 = ~a956 & a926;
assign a960 = a958 & l116;
assign a962 = a960 & a954;
assign a964 = ~a942 & a940;
assign a966 = ~a964 & a938;
assign a968 = a966 & l108;
assign a970 = a944 & a934;
assign a972 = ~a970 & a932;
assign a974 = a972 & l102;
assign a976 = ~a974 & ~a968;
assign a978 = a976 & ~l130;
assign a980 = a978 & a962;
assign a982 = a976 & l130;
assign a984 = ~a982 & ~a980;
assign a986 = a984 & l98;
assign a988 = a980 & l118;
assign a990 = l180 & l178;
assign a992 = a990 & l176;
assign a994 = ~l190 & ~l188;
assign a996 = a994 & l186;
assign a998 = a996 & l184;
assign a1000 = a998 & ~l182;
assign a1002 = a1000 & a992;
assign a1004 = ~a1002 & l436;
assign a1006 = a1002 & ~l436;
assign a1008 = ~a1006 & ~a1004;
assign a1010 = ~a1008 & a982;
assign a1012 = ~a1010 & ~a988;
assign a1014 = a1012 & ~a986;
assign a1016 = a984 & l100;
assign a1018 = a980 & l120;
assign a1020 = ~l180 & l178;
assign a1022 = l190 & l188;
assign a1024 = a1022 & ~l186;
assign a1026 = a1024 & ~l184;
assign a1028 = a1026 & l182;
assign a1030 = a1028 & l176;
assign a1032 = a1030 & a1020;
assign a1034 = ~a1032 & l434;
assign a1036 = a1032 & ~l434;
assign a1038 = ~a1036 & ~a1034;
assign a1040 = ~a1038 & a982;
assign a1042 = ~a1040 & ~a1018;
assign a1044 = a1042 & ~a1016;
assign a1046 = ~a976 & ~a972;
assign a1048 = a978 & ~a962;
assign a1050 = ~a1048 & l102;
assign a1052 = a1050 & ~a1046;
assign a1054 = ~a1052 & a984;
assign a1056 = a984 & l104;
assign a1058 = a980 & l112;
assign a1060 = l180 & ~l178;
assign a1062 = a1024 & l184;
assign a1064 = a1062 & l182;
assign a1066 = a1064 & ~l176;
assign a1068 = a1066 & a1060;
assign a1070 = ~a1068 & l432;
assign a1072 = a1068 & ~l432;
assign a1074 = ~a1072 & ~a1070;
assign a1076 = ~a1074 & a982;
assign a1078 = ~a1076 & ~a1058;
assign a1080 = a1078 & ~a1056;
assign a1082 = a984 & l106;
assign a1084 = a980 & l114;
assign a1086 = l190 & ~l188;
assign a1088 = a1086 & l186;
assign a1090 = a1088 & ~l184;
assign a1092 = a1090 & ~l182;
assign a1094 = a1092 & a992;
assign a1096 = ~a1094 & l174;
assign a1098 = a1094 & ~l174;
assign a1100 = ~a1098 & ~a1096;
assign a1102 = ~a1100 & a982;
assign a1104 = ~a1102 & ~a1084;
assign a1106 = a1104 & ~a1082;
assign a1108 = ~a976 & ~a966;
assign a1110 = ~a1048 & l108;
assign a1112 = a1110 & ~a1108;
assign a1114 = ~a1112 & a984;
assign a1116 = ~a904 & ~a898;
assign a1118 = a1116 & ~a892;
assign a1120 = a804 & ~a600;
assign a1122 = a1120 & a604;
assign a1124 = a800 & ~a644;
assign a1126 = a1124 & a642;
assign a1128 = ~a1126 & ~a1122;
assign a1130 = a794 & ~a516;
assign a1132 = a1130 & a512;
assign a1134 = ~a1132 & a1128;
assign a1136 = a790 & ~a556;
assign a1138 = a1136 & a554;
assign a1140 = ~a1138 & a1134;
assign a1142 = a1140 & a604;
assign a1144 = a852 & ~a812;
assign a1146 = a1144 & a1142;
assign a1148 = ~a1146 & a1140;
assign a1150 = a1148 & a642;
assign a1152 = ~a1150 & ~a858;
assign a1154 = ~a1152 & a884;
assign a1156 = ~a1154 & a1118;
assign a1158 = a1156 & ~a878;
assign a1160 = a884 & ~a858;
assign a1162 = a1160 & a1150;
assign a1164 = ~a1162 & a1148;
assign a1166 = a1164 & a512;
assign a1168 = a916 & ~a890;
assign a1170 = a1168 & a1166;
assign a1172 = ~a1170 & a1164;
assign a1174 = a1172 & a554;
assign a1176 = a948 & ~a922;
assign a1178 = a1176 & a1174;
assign a1180 = ~a1178 & a1172;
assign a1182 = a1180 & a508;
assign a1184 = ~a980 & a954;
assign a1186 = ~a980 & a960;
assign a1188 = a1186 & a1184;
assign a1190 = ~a976 & l130;
assign a1192 = ~a1190 & ~l132;
assign a1194 = a1192 & a1188;
assign a1196 = ~a1194 & a1186;
assign a1198 = a1196 & ~a1184;
assign a1200 = ~a1198 & a1182;
assign a1202 = a1200 & i14;
assign a1204 = ~a1200 & l112;
assign a1206 = ~a1204 & ~a1202;
assign a1208 = a1200 & i12;
assign a1210 = ~a1200 & l114;
assign a1212 = ~a1210 & ~a1208;
assign a1214 = ~a1198 & ~a1182;
assign a1216 = a1198 & a1182;
assign a1218 = a1216 & i14;
assign a1220 = ~a1216 & l118;
assign a1222 = ~a1220 & ~a1218;
assign a1224 = a1216 & i12;
assign a1226 = ~a1216 & l120;
assign a1228 = ~a1226 & ~a1224;
assign a1230 = ~a1194 & a1184;
assign a1232 = a1230 & ~a1186;
assign a1234 = ~a1232 & ~a1216;
assign a1236 = ~a872 & ~a866;
assign a1238 = a1236 & ~a860;
assign a1240 = ~a1142 & ~a812;
assign a1242 = ~a1240 & a852;
assign a1244 = ~a1242 & a1238;
assign a1246 = a1244 & ~a846;
assign a1248 = ~a936 & ~a930;
assign a1250 = a1248 & ~a924;
assign a1252 = ~a1166 & ~a890;
assign a1254 = ~a1252 & a916;
assign a1256 = ~a1254 & a1250;
assign a1258 = a1256 & ~a910;
assign a1260 = ~a970 & ~a964;
assign a1262 = a1260 & ~a956;
assign a1264 = ~a1174 & ~a922;
assign a1266 = ~a1264 & a948;
assign a1268 = ~a1266 & a1262;
assign a1270 = a1268 & ~a942;
assign a1272 = a1192 & ~a1188;
assign a1274 = ~a1190 & l132;
assign a1276 = a1230 & a1196;
assign a1278 = ~l136 & ~l134;
assign a1280 = ~l140 & ~l138;
assign a1282 = a1280 & a1278;
assign a1284 = ~l144 & ~l142;
assign a1286 = l150 & l148;
assign a1288 = a1286 & l146;
assign a1290 = a1288 & a1284;
assign a1292 = a1290 & a1282;
assign a1294 = l136 & l134;
assign a1296 = a1294 & l138;
assign a1298 = a1296 & l140;
assign a1300 = a1298 & l142;
assign a1302 = a1300 & l144;
assign a1304 = a1302 & l146;
assign a1306 = a1304 & l148;
assign a1308 = a1306 & l150;
assign a1310 = ~a1308 & ~a1292;
assign a1312 = l154 & ~l152;
assign a1314 = ~l154 & l152;
assign a1316 = ~a1314 & ~a1312;
assign a1318 = ~a1316 & ~a1310;
assign a1320 = a1316 & a1310;
assign a1322 = ~a1320 & ~a1318;
assign a1324 = ~a1306 & ~l150;
assign a1326 = ~a1324 & ~a1308;
assign a1328 = a1326 & ~a1292;
assign a1330 = a1328 & ~l156;
assign a1332 = ~a1328 & l156;
assign a1334 = ~a1332 & ~a1330;
assign a1336 = ~a1304 & ~l148;
assign a1338 = ~a1336 & ~a1306;
assign a1340 = a1338 & ~a1292;
assign a1342 = a1340 & ~l158;
assign a1344 = ~a1292 & ~l134;
assign a1346 = ~a1344 & l160;
assign a1348 = ~l162 & l144;
assign a1350 = l162 & ~l144;
assign a1352 = ~a1350 & ~a1348;
assign a1354 = ~a1352 & ~a1300;
assign a1356 = ~a1294 & ~l138;
assign a1358 = ~a1356 & ~a1296;
assign a1360 = a1358 & ~l164;
assign a1362 = ~l166 & l142;
assign a1364 = l166 & ~l142;
assign a1366 = ~a1364 & ~a1362;
assign a1368 = a1366 & a1298;
assign a1370 = ~a1368 & ~a1360;
assign a1372 = a1370 & ~a1354;
assign a1374 = a1372 & ~a1346;
assign a1376 = a1352 & a1300;
assign a1378 = ~a1294 & ~a1278;
assign a1380 = a1378 & ~l168;
assign a1382 = ~a1378 & l168;
assign a1384 = ~a1382 & ~a1380;
assign a1386 = ~a1366 & ~a1298;
assign a1388 = ~a1386 & a1384;
assign a1390 = a1388 & ~a1376;
assign a1392 = a1344 & ~l160;
assign a1394 = ~a1358 & l164;
assign a1396 = ~l170 & l140;
assign a1398 = l170 & ~l140;
assign a1400 = ~a1398 & ~a1396;
assign a1402 = a1400 & a1296;
assign a1404 = ~a1400 & ~a1296;
assign a1406 = ~a1404 & ~a1402;
assign a1408 = a1406 & ~a1394;
assign a1410 = a1408 & ~a1392;
assign a1412 = a1410 & a1390;
assign a1414 = a1412 & a1374;
assign a1416 = a1414 & ~a1342;
assign a1418 = ~a1302 & ~l146;
assign a1420 = ~a1418 & ~a1304;
assign a1422 = a1420 & ~a1292;
assign a1424 = a1422 & ~l172;
assign a1426 = ~a1422 & l172;
assign a1428 = ~a1426 & ~a1424;
assign a1430 = ~a1340 & l158;
assign a1432 = ~a1430 & a1428;
assign a1434 = a1432 & a1416;
assign a1436 = a1434 & a1334;
assign a1438 = a1436 & ~a1322;
assign a1440 = ~a1438 & ~a1276;
assign a1442 = ~a1440 & a1274;
assign a1444 = ~l160 & l134;
assign a1446 = l160 & ~l134;
assign a1448 = ~a1446 & ~a1444;
assign a1450 = ~l168 & l136;
assign a1452 = l168 & ~l136;
assign a1454 = ~a1452 & ~a1450;
assign a1456 = a1454 & a1448;
assign a1458 = ~l164 & l138;
assign a1460 = l164 & ~l138;
assign a1462 = ~a1460 & ~a1458;
assign a1464 = a1400 & a1366;
assign a1466 = a1464 & a1462;
assign a1468 = a1466 & a1456;
assign a1470 = ~l172 & l146;
assign a1472 = l172 & ~l146;
assign a1474 = ~a1472 & ~a1470;
assign a1476 = a1474 & a1352;
assign a1478 = ~l158 & l148;
assign a1480 = l158 & ~l148;
assign a1482 = ~a1480 & ~a1478;
assign a1484 = ~l156 & l150;
assign a1486 = l156 & ~l150;
assign a1488 = ~a1486 & ~a1484;
assign a1490 = a1488 & a1316;
assign a1492 = a1490 & a1482;
assign a1494 = a1492 & a1476;
assign a1496 = a1494 & a1468;
assign a1498 = ~a1496 & ~a1276;
assign a1500 = ~a1498 & ~l132;
assign a1504 = ~a1292 & a1274;
assign a1506 = a1504 & ~l134;
assign a1508 = ~a1274 & l134;
assign a1510 = ~a1508 & ~a1506;
assign a1512 = a1504 & a1378;
assign a1514 = ~a1274 & l136;
assign a1516 = ~a1514 & ~a1512;
assign a1518 = a1504 & a1358;
assign a1520 = ~a1274 & l138;
assign a1522 = ~a1520 & ~a1518;
assign a1524 = ~a1296 & ~l140;
assign a1526 = ~a1524 & ~a1298;
assign a1528 = a1526 & a1504;
assign a1530 = ~a1274 & l140;
assign a1532 = ~a1530 & ~a1528;
assign a1534 = ~a1298 & ~l142;
assign a1536 = ~a1534 & ~a1300;
assign a1538 = a1536 & a1504;
assign a1540 = ~a1274 & l142;
assign a1542 = ~a1540 & ~a1538;
assign a1544 = ~a1300 & ~l144;
assign a1546 = ~a1544 & ~a1302;
assign a1548 = a1546 & a1504;
assign a1550 = ~a1274 & l144;
assign a1552 = ~a1550 & ~a1548;
assign a1554 = a1504 & a1420;
assign a1556 = ~a1274 & l146;
assign a1558 = ~a1556 & ~a1554;
assign a1560 = a1504 & a1338;
assign a1562 = ~a1274 & l148;
assign a1564 = ~a1562 & ~a1560;
assign a1566 = a1504 & a1326;
assign a1568 = ~a1274 & l150;
assign a1570 = ~a1568 & ~a1566;
assign a1572 = ~l168 & ~l160;
assign a1574 = ~l170 & ~l164;
assign a1576 = a1574 & a1572;
assign a1578 = ~l166 & ~l162;
assign a1580 = l158 & l156;
assign a1582 = a1580 & l172;
assign a1584 = a1582 & a1578;
assign a1586 = a1584 & a1576;
assign a1588 = l168 & l160;
assign a1590 = a1588 & l164;
assign a1592 = a1590 & l170;
assign a1594 = a1592 & l166;
assign a1596 = a1594 & l162;
assign a1598 = a1596 & l172;
assign a1600 = a1598 & l158;
assign a1602 = a1600 & l156;
assign a1604 = ~a1602 & ~a1586;
assign a1606 = ~a1604 & a1276;
assign a1608 = a1606 & l152;
assign a1610 = ~a1606 & ~l152;
assign a1614 = ~a1310 & a1274;
assign a1616 = a1614 & l154;
assign a1618 = ~a1614 & ~l154;
assign a1622 = a1600 & a1276;
assign a1624 = ~a1622 & ~l156;
assign a1628 = ~a1586 & a1276;
assign a1630 = ~a1598 & ~l158;
assign a1632 = ~a1630 & ~a1600;
assign a1634 = a1632 & a1628;
assign a1636 = ~a1276 & l158;
assign a1638 = ~a1636 & ~a1634;
assign a1640 = a1628 & ~l160;
assign a1642 = ~a1276 & l160;
assign a1644 = ~a1642 & ~a1640;
assign a1646 = ~a1594 & ~l162;
assign a1648 = ~a1646 & ~a1596;
assign a1650 = a1648 & a1628;
assign a1652 = ~a1276 & l162;
assign a1654 = ~a1652 & ~a1650;
assign a1656 = ~a1588 & ~l164;
assign a1658 = ~a1656 & ~a1590;
assign a1660 = a1658 & a1628;
assign a1662 = ~a1276 & l164;
assign a1664 = ~a1662 & ~a1660;
assign a1666 = ~a1592 & ~l166;
assign a1668 = ~a1666 & ~a1594;
assign a1670 = a1668 & a1628;
assign a1672 = ~a1276 & l166;
assign a1674 = ~a1672 & ~a1670;
assign a1676 = ~a1588 & ~a1572;
assign a1678 = a1676 & a1628;
assign a1680 = ~a1276 & l168;
assign a1682 = ~a1680 & ~a1678;
assign a1684 = ~a1590 & ~l170;
assign a1686 = ~a1684 & ~a1592;
assign a1688 = a1686 & a1628;
assign a1690 = ~a1276 & l170;
assign a1692 = ~a1690 & ~a1688;
assign a1694 = ~a1596 & ~l172;
assign a1696 = ~a1694 & ~a1598;
assign a1698 = a1696 & a1628;
assign a1700 = ~a1276 & l172;
assign a1702 = ~a1700 & ~a1698;
assign a1704 = ~a1274 & ~a1194;
assign a1706 = a1704 & l174;
assign a1708 = a1194 & l114;
assign a1710 = a1274 & l272;
assign a1712 = ~a1710 & ~a1708;
assign a1714 = a1712 & ~a1706;
assign a1716 = l306 & l218;
assign a1718 = ~l306 & ~l218;
assign a1720 = ~a1718 & ~a1716;
assign a1722 = l262 & ~l230;
assign a1724 = ~l262 & l230;
assign a1726 = ~a1724 & ~a1722;
assign a1728 = a1726 & a1720;
assign a1730 = ~a1726 & ~a1720;
assign a1732 = ~a1730 & ~a1728;
assign a1734 = l394 & ~l388;
assign a1736 = ~l394 & l388;
assign a1738 = ~a1736 & ~a1734;
assign a1740 = a1738 & l292;
assign a1742 = ~a1738 & ~l292;
assign a1744 = ~a1742 & ~a1740;
assign a1746 = a1744 & ~a1732;
assign a1748 = ~a1744 & a1732;
assign a1750 = ~a1748 & ~a1746;
assign a1752 = ~l328 & l200;
assign a1754 = l328 & ~l200;
assign a1756 = ~a1754 & ~a1752;
assign a1758 = a1756 & l276;
assign a1760 = ~a1756 & ~l276;
assign a1762 = ~a1760 & ~a1758;
assign a1764 = ~l322 & l286;
assign a1766 = l322 & ~l286;
assign a1768 = ~a1766 & ~a1764;
assign a1770 = l424 & ~l316;
assign a1772 = ~l424 & l316;
assign a1774 = ~a1772 & ~a1770;
assign a1776 = a1774 & ~a1768;
assign a1778 = ~a1774 & a1768;
assign a1780 = ~a1778 & ~a1776;
assign a1782 = ~a1780 & a1762;
assign a1784 = a1780 & ~a1762;
assign a1786 = ~a1784 & ~a1782;
assign a1788 = a1786 & ~a1750;
assign a1790 = ~a1786 & a1750;
assign a1792 = ~a1790 & ~a1788;
assign a1794 = a1792 & a1274;
assign a1796 = a1704 & l176;
assign a1798 = ~a1796 & ~a1794;
assign a1800 = ~l292 & l212;
assign a1802 = l292 & ~l212;
assign a1804 = ~a1802 & ~a1800;
assign a1806 = a1804 & l302;
assign a1808 = ~a1804 & ~l302;
assign a1810 = ~a1808 & ~a1806;
assign a1812 = ~l394 & l204;
assign a1814 = l394 & ~l204;
assign a1816 = ~a1814 & ~a1812;
assign a1818 = l312 & ~l258;
assign a1820 = ~l312 & l258;
assign a1822 = ~a1820 & ~a1818;
assign a1824 = a1822 & ~a1816;
assign a1826 = ~a1822 & a1816;
assign a1828 = ~a1826 & ~a1824;
assign a1830 = ~a1828 & a1810;
assign a1832 = a1828 & ~a1810;
assign a1834 = ~a1832 & ~a1830;
assign a1836 = l196 & ~l192;
assign a1838 = ~l196 & l192;
assign a1840 = ~a1838 & ~a1836;
assign a1842 = l428 & ~l230;
assign a1844 = ~l428 & l230;
assign a1846 = ~a1844 & ~a1842;
assign a1848 = a1846 & ~a1840;
assign a1850 = ~a1846 & a1840;
assign a1852 = ~a1850 & ~a1848;
assign a1854 = ~a1852 & a1762;
assign a1856 = a1852 & ~a1762;
assign a1858 = ~a1856 & ~a1854;
assign a1860 = a1858 & ~a1834;
assign a1862 = ~a1858 & a1834;
assign a1864 = ~a1862 & ~a1860;
assign a1866 = a1864 & a1274;
assign a1868 = a1704 & l178;
assign a1870 = ~a1868 & ~a1866;
assign a1872 = l404 & ~l296;
assign a1874 = ~l404 & l296;
assign a1876 = ~a1874 & ~a1872;
assign a1878 = a1876 & l338;
assign a1880 = ~a1876 & ~l338;
assign a1882 = ~a1880 & ~a1878;
assign a1884 = a1882 & ~a1828;
assign a1886 = ~a1882 & a1828;
assign a1888 = ~a1886 & ~a1884;
assign a1890 = ~l388 & l202;
assign a1892 = l388 & ~l202;
assign a1894 = ~a1892 & ~a1890;
assign a1896 = a1894 & l226;
assign a1898 = ~a1894 & ~l226;
assign a1900 = ~a1898 & ~a1896;
assign a1902 = l306 & ~l286;
assign a1904 = ~l306 & l286;
assign a1906 = ~a1904 & ~a1902;
assign a1908 = l420 & ~l280;
assign a1910 = ~l420 & l280;
assign a1912 = ~a1910 & ~a1908;
assign a1914 = a1912 & ~a1906;
assign a1916 = ~a1912 & a1906;
assign a1918 = ~a1916 & ~a1914;
assign a1920 = ~a1918 & a1900;
assign a1922 = a1918 & ~a1900;
assign a1924 = ~a1922 & ~a1920;
assign a1926 = a1924 & ~a1888;
assign a1928 = ~a1924 & a1888;
assign a1930 = ~a1928 & ~a1926;
assign a1932 = a1930 & a1274;
assign a1934 = a1704 & l180;
assign a1936 = ~a1934 & ~a1932;
assign a1938 = ~l404 & l206;
assign a1940 = l404 & ~l206;
assign a1942 = ~a1940 & ~a1938;
assign a1944 = ~l272 & l234;
assign a1946 = l272 & ~l234;
assign a1948 = ~a1946 & ~a1944;
assign a1950 = a1948 & ~a1942;
assign a1952 = ~a1948 & a1942;
assign a1954 = ~a1952 & ~a1950;
assign a1956 = l338 & l208;
assign a1958 = ~l338 & ~l208;
assign a1960 = ~a1958 & ~a1956;
assign a1962 = ~l398 & l328;
assign a1964 = l398 & ~l328;
assign a1966 = ~a1964 & ~a1962;
assign a1968 = a1966 & a1960;
assign a1970 = ~a1966 & ~a1960;
assign a1972 = ~a1970 & ~a1968;
assign a1974 = a1972 & ~a1954;
assign a1976 = ~a1972 & a1954;
assign a1978 = ~a1976 & ~a1974;
assign a1980 = ~l280 & l210;
assign a1982 = l280 & ~l210;
assign a1984 = ~a1982 & ~a1980;
assign a1986 = a1984 & l322;
assign a1988 = ~a1984 & ~l322;
assign a1990 = ~a1988 & ~a1986;
assign a1992 = ~l416 & l262;
assign a1994 = l416 & ~l262;
assign a1996 = ~a1994 & ~a1992;
assign a1998 = l312 & ~l286;
assign a2000 = ~l312 & l286;
assign a2002 = ~a2000 & ~a1998;
assign a2004 = a2002 & ~a1996;
assign a2006 = ~a2002 & a1996;
assign a2008 = ~a2006 & ~a2004;
assign a2010 = ~a2008 & a1990;
assign a2012 = a2008 & ~a1990;
assign a2014 = ~a2012 & ~a2010;
assign a2016 = a2014 & ~a1978;
assign a2018 = ~a2014 & a1978;
assign a2020 = ~a2018 & ~a2016;
assign a2022 = a2020 & a1274;
assign a2024 = a1704 & l182;
assign a2026 = ~a2024 & ~a2022;
assign a2028 = ~l412 & l272;
assign a2030 = l412 & ~l272;
assign a2032 = ~a2030 & ~a2028;
assign a2034 = ~a2032 & a1732;
assign a2036 = a2032 & ~a1732;
assign a2038 = ~a2036 & ~a2034;
assign a2040 = ~l316 & l296;
assign a2042 = l316 & ~l296;
assign a2044 = ~a2042 & ~a2040;
assign a2046 = ~l332 & l216;
assign a2048 = l332 & ~l216;
assign a2050 = ~a2048 & ~a2046;
assign a2052 = a2050 & l398;
assign a2054 = ~a2050 & ~l398;
assign a2056 = ~a2054 & ~a2052;
assign a2058 = a2056 & ~a2044;
assign a2060 = ~a2056 & a2044;
assign a2062 = ~a2060 & ~a2058;
assign a2064 = l194 & l192;
assign a2066 = ~l194 & ~l192;
assign a2068 = ~a2066 & ~a2064;
assign a2070 = ~a2068 & a1960;
assign a2072 = a2068 & ~a1960;
assign a2074 = ~a2072 & ~a2070;
assign a2076 = ~a2074 & a2062;
assign a2078 = a2074 & ~a2062;
assign a2080 = ~a2078 & ~a2076;
assign a2082 = a2080 & ~a2038;
assign a2084 = ~a2080 & a2038;
assign a2086 = ~a2084 & ~a2082;
assign a2088 = a2086 & a1274;
assign a2090 = a1704 & l184;
assign a2092 = ~a2090 & ~a2088;
assign a2094 = l198 & l196;
assign a2096 = ~l198 & ~l196;
assign a2098 = ~a2096 & ~a2094;
assign a2100 = ~a2098 & l226;
assign a2102 = a2098 & ~l226;
assign a2104 = ~a2102 & ~a2100;
assign a2106 = a2104 & ~a1990;
assign a2108 = ~a2104 & a1990;
assign a2110 = ~a2108 & ~a2106;
assign a2112 = l302 & ~l276;
assign a2114 = ~l302 & l276;
assign a2116 = ~a2114 & ~a2112;
assign a2118 = ~l408 & l234;
assign a2120 = l408 & ~l234;
assign a2122 = ~a2120 & ~a2118;
assign a2124 = a2122 & ~a2116;
assign a2126 = ~a2122 & a2116;
assign a2128 = ~a2126 & ~a2124;
assign a2130 = ~a2128 & a2062;
assign a2132 = a2128 & ~a2062;
assign a2134 = ~a2132 & ~a2130;
assign a2136 = a2134 & ~a2110;
assign a2138 = ~a2134 & a2110;
assign a2140 = ~a2138 & ~a2136;
assign a2142 = a2140 & a1274;
assign a2144 = a1704 & l186;
assign a2146 = ~a2144 & ~a2142;
assign a2148 = l198 & ~l194;
assign a2150 = ~l198 & l194;
assign a2152 = ~a2150 & ~a2148;
assign a2154 = a2152 & l332;
assign a2156 = ~a2152 & ~l332;
assign a2158 = ~a2156 & ~a2154;
assign a2160 = a2158 & ~a1900;
assign a2162 = ~a2158 & a1900;
assign a2164 = ~a2162 & ~a2160;
assign a2166 = l268 & ~l258;
assign a2168 = ~l268 & l258;
assign a2170 = ~a2168 & ~a2166;
assign a2172 = ~a2170 & a1954;
assign a2174 = a2170 & ~a1954;
assign a2176 = ~a2174 & ~a2172;
assign a2178 = a2176 & ~a1810;
assign a2180 = ~a2176 & a1810;
assign a2182 = ~a2180 & ~a2178;
assign a2184 = a2182 & ~a2164;
assign a2186 = ~a2182 & a2164;
assign a2188 = ~a2186 & ~a2184;
assign a2190 = a2188 & a1274;
assign a2192 = a1704 & l188;
assign a2194 = ~a2192 & ~a2190;
assign a2196 = ~l202 & l200;
assign a2198 = l202 & ~l200;
assign a2200 = ~a2198 & ~a2196;
assign a2202 = a2200 & a2098;
assign a2204 = ~a2200 & ~a2098;
assign a2206 = ~a2204 & ~a2202;
assign a2208 = a2206 & a2068;
assign a2210 = ~a2206 & ~a2068;
assign a2212 = ~a2210 & ~a2208;
assign a2214 = ~l206 & l204;
assign a2216 = l206 & ~l204;
assign a2218 = ~a2216 & ~a2214;
assign a2220 = l210 & ~l208;
assign a2222 = ~l210 & l208;
assign a2224 = ~a2222 & ~a2220;
assign a2226 = ~a2224 & a2218;
assign a2228 = a2224 & ~a2218;
assign a2230 = ~a2228 & ~a2226;
assign a2232 = ~l214 & l212;
assign a2234 = l214 & ~l212;
assign a2236 = ~a2234 & ~a2232;
assign a2238 = l218 & ~l216;
assign a2240 = ~l218 & l216;
assign a2242 = ~a2240 & ~a2238;
assign a2244 = ~a2242 & a2236;
assign a2246 = a2242 & ~a2236;
assign a2248 = ~a2246 & ~a2244;
assign a2250 = ~a2248 & a2230;
assign a2252 = a2248 & ~a2230;
assign a2254 = ~a2252 & ~a2250;
assign a2256 = a2254 & ~a2212;
assign a2258 = ~a2254 & a2212;
assign a2260 = ~a2258 & ~a2256;
assign a2262 = a2260 & a1274;
assign a2264 = a1704 & l190;
assign a2266 = ~a2264 & ~a2262;
assign a2268 = i24 & i22;
assign a2270 = ~a2268 & i20;
assign a2274 = a2272 & ~l220;
assign a2276 = a2274 & i26;
assign a2278 = a2276 & i16;
assign a2280 = ~l222 & ~i16;
assign a2282 = a2280 & a2276;
assign a2284 = a2282 & i30;
assign a2286 = ~a2284 & ~i28;
assign a2288 = a2286 & ~a2278;
assign a2290 = a2288 & l192;
assign a2292 = a2274 & ~i16;
assign a2294 = ~a2292 & i28;
assign a2296 = a2294 & ~i20;
assign a2298 = i32 & i30;
assign a2300 = a2298 & a2296;
assign a2302 = ~a2300 & ~a2288;
assign a2304 = a2300 & l402;
assign a2306 = ~a2304 & ~a2302;
assign a2308 = a2306 & ~a2290;
assign a2310 = a2288 & l194;
assign a2312 = a2300 & l392;
assign a2314 = ~a2312 & ~a2310;
assign a2316 = a2288 & l196;
assign a2318 = a2300 & l386;
assign a2320 = ~a2318 & ~a2316;
assign a2322 = a2288 & l198;
assign a2324 = a2300 & l342;
assign a2326 = ~a2324 & ~a2302;
assign a2328 = a2326 & ~a2322;
assign a2330 = a2288 & l200;
assign a2332 = a2300 & l336;
assign a2334 = ~a2332 & ~a2302;
assign a2336 = a2334 & ~a2330;
assign a2338 = a2288 & l202;
assign a2340 = a2300 & l326;
assign a2342 = ~a2340 & ~a2302;
assign a2344 = a2342 & ~a2338;
assign a2346 = a2288 & l204;
assign a2348 = a2300 & l320;
assign a2350 = ~a2348 & ~a2302;
assign a2352 = a2350 & ~a2346;
assign a2354 = a2288 & l206;
assign a2356 = a2300 & l310;
assign a2358 = ~a2356 & ~a2302;
assign a2360 = a2358 & ~a2354;
assign a2362 = a2288 & l208;
assign a2364 = a2300 & l300;
assign a2366 = ~a2364 & ~a2362;
assign a2368 = a2288 & l210;
assign a2370 = a2300 & l290;
assign a2372 = ~a2370 & ~a2302;
assign a2374 = a2372 & ~a2368;
assign a2376 = a2288 & l212;
assign a2378 = a2300 & l284;
assign a2380 = ~a2378 & ~a2302;
assign a2382 = a2380 & ~a2376;
assign a2384 = a2288 & l214;
assign a2386 = a2300 & l266;
assign a2388 = ~a2386 & ~a2302;
assign a2390 = a2388 & ~a2384;
assign a2392 = a2288 & l216;
assign a2394 = a2300 & l256;
assign a2396 = ~a2394 & ~a2302;
assign a2398 = a2396 & ~a2392;
assign a2400 = a2288 & l218;
assign a2402 = a2300 & l224;
assign a2404 = ~a2402 & ~a2302;
assign a2406 = a2404 & ~a2400;
assign a2408 = ~a2270 & i34;
assign a2410 = a2408 & i36;
assign a2412 = a2410 & l238;
assign a2414 = ~a2410 & l222;
assign a2416 = ~a2414 & ~a2412;
assign a2418 = a2410 & l226;
assign a2420 = ~a2410 & l224;
assign a2422 = ~a2420 & ~a2418;
assign a2424 = a2288 & l226;
assign a2426 = a2300 & l228;
assign a2428 = ~a2426 & ~a2424;
assign a2430 = a2410 & l230;
assign a2432 = ~a2410 & l228;
assign a2434 = ~a2432 & ~a2430;
assign a2436 = a2288 & l230;
assign a2438 = a2300 & l232;
assign a2440 = ~a2438 & ~a2302;
assign a2442 = a2440 & ~a2436;
assign a2444 = a2410 & l234;
assign a2446 = ~a2410 & l232;
assign a2448 = ~a2446 & ~a2444;
assign a2450 = a2288 & l234;
assign a2452 = a2300 & l236;
assign a2454 = ~a2452 & ~a2302;
assign a2456 = a2454 & ~a2450;
assign a2458 = a2410 & l200;
assign a2460 = ~a2410 & l236;
assign a2462 = ~a2460 & ~a2458;
assign a2464 = ~i32 & i26;
assign a2466 = a2464 & ~i30;
assign a2468 = i24 & i20;
assign a2470 = a2468 & i36;
assign a2472 = a2292 & ~i28;
assign a2474 = a2472 & i34;
assign a2476 = a2474 & a2470;
assign a2478 = a2476 & a2466;
assign a2480 = a2478 & i38;
assign a2482 = ~a2292 & ~i28;
assign a2484 = a2482 & ~a2278;
assign a2486 = a2484 & l238;
assign a2488 = a2300 & l240;
assign a2490 = ~a2488 & ~a2486;
assign a2492 = a2490 & ~a2480;
assign a2494 = a2410 & l242;
assign a2496 = ~a2410 & l240;
assign a2498 = ~a2496 & ~a2494;
assign a2500 = ~a2484 & ~a2478;
assign a2502 = a2500 & ~a2300;
assign a2504 = a2478 & i40;
assign a2506 = a2484 & l242;
assign a2508 = a2300 & l244;
assign a2510 = ~a2508 & ~a2506;
assign a2512 = a2510 & ~a2504;
assign a2514 = a2512 & ~a2502;
assign a2516 = a2410 & l246;
assign a2518 = ~a2410 & l244;
assign a2520 = ~a2518 & ~a2516;
assign a2522 = a2478 & i42;
assign a2524 = a2484 & l246;
assign a2526 = a2300 & l248;
assign a2528 = ~a2526 & ~a2524;
assign a2530 = a2528 & ~a2522;
assign a2532 = a2530 & ~a2502;
assign a2534 = a2410 & l250;
assign a2536 = ~a2410 & l248;
assign a2538 = ~a2536 & ~a2534;
assign a2540 = a2484 & l250;
assign a2542 = a2300 & l252;
assign a2544 = ~a2542 & ~a2540;
assign a2546 = a2544 & ~a2502;
assign a2548 = a2410 & l254;
assign a2550 = ~a2410 & l252;
assign a2552 = ~a2550 & ~a2548;
assign a2554 = a2484 & l254;
assign a2556 = a2300 & i44;
assign a2558 = ~a2556 & ~a2554;
assign a2560 = a2558 & ~a2502;
assign a2562 = a2410 & l258;
assign a2564 = ~a2410 & l256;
assign a2566 = ~a2564 & ~a2562;
assign a2568 = a2288 & l258;
assign a2570 = a2300 & l260;
assign a2572 = ~a2570 & ~a2302;
assign a2574 = a2572 & ~a2568;
assign a2576 = a2410 & l262;
assign a2578 = ~a2410 & l260;
assign a2580 = ~a2578 & ~a2576;
assign a2582 = a2288 & l262;
assign a2584 = a2300 & l264;
assign a2586 = ~a2584 & ~a2302;
assign a2588 = a2586 & ~a2582;
assign a2590 = a2410 & l198;
assign a2592 = ~a2410 & l264;
assign a2594 = ~a2592 & ~a2590;
assign a2596 = a2410 & l268;
assign a2598 = ~a2410 & l266;
assign a2600 = ~a2598 & ~a2596;
assign a2602 = a2288 & l268;
assign a2604 = a2300 & l270;
assign a2606 = ~a2604 & ~a2602;
assign a2608 = a2410 & l272;
assign a2610 = ~a2410 & l270;
assign a2612 = ~a2610 & ~a2608;
assign a2614 = a2288 & l272;
assign a2616 = a2300 & l274;
assign a2618 = ~a2616 & ~a2302;
assign a2620 = a2618 & ~a2614;
assign a2622 = a2410 & l276;
assign a2624 = ~a2410 & l274;
assign a2626 = ~a2624 & ~a2622;
assign a2628 = a2288 & l276;
assign a2630 = a2300 & l278;
assign a2632 = ~a2630 & ~a2302;
assign a2634 = a2632 & ~a2628;
assign a2636 = a2410 & l280;
assign a2638 = ~a2410 & l278;
assign a2640 = ~a2638 & ~a2636;
assign a2642 = a2288 & l280;
assign a2644 = a2300 & l282;
assign a2646 = ~a2644 & ~a2302;
assign a2648 = a2646 & ~a2642;
assign a2650 = a2410 & l192;
assign a2652 = ~a2410 & l282;
assign a2654 = ~a2652 & ~a2650;
assign a2656 = a2410 & l286;
assign a2658 = ~a2410 & l284;
assign a2660 = ~a2658 & ~a2656;
assign a2662 = a2288 & l286;
assign a2664 = a2300 & l288;
assign a2666 = ~a2664 & ~a2662;
assign a2668 = a2410 & l216;
assign a2670 = ~a2410 & l288;
assign a2672 = ~a2670 & ~a2668;
assign a2674 = a2410 & l292;
assign a2676 = ~a2410 & l290;
assign a2678 = ~a2676 & ~a2674;
assign a2680 = a2288 & l292;
assign a2682 = a2300 & l294;
assign a2684 = ~a2682 & ~a2302;
assign a2686 = a2684 & ~a2680;
assign a2688 = a2410 & l296;
assign a2690 = ~a2410 & l294;
assign a2692 = ~a2690 & ~a2688;
assign a2694 = a2288 & l296;
assign a2696 = a2300 & l298;
assign a2698 = ~a2696 & ~a2694;
assign a2700 = a2410 & l206;
assign a2702 = ~a2410 & l298;
assign a2704 = ~a2702 & ~a2700;
assign a2706 = a2410 & l302;
assign a2708 = ~a2410 & l300;
assign a2710 = ~a2708 & ~a2706;
assign a2712 = a2288 & l302;
assign a2714 = a2300 & l304;
assign a2716 = ~a2714 & ~a2302;
assign a2718 = a2716 & ~a2712;
assign a2720 = a2410 & l306;
assign a2722 = ~a2410 & l304;
assign a2724 = ~a2722 & ~a2720;
assign a2726 = a2288 & l306;
assign a2728 = a2300 & l308;
assign a2730 = ~a2728 & ~a2726;
assign a2732 = a2410 & l210;
assign a2734 = ~a2410 & l308;
assign a2736 = ~a2734 & ~a2732;
assign a2738 = a2410 & l312;
assign a2740 = ~a2410 & l310;
assign a2742 = ~a2740 & ~a2738;
assign a2744 = a2288 & l312;
assign a2746 = a2300 & l314;
assign a2748 = ~a2746 & ~a2302;
assign a2750 = a2748 & ~a2744;
assign a2752 = a2410 & l316;
assign a2754 = ~a2410 & l314;
assign a2756 = ~a2754 & ~a2752;
assign a2758 = a2288 & l316;
assign a2760 = a2300 & l318;
assign a2762 = ~a2760 & ~a2758;
assign a2764 = a2410 & l202;
assign a2766 = ~a2410 & l318;
assign a2768 = ~a2766 & ~a2764;
assign a2770 = a2410 & l322;
assign a2772 = ~a2410 & l320;
assign a2774 = ~a2772 & ~a2770;
assign a2776 = a2288 & l322;
assign a2778 = a2300 & l324;
assign a2780 = ~a2778 & ~a2302;
assign a2782 = a2780 & ~a2776;
assign a2784 = a2410 & l194;
assign a2786 = ~a2410 & l324;
assign a2788 = ~a2786 & ~a2784;
assign a2790 = a2410 & l328;
assign a2792 = ~a2410 & l326;
assign a2794 = ~a2792 & ~a2790;
assign a2796 = a2288 & l328;
assign a2798 = a2300 & l330;
assign a2800 = ~a2798 & ~a2302;
assign a2802 = a2800 & ~a2796;
assign a2804 = a2410 & l332;
assign a2806 = ~a2410 & l330;
assign a2808 = ~a2806 & ~a2804;
assign a2810 = a2288 & l332;
assign a2812 = a2300 & l334;
assign a2814 = ~a2812 & ~a2302;
assign a2816 = a2814 & ~a2810;
assign a2818 = a2410 & l204;
assign a2820 = ~a2410 & l334;
assign a2822 = ~a2820 & ~a2818;
assign a2824 = a2410 & l338;
assign a2826 = ~a2410 & l336;
assign a2828 = ~a2826 & ~a2824;
assign a2830 = a2288 & l338;
assign a2832 = a2300 & l340;
assign a2834 = ~a2832 & ~a2302;
assign a2836 = a2834 & ~a2830;
assign a2838 = a2410 & l196;
assign a2840 = ~a2410 & l340;
assign a2842 = ~a2840 & ~a2838;
assign a2844 = a2410 & l344;
assign a2846 = ~a2410 & l342;
assign a2848 = ~a2846 & ~a2844;
assign a2850 = ~i48 & ~i46;
assign a2852 = ~i52 & ~i50;
assign a2854 = a2852 & a2850;
assign a2856 = i58 & i56;
assign a2858 = a2856 & i54;
assign a2860 = i64 & ~i62;
assign a2862 = a2860 & ~i60;
assign a2864 = a2862 & ~a2858;
assign a2866 = a2864 & a2854;
assign a2868 = ~a2866 & a2478;
assign a2870 = a2484 & l344;
assign a2872 = a2300 & l346;
assign a2874 = ~a2872 & ~a2870;
assign a2876 = a2874 & ~a2868;
assign a2878 = a2876 & ~a2502;
assign a2880 = a2410 & l348;
assign a2882 = ~a2410 & l346;
assign a2884 = ~a2882 & ~a2880;
assign a2886 = a2478 & i66;
assign a2888 = a2484 & l348;
assign a2890 = a2300 & l350;
assign a2892 = ~a2890 & ~a2888;
assign a2894 = a2892 & ~a2886;
assign a2896 = a2410 & l352;
assign a2898 = ~a2410 & l350;
assign a2900 = ~a2898 & ~a2896;
assign a2902 = a2484 & l352;
assign a2904 = a2300 & l354;
assign a2906 = ~a2904 & ~a2902;
assign a2908 = a2906 & ~a2502;
assign a2910 = a2410 & l356;
assign a2912 = ~a2410 & l354;
assign a2914 = ~a2912 & ~a2910;
assign a2916 = a2484 & l356;
assign a2918 = a2300 & l358;
assign a2920 = ~a2918 & ~a2916;
assign a2922 = a2920 & ~a2502;
assign a2924 = a2410 & l360;
assign a2926 = ~a2410 & l358;
assign a2928 = ~a2926 & ~a2924;
assign a2930 = a2484 & l360;
assign a2932 = a2300 & l362;
assign a2934 = ~a2932 & ~a2930;
assign a2936 = a2934 & ~a2502;
assign a2938 = a2410 & l364;
assign a2940 = ~a2410 & l362;
assign a2942 = ~a2940 & ~a2938;
assign a2944 = a2484 & l364;
assign a2946 = a2300 & l366;
assign a2948 = ~a2946 & ~a2944;
assign a2950 = a2948 & ~a2502;
assign a2952 = a2410 & l368;
assign a2954 = ~a2410 & l366;
assign a2956 = ~a2954 & ~a2952;
assign a2958 = a2484 & l368;
assign a2960 = a2300 & l370;
assign a2962 = ~a2960 & ~a2958;
assign a2964 = a2962 & ~a2502;
assign a2966 = a2410 & l372;
assign a2968 = ~a2410 & l370;
assign a2970 = ~a2968 & ~a2966;
assign a2972 = a2484 & l372;
assign a2974 = a2300 & l374;
assign a2976 = ~a2974 & ~a2972;
assign a2978 = a2410 & l376;
assign a2980 = ~a2410 & l374;
assign a2982 = ~a2980 & ~a2978;
assign a2984 = a2484 & l376;
assign a2986 = a2300 & l378;
assign a2988 = ~a2986 & ~a2984;
assign a2990 = a2988 & ~a2502;
assign a2992 = a2410 & l380;
assign a2994 = ~a2410 & l378;
assign a2996 = ~a2994 & ~a2992;
assign a2998 = a2484 & l380;
assign a3000 = a2300 & l382;
assign a3002 = ~a3000 & ~a2998;
assign a3004 = a3002 & ~a2502;
assign a3006 = a2410 & l384;
assign a3008 = ~a2410 & l382;
assign a3010 = ~a3008 & ~a3006;
assign a3012 = a2484 & l384;
assign a3014 = a2300 & l222;
assign a3016 = ~a3014 & ~a3012;
assign a3018 = a3016 & ~a2502;
assign a3020 = a2410 & l388;
assign a3022 = ~a2410 & l386;
assign a3024 = ~a3022 & ~a3020;
assign a3026 = a2288 & l388;
assign a3028 = a2300 & l390;
assign a3030 = ~a3028 & ~a2302;
assign a3032 = a3030 & ~a3026;
assign a3034 = a2410 & l208;
assign a3036 = ~a2410 & l390;
assign a3038 = ~a3036 & ~a3034;
assign a3040 = a2410 & l394;
assign a3042 = ~a2410 & l392;
assign a3044 = ~a3042 & ~a3040;
assign a3046 = a2288 & l394;
assign a3048 = a2300 & l396;
assign a3050 = ~a3048 & ~a2302;
assign a3052 = a3050 & ~a3046;
assign a3054 = a2410 & l398;
assign a3056 = ~a2410 & l396;
assign a3058 = ~a3056 & ~a3054;
assign a3060 = a2288 & l398;
assign a3062 = a2300 & l400;
assign a3064 = ~a3062 & ~a2302;
assign a3066 = a3064 & ~a3060;
assign a3068 = a2410 & l212;
assign a3070 = ~a2410 & l400;
assign a3072 = ~a3070 & ~a3068;
assign a3074 = a2410 & l404;
assign a3076 = ~a2410 & l402;
assign a3078 = ~a3076 & ~a3074;
assign a3080 = a2288 & l404;
assign a3082 = a2300 & l406;
assign a3084 = ~a3082 & ~a2302;
assign a3086 = a3084 & ~a3080;
assign a3088 = a2410 & l218;
assign a3090 = ~a2410 & l406;
assign a3092 = ~a3090 & ~a3088;
assign a3094 = a2288 & l408;
assign a3096 = a2300 & l410;
assign a3098 = ~a3096 & ~a2302;
assign a3100 = a3098 & ~a3094;
assign a3102 = a2410 & l214;
assign a3104 = ~a2410 & l410;
assign a3106 = ~a3104 & ~a3102;
assign a3108 = a2288 & l412;
assign a3110 = a2300 & l414;
assign a3112 = ~a3110 & ~a2302;
assign a3114 = a3112 & ~a3108;
assign a3116 = a2410 & l408;
assign a3118 = ~a2410 & l414;
assign a3120 = ~a3118 & ~a3116;
assign a3122 = a2288 & l416;
assign a3124 = a2300 & l418;
assign a3126 = ~a3124 & ~a3122;
assign a3128 = a2410 & l412;
assign a3130 = ~a2410 & l418;
assign a3132 = ~a3130 & ~a3128;
assign a3134 = a2288 & l420;
assign a3136 = a2300 & l422;
assign a3138 = ~a3136 & ~a2302;
assign a3140 = a3138 & ~a3134;
assign a3142 = a2410 & l424;
assign a3144 = ~a2410 & l422;
assign a3146 = ~a3144 & ~a3142;
assign a3148 = a2288 & l424;
assign a3150 = a2300 & l426;
assign a3152 = ~a3150 & ~a2302;
assign a3154 = a3152 & ~a3148;
assign a3156 = a2410 & l416;
assign a3158 = ~a2410 & l426;
assign a3160 = ~a3158 & ~a3156;
assign a3162 = a2288 & l428;
assign a3164 = a2300 & l430;
assign a3166 = ~a3164 & ~a2302;
assign a3168 = a3166 & ~a3162;
assign a3170 = a2410 & l420;
assign a3172 = ~a2410 & l430;
assign a3174 = ~a3172 & ~a3170;
assign a3176 = a1704 & l432;
assign a3178 = a1194 & l112;
assign a3180 = a1274 & l276;
assign a3182 = ~a3180 & ~a3178;
assign a3184 = a3182 & ~a3176;
assign a3186 = a1704 & l434;
assign a3188 = a1194 & l120;
assign a3190 = a1274 & l296;
assign a3192 = ~a3190 & ~a3188;
assign a3194 = a3192 & ~a3186;
assign a3196 = a1704 & l436;
assign a3198 = a1194 & l118;
assign a3200 = a1274 & l206;
assign a3202 = ~a3200 & ~a3198;
assign a3204 = a3202 & ~a3196;
assign p0 = a470;

assert property (~p0);

endmodule
