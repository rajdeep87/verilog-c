module m6s17 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134;

output p0;

wire na404,na418,na502,na566,na578,na590,na602,na614,na646,na658,na670,na706,na712,na718,na724,
na1724,na1764,na1770,na1888,na1908,na1932,na1952,na1958,na1976,na1982,na1990,na2000,na2006,na2012,na2018,
na2024,na2030,na2036,na2042,na2048,na2054,na2060,na2066,na2072,na2078,na2086,na2092,na2098,na2106,na2112,
na2118,na2138,na2144,na2402,na2418,na2718,na2724,na2750,na2754,na2758,na2762,na2766,na2772,na2778,na2784,
na2790,na2796,na2802,na2808,na2814,na2820,na2824,na2830,na2836,na2842,na2848,na2854,na2858,na2864,na2868,
na2876,na2884,na2892,na2900,na2906,na2912,na2918,na2924,na2190,na2958,na2316,na2970,na2976,na2986,na2998,
a4188,c1,na4194,a4374,a4510,a4586,a4672,a4708,a4784,a4830,a4866,na4872,na4884,na4890,na4902,
na4914,na4926,na4938,na4950,na4962,a4964,a4986,a4992,a5304,a5336,a5366,a5368,a5376,na5392,na5416,
a5418,a5422,a5428,a5432,a5458,a5486,na5494,a392,a394,a396,a398,a400,a402,a404,a406,
a408,a410,a412,a414,a416,a418,a420,a422,a424,a426,a428,a430,a432,a434,a436,
a438,a440,a442,a444,a446,a448,a450,a452,a454,a456,a458,a460,a462,a464,a466,
a468,a470,a472,a474,a476,a478,a480,a482,a484,a486,a488,a490,a492,a494,a496,
a498,a500,a502,a504,a506,a508,a510,a512,a514,a516,a518,a520,a522,a524,a526,
a528,a530,a532,a534,a536,a538,a540,a542,a544,a546,a548,a550,a552,a554,a556,
a558,a560,a562,a564,a566,a568,a570,a572,a574,a576,a578,a580,a582,a584,a586,
a588,a590,a592,a594,a596,a598,a600,a602,a604,a606,a608,a610,a612,a614,a616,
a618,a620,a622,a624,a626,a628,a630,a632,a634,a636,a638,a640,a642,a644,a646,
a648,a650,a652,a654,a656,a658,a660,a662,a664,a666,a668,a670,a672,a674,a676,
a678,a680,a682,a684,a686,a688,a690,a692,a694,a696,a698,a700,a702,a704,a706,
a708,a710,a712,a714,a716,a718,a720,a722,a724,a726,a728,a730,a732,a734,a736,
a738,a740,a742,a744,a746,a748,a750,a752,a754,a756,a758,a760,a762,a764,a766,
a768,a770,a772,a774,a776,a778,a780,a782,a784,a786,a788,a790,a792,a794,a796,
a798,a800,a802,a804,a806,a808,a810,a812,a814,a816,a818,a820,a822,a824,a826,
a828,a830,a832,a834,a836,a838,a840,a842,a844,a846,a848,a850,a852,a854,a856,
a858,a860,a862,a864,a866,a868,a870,a872,a874,a876,a878,a880,a882,a884,a886,
a888,a890,a892,a894,a896,a898,a900,a902,a904,a906,a908,a910,a912,a914,a916,
a918,a920,a922,a924,a926,a928,a930,a932,a934,a936,a938,a940,a942,a944,a946,
a948,a950,a952,a954,a956,a958,a960,a962,a964,a966,a968,a970,a972,a974,a976,
a978,a980,a982,a984,a986,a988,a990,a992,a994,a996,a998,a1000,a1002,a1004,a1006,
a1008,a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,
a1038,a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,a1062,a1064,a1066,
a1068,a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,a1092,a1094,a1096,
a1098,a1100,a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,a1124,a1126,
a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,a1154,a1156,
a1158,a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,a1178,a1180,a1182,a1184,a1186,
a1188,a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,
a1218,a1220,a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,
a1248,a1250,a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,a1268,a1270,a1272,a1274,a1276,
a1278,a1280,a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,
a1308,a1310,a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,a1334,a1336,
a1338,a1340,a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,
a1368,a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,a1388,a1390,a1392,a1394,a1396,
a1398,a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1426,
a1428,a1430,a1432,a1434,a1436,a1438,a1440,a1442,a1444,a1446,a1448,a1450,a1452,a1454,a1456,
a1458,a1460,a1462,a1464,a1466,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1482,a1484,a1486,
a1488,a1490,a1492,a1494,a1496,a1498,a1500,a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,
a1518,a1520,a1522,a1524,a1526,a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,
a1548,a1550,a1552,a1554,a1556,a1558,a1560,a1562,a1564,a1566,a1568,a1570,a1572,a1574,a1576,
a1578,a1580,a1582,a1584,a1586,a1588,a1590,a1592,a1594,a1596,a1598,a1600,a1602,a1604,a1606,
a1608,a1610,a1612,a1614,a1616,a1618,a1620,a1622,a1624,a1626,a1628,a1630,a1632,a1634,a1636,
a1638,a1640,a1642,a1644,a1646,a1648,a1650,a1652,a1654,a1656,a1658,a1660,a1662,a1664,a1666,
a1668,a1670,a1672,a1674,a1676,a1678,a1680,a1682,a1684,a1686,a1688,a1690,a1692,a1694,a1696,
a1698,a1700,a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,
a1728,a1730,a1732,a1734,a1736,a1738,a1740,a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,
a1758,a1760,a1762,a1764,a1766,a1768,a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,
a1788,a1790,a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,
a1818,a1820,a1822,a1824,a1826,a1828,a1830,a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,
a1848,a1850,a1852,a1854,a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,
a1878,a1880,a1882,a1884,a1886,a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,
a1908,a1910,a1912,a1914,a1916,a1918,a1920,a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,
a1938,a1940,a1942,a1944,a1946,a1948,a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,
a1968,a1970,a1972,a1974,a1976,a1978,a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,
a1998,a2000,a2002,a2004,a2006,a2008,a2010,a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,
a2028,a2030,a2032,a2034,a2036,a2038,a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,
a2058,a2060,a2062,a2064,a2066,a2068,a2070,a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,
a2088,a2090,a2092,a2094,a2096,a2098,a2100,a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,
a2118,a2120,a2122,a2124,a2126,a2128,a2130,a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,
a2148,a2150,a2152,a2154,a2156,a2158,a2160,a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,
a2178,a2180,a2182,a2184,a2186,a2188,a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,
a2208,a2210,a2212,a2214,a2216,a2218,a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,
a2238,a2240,a2242,a2244,a2246,a2248,a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,
a2268,a2270,a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,
a2298,a2300,a2302,a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,
a2328,a2330,a2332,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,
a2358,a2360,a2362,a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,
a2388,a2390,a2392,a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,
a2418,a2420,a2422,a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,
a2448,a2450,a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,
a2478,a2480,a2482,a2484,a2486,a2488,a2490,a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,
a2508,a2510,a2512,a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,
a2538,a2540,a2542,a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,
a2568,a2570,a2572,a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,
a2598,a2600,a2602,a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,
a2628,a2630,a2632,a2634,a2636,a2638,a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,
a2658,a2660,a2662,a2664,a2666,a2668,a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,
a2688,a2690,a2692,a2694,a2696,a2698,a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,
a2718,a2720,a2722,a2724,a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,
a2748,a2750,a2752,a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,
a2778,a2780,a2782,a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,
a2808,a2810,a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,
a2838,a2840,a2842,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,
a2868,a2870,a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,
a2898,a2900,a2902,a2904,a2906,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,
a2928,a2930,a2932,a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,
a2958,a2960,a2962,a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,
a2988,a2990,a2992,a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,
a3018,a3020,a3022,a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,
a3048,a3050,a3052,a3054,a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,
a3078,a3080,a3082,a3084,a3086,a3088,a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,
a3108,a3110,a3112,a3114,a3116,a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,
a3138,a3140,a3142,a3144,a3146,a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,
a3168,a3170,a3172,a3174,a3176,a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,
a3198,a3200,a3202,a3204,a3206,a3208,a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,
a3228,a3230,a3232,a3234,a3236,a3238,a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,
a3258,a3260,a3262,a3264,a3266,a3268,a3270,a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,
a3288,a3290,a3292,a3294,a3296,a3298,a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,
a3318,a3320,a3322,a3324,a3326,a3328,a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,
a3348,a3350,a3352,a3354,a3356,a3358,a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,
a3378,a3380,a3382,a3384,a3386,a3388,a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,
a3408,a3410,a3412,a3414,a3416,a3418,a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,
a3438,a3440,a3442,a3444,a3446,a3448,a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,
a3468,a3470,a3472,a3474,a3476,a3478,a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,
a3498,a3500,a3502,a3504,a3506,a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,
a3528,a3530,a3532,a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,
a3558,a3560,a3562,a3564,a3566,a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,
a3588,a3590,a3592,a3594,a3596,a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,
a3618,a3620,a3622,a3624,a3626,a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,
a3648,a3650,a3652,a3654,a3656,a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,
a3678,a3680,a3682,a3684,a3686,a3688,a3690,a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,
a3708,a3710,a3712,a3714,a3716,a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,
a3738,a3740,a3742,a3744,a3746,a3748,a3750,a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,
a3768,a3770,a3772,a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,
a3798,a3800,a3802,a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,
a3828,a3830,a3832,a3834,a3836,a3838,a3840,a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,
a3858,a3860,a3862,a3864,a3866,a3868,a3870,a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,
a3888,a3890,a3892,a3894,a3896,a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,
a3918,a3920,a3922,a3924,a3926,a3928,a3930,a3932,a3934,a3936,a3938,a3940,a3942,a3944,a3946,
a3948,a3950,a3952,a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,
a3978,a3980,a3982,a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,
a4008,a4010,a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,
a4038,a4040,a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,
a4068,a4070,a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,a4096,
a4098,a4100,a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4124,a4126,
a4128,a4130,a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,a4152,a4154,a4156,
a4158,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,a4184,a4186,
a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,a4214,a4216,a4218,
a4220,a4222,a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,a4244,a4246,a4248,
a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,a4274,a4276,a4278,
a4280,a4282,a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,a4306,a4308,
a4310,a4312,a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,a4334,a4336,a4338,
a4340,a4342,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,a4368,
a4370,a4372,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,a4394,a4396,a4398,a4400,
a4402,a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,
a4432,a4434,a4436,a4438,a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,a4458,a4460,
a4462,a4464,a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4482,a4484,a4486,a4488,a4490,
a4492,a4494,a4496,a4498,a4500,a4502,a4504,a4506,a4508,a4512,a4514,a4516,a4518,a4520,a4522,
a4524,a4526,a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,
a4554,a4556,a4558,a4560,a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,a4578,a4580,a4582,
a4584,a4588,a4590,a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,a4612,a4614,
a4616,a4618,a4620,a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,a4642,a4644,
a4646,a4648,a4650,a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,a4674,a4676,
a4678,a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,a4696,a4698,a4700,a4702,a4704,a4706,
a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,a4726,a4728,a4730,a4732,a4734,a4736,a4738,
a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,a4756,a4758,a4760,a4762,a4764,a4766,a4768,
a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4786,a4788,a4790,a4792,a4794,a4796,a4798,a4800,
a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,a4818,a4820,a4822,a4824,a4826,a4828,a4832,
a4834,a4836,a4838,a4840,a4842,a4844,a4846,a4848,a4850,a4852,a4854,a4856,a4858,a4860,a4862,
a4864,a4868,a4870,a4872,a4874,a4876,a4878,a4880,a4882,a4884,a4886,a4888,a4890,a4892,a4894,
a4896,a4898,a4900,a4902,a4904,a4906,a4908,a4910,a4912,a4914,a4916,a4918,a4920,a4922,a4924,
a4926,a4928,a4930,a4932,a4934,a4936,a4938,a4940,a4942,a4944,a4946,a4948,a4950,a4952,a4954,
a4956,a4958,a4960,a4962,a4966,a4968,a4970,a4972,a4974,a4976,a4978,a4980,a4982,a4984,a4988,
a4990,a4994,a4996,a4998,a5000,a5002,a5004,a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,
a5022,a5024,a5026,a5028,a5030,a5032,a5034,a5036,a5038,a5040,a5042,a5044,a5046,a5048,a5050,
a5052,a5054,a5056,a5058,a5060,a5062,a5064,a5066,a5068,a5070,a5072,a5074,a5076,a5078,a5080,
a5082,a5084,a5086,a5088,a5090,a5092,a5094,a5096,a5098,a5100,a5102,a5104,a5106,a5108,a5110,
a5112,a5114,a5116,a5118,a5120,a5122,a5124,a5126,a5128,a5130,a5132,a5134,a5136,a5138,a5140,
a5142,a5144,a5146,a5148,a5150,a5152,a5154,a5156,a5158,a5160,a5162,a5164,a5166,a5168,a5170,
a5172,a5174,a5176,a5178,a5180,a5182,a5184,a5186,a5188,a5190,a5192,a5194,a5196,a5198,a5200,
a5202,a5204,a5206,a5208,a5210,a5212,a5214,a5216,a5218,a5220,a5222,a5224,a5226,a5228,a5230,
a5232,a5234,a5236,a5238,a5240,a5242,a5244,a5246,a5248,a5250,a5252,a5254,a5256,a5258,a5260,
a5262,a5264,a5266,a5268,a5270,a5272,a5274,a5276,a5278,a5280,a5282,a5284,a5286,a5288,a5290,
a5292,a5294,a5296,a5298,a5300,a5302,a5306,a5308,a5310,a5312,a5314,a5316,a5318,a5320,a5322,
a5324,a5326,a5328,a5330,a5332,a5334,a5338,a5340,a5342,a5344,a5346,a5348,a5350,a5352,a5354,
a5356,a5358,a5360,a5362,a5364,a5370,a5372,a5374,a5378,a5380,a5382,a5384,a5386,a5388,a5390,
a5392,a5394,a5396,a5398,a5400,a5402,a5404,a5406,a5408,a5410,a5412,a5414,a5416,a5420,a5424,
a5426,a5430,a5434,a5436,a5438,a5440,a5442,a5444,a5446,a5448,a5450,a5452,a5454,a5456,a5460,
a5462,a5464,a5466,a5468,a5470,a5472,a5474,a5476,a5478,a5480,a5482,a5484,a5488,a5490,a5492,
a5494,a5496,a5498,a5500,a5502,a5504,a5506,a5508,a5510,a5512,a5514,a5516,a5518,a5520,a5522,
a5524,a5526,a5528,a5530,a5532,a5534,a5536,a5538,a5540,a5542,a5544,a5546,a5548,a5550,a5552,
a5554,a5556,a5558,a5560,a5562,p0;

reg l136,l138,l140,l142,l144,l146,l148,l150,l152,l154,l156,l158,l160,l162,l164,
l166,l168,l170,l172,l174,l176,l178,l180,l182,l184,l186,l188,l190,l192,l194,
l196,l198,l200,l202,l204,l206,l208,l210,l212,l214,l216,l218,l220,l222,l224,
l226,l228,l230,l232,l234,l236,l238,l240,l242,l244,l246,l248,l250,l252,l254,
l256,l258,l260,l262,l264,l266,l268,l270,l272,l274,l276,l278,l280,l282,l284,
l286,l288,l290,l292,l294,l296,l298,l300,l302,l304,l306,l308,l310,l312,l314,
l316,l318,l320,l322,l324,l326,l328,l330,l332,l334,l336,l338,l340,l342,l344,
l346,l348,l350,l352,l354,l356,l358,l360,l362,l364,l366,l368,l370,l372,l374,
l376,l378,l380,l382,l384,l386,l388,l390;

initial
begin
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
end

always @(posedge na404)
   l136 <= na404;

always @(posedge na418)
   l138 <= na418;

always @(posedge na502)
   l140 <= na502;

always @(posedge na566)
   l142 <= na566;

always @(posedge na578)
   l144 <= na578;

always @(posedge na590)
   l146 <= na590;

always @(posedge na602)
   l148 <= na602;

always @(posedge na614)
   l150 <= na614;

always @(posedge na646)
   l152 <= na646;

always @(posedge na658)
   l154 <= na658;

always @(posedge na670)
   l156 <= na670;

always @(posedge na706)
   l158 <= na706;

always @(posedge na712)
   l160 <= na712;

always @(posedge na718)
   l162 <= na718;

always @(posedge na724)
   l164 <= na724;

always @(posedge na1724)
   l166 <= na1724;

always @(posedge na1764)
   l168 <= na1764;

always @(posedge na1770)
   l170 <= na1770;

always @(posedge na1888)
   l172 <= na1888;

always @(posedge na1908)
   l174 <= na1908;

always @(posedge na1932)
   l176 <= na1932;

always @(posedge na1952)
   l178 <= na1952;

always @(posedge na1958)
   l180 <= na1958;

always @(posedge na1976)
   l182 <= na1976;

always @(posedge na1982)
   l184 <= na1982;

always @(posedge na1990)
   l186 <= na1990;

always @(posedge na2000)
   l188 <= na2000;

always @(posedge na2006)
   l190 <= na2006;

always @(posedge na2012)
   l192 <= na2012;

always @(posedge na2018)
   l194 <= na2018;

always @(posedge na2024)
   l196 <= na2024;

always @(posedge na2030)
   l198 <= na2030;

always @(posedge na2036)
   l200 <= na2036;

always @(posedge na2042)
   l202 <= na2042;

always @(posedge na2048)
   l204 <= na2048;

always @(posedge na2054)
   l206 <= na2054;

always @(posedge na2060)
   l208 <= na2060;

always @(posedge na2066)
   l210 <= na2066;

always @(posedge na2072)
   l212 <= na2072;

always @(posedge na2078)
   l214 <= na2078;

always @(posedge na2086)
   l216 <= na2086;

always @(posedge na2092)
   l218 <= na2092;

always @(posedge na2098)
   l220 <= na2098;

always @(posedge na2106)
   l222 <= na2106;

always @(posedge na2112)
   l224 <= na2112;

always @(posedge na2118)
   l226 <= na2118;

always @(posedge na2138)
   l228 <= na2138;

always @(posedge na2144)
   l230 <= na2144;

always @(posedge na2402)
   l232 <= na2402;

always @(posedge na2418)
   l234 <= na2418;

always @(posedge na2718)
   l236 <= na2718;

always @(posedge na2724)
   l238 <= na2724;

always @(posedge na2750)
   l240 <= na2750;

always @(posedge i16)
   l242 <= i16;

always @(posedge na2754)
   l244 <= na2754;

always @(posedge na2758)
   l246 <= na2758;

always @(posedge na2762)
   l248 <= na2762;

always @(posedge na2766)
   l250 <= na2766;

always @(posedge na2772)
   l252 <= na2772;

always @(posedge na2778)
   l254 <= na2778;

always @(posedge na2784)
   l256 <= na2784;

always @(posedge na2790)
   l258 <= na2790;

always @(posedge na2796)
   l260 <= na2796;

always @(posedge na2802)
   l262 <= na2802;

always @(posedge na2808)
   l264 <= na2808;

always @(posedge na2814)
   l266 <= na2814;

always @(posedge na2820)
   l268 <= na2820;

always @(posedge na2824)
   l270 <= na2824;

always @(posedge na2830)
   l272 <= na2830;

always @(posedge na2836)
   l274 <= na2836;

always @(posedge na2842)
   l276 <= na2842;

always @(posedge na2848)
   l278 <= na2848;

always @(posedge na2854)
   l280 <= na2854;

always @(posedge na2858)
   l282 <= na2858;

always @(posedge na2864)
   l284 <= na2864;

always @(posedge na2868)
   l286 <= na2868;

always @(posedge na2876)
   l288 <= na2876;

always @(posedge na2884)
   l290 <= na2884;

always @(posedge na2892)
   l292 <= na2892;

always @(posedge na2900)
   l294 <= na2900;

always @(posedge na2906)
   l296 <= na2906;

always @(posedge na2912)
   l298 <= na2912;

always @(posedge na2918)
   l300 <= na2918;

always @(posedge na2924)
   l302 <= na2924;

always @(posedge na2190)
   l304 <= na2190;

always @(posedge na2958)
   l306 <= na2958;

always @(posedge na2316)
   l308 <= na2316;

always @(posedge na2970)
   l310 <= na2970;

always @(posedge na2976)
   l312 <= na2976;

always @(posedge na2986)
   l314 <= na2986;

always @(posedge na2998)
   l316 <= na2998;

always @(posedge a4188)
   l318 <= a4188;

always @(posedge c1)
   l320 <= c1;

always @(posedge na4194)
   l322 <= na4194;

always @(posedge a4374)
   l324 <= a4374;

always @(posedge a4510)
   l326 <= a4510;

always @(posedge a4586)
   l328 <= a4586;

always @(posedge a4672)
   l330 <= a4672;

always @(posedge a4708)
   l332 <= a4708;

always @(posedge a4784)
   l334 <= a4784;

always @(posedge a4830)
   l336 <= a4830;

always @(posedge a4866)
   l338 <= a4866;

always @(posedge na4872)
   l340 <= na4872;

always @(posedge na4884)
   l342 <= na4884;

always @(posedge na4890)
   l344 <= na4890;

always @(posedge na4902)
   l346 <= na4902;

always @(posedge na4914)
   l348 <= na4914;

always @(posedge na4926)
   l350 <= na4926;

always @(posedge na4938)
   l352 <= na4938;

always @(posedge na4950)
   l354 <= na4950;

always @(posedge na4962)
   l356 <= na4962;

always @(posedge a4964)
   l358 <= a4964;

always @(posedge a4986)
   l360 <= a4986;

always @(posedge a4992)
   l362 <= a4992;

always @(posedge a5304)
   l364 <= a5304;

always @(posedge a5336)
   l366 <= a5336;

always @(posedge a5366)
   l368 <= a5366;

always @(posedge a5368)
   l370 <= a5368;

always @(posedge a5376)
   l372 <= a5376;

always @(posedge na5392)
   l374 <= na5392;

always @(posedge na5416)
   l376 <= na5416;

always @(posedge a5418)
   l378 <= a5418;

always @(posedge a5422)
   l380 <= a5422;

always @(posedge a5428)
   l382 <= a5428;

always @(posedge a5432)
   l384 <= a5432;

always @(posedge a5458)
   l386 <= a5458;

always @(posedge a5486)
   l388 <= a5486;

always @(posedge na5494)
   l390 <= na5494;


assign na404 = ~a404;
assign na418 = ~a418;
assign na502 = ~a502;
assign na566 = ~a566;
assign na578 = ~a578;
assign na590 = ~a590;
assign na602 = ~a602;
assign na614 = ~a614;
assign na646 = ~a646;
assign na658 = ~a658;
assign na670 = ~a670;
assign na706 = ~a706;
assign na712 = ~a712;
assign na718 = ~a718;
assign na724 = ~a724;
assign na1724 = ~a1724;
assign na1764 = ~a1764;
assign na1770 = ~a1770;
assign na1888 = ~a1888;
assign na1908 = ~a1908;
assign na1932 = ~a1932;
assign na1952 = ~a1952;
assign na1958 = ~a1958;
assign na1976 = ~a1976;
assign na1982 = ~a1982;
assign na1990 = ~a1990;
assign na2000 = ~a2000;
assign na2006 = ~a2006;
assign na2012 = ~a2012;
assign na2018 = ~a2018;
assign na2024 = ~a2024;
assign na2030 = ~a2030;
assign na2036 = ~a2036;
assign na2042 = ~a2042;
assign na2048 = ~a2048;
assign na2054 = ~a2054;
assign na2060 = ~a2060;
assign na2066 = ~a2066;
assign na2072 = ~a2072;
assign na2078 = ~a2078;
assign na2086 = ~a2086;
assign na2092 = ~a2092;
assign na2098 = ~a2098;
assign na2106 = ~a2106;
assign na2112 = ~a2112;
assign na2118 = ~a2118;
assign na2138 = ~a2138;
assign na2144 = ~a2144;
assign na2402 = ~a2402;
assign na2418 = ~a2418;
assign na2718 = ~a2718;
assign na2724 = ~a2724;
assign na2750 = ~a2750;
assign na2754 = ~a2754;
assign na2758 = ~a2758;
assign na2762 = ~a2762;
assign na2766 = ~a2766;
assign na2772 = ~a2772;
assign na2778 = ~a2778;
assign na2784 = ~a2784;
assign na2790 = ~a2790;
assign na2796 = ~a2796;
assign na2802 = ~a2802;
assign na2808 = ~a2808;
assign na2814 = ~a2814;
assign na2820 = ~a2820;
assign na2824 = ~a2824;
assign na2830 = ~a2830;
assign na2836 = ~a2836;
assign na2842 = ~a2842;
assign na2848 = ~a2848;
assign na2854 = ~a2854;
assign na2858 = ~a2858;
assign na2864 = ~a2864;
assign na2868 = ~a2868;
assign na2876 = ~a2876;
assign na2884 = ~a2884;
assign na2892 = ~a2892;
assign na2900 = ~a2900;
assign na2906 = ~a2906;
assign na2912 = ~a2912;
assign na2918 = ~a2918;
assign na2924 = ~a2924;
assign na2190 = ~a2190;
assign na2958 = ~a2958;
assign na2316 = ~a2316;
assign na2970 = ~a2970;
assign na2976 = ~a2976;
assign na2986 = ~a2986;
assign na2998 = ~a2998;
assign a4188 = a4186 & a3888;
assign c1 = 1;
assign na4194 = ~a4194;
assign a4374 = a4372 & a4292;
assign a4510 = a4508 & a4398;
assign a4586 = a4584 & a4552;
assign a4672 = a4670 & a4612;
assign a4708 = a4706 & a4360;
assign a4784 = a4782 & a4722;
assign a4830 = a4828 & a4804;
assign a4866 = a4864 & a4836;
assign na4872 = ~a4872;
assign na4884 = ~a4884;
assign na4890 = ~a4890;
assign na4902 = ~a4902;
assign na4914 = ~a4914;
assign na4926 = ~a4926;
assign na4938 = ~a4938;
assign na4950 = ~a4950;
assign na4962 = ~a4962;
assign a4964 = a4956 & ~a1942;
assign a4986 = a4984 & a4982;
assign a4992 = a4990 & a4046;
assign a5304 = a5302 & a5172;
assign a5336 = a5334 & a5330;
assign a5366 = a5364 & a5356;
assign a5368 = ~a1942 & a664;
assign a5376 = a5374 & a5078;
assign na5392 = ~a5392;
assign na5416 = ~a5416;
assign a5418 = ~a1942 & a608;
assign a5422 = ~a5420 & a5172;
assign a5428 = a5426 & a5362;
assign a5432 = ~a5430 & a5356;
assign a5458 = ~a5456 & ~a5442;
assign a5486 = a5484 & ~a5464;
assign na5494 = ~a5494;
assign a392 = l136 & i2;
assign a394 = ~l388 & l320;
assign a396 = ~l320 & i128;
assign a398 = ~a396 & ~a394;
assign a400 = ~a398 & ~l386;
assign a402 = a400 & ~a392;
assign a404 = a402 & ~l390;
assign a406 = l176 & i28;
assign a408 = l314 & i72;
assign a410 = ~a408 & ~a392;
assign a412 = a410 & a406;
assign a414 = ~a410 & i70;
assign a416 = a414 & l138;
assign a418 = ~a416 & ~a412;
assign a420 = ~a392 & l138;
assign a422 = ~a420 & l140;
assign a424 = ~l148 & ~l146;
assign a426 = a424 & ~l144;
assign a428 = a426 & l142;
assign a430 = ~l148 & l146;
assign a432 = a430 & ~l144;
assign a434 = a432 & i4;
assign a436 = ~a434 & ~a428;
assign a438 = a430 & l144;
assign a440 = a438 & i6;
assign a442 = a424 & l144;
assign a444 = a442 & i8;
assign a446 = ~a444 & ~a440;
assign a448 = a446 & a436;
assign a450 = a448 & ~l150;
assign a452 = a426 & l152;
assign a454 = a432 & i10;
assign a456 = ~a454 & ~a452;
assign a458 = a438 & i12;
assign a460 = a442 & i14;
assign a462 = ~a460 & ~a458;
assign a464 = a462 & a456;
assign a466 = ~a464 & l154;
assign a468 = ~a448 & l150;
assign a470 = ~a468 & ~a466;
assign a472 = ~a470 & ~a450;
assign a474 = ~a472 & l156;
assign a476 = a472 & ~l156;
assign a478 = ~a476 & ~a474;
assign a480 = a426 & l158;
assign a482 = a432 & l160;
assign a484 = ~a482 & ~a480;
assign a486 = a438 & l162;
assign a488 = a442 & l164;
assign a490 = ~a488 & ~a486;
assign a492 = a490 & a484;
assign a494 = ~a492 & a478;
assign a496 = a492 & ~a478;
assign a498 = ~a496 & ~a494;
assign a500 = ~a498 & a420;
assign a502 = ~a500 & ~a422;
assign a504 = ~l176 & ~l138;
assign a506 = ~a504 & ~a392;
assign a508 = ~l350 & ~l348;
assign a510 = a508 & ~l346;
assign a512 = a510 & l152;
assign a514 = a508 & l346;
assign a516 = a514 & i10;
assign a518 = ~a516 & ~a512;
assign a520 = ~l350 & l348;
assign a522 = a520 & ~l346;
assign a524 = a522 & i14;
assign a526 = a520 & l346;
assign a528 = a526 & i12;
assign a530 = ~a528 & ~a524;
assign a532 = a530 & a518;
assign a534 = ~a532 & l354;
assign a536 = a510 & l142;
assign a538 = a514 & i4;
assign a540 = ~a538 & ~a536;
assign a542 = a522 & i8;
assign a544 = a526 & i6;
assign a546 = ~a544 & ~a542;
assign a548 = a546 & a540;
assign a550 = a548 & ~l352;
assign a552 = ~a548 & l352;
assign a554 = ~a552 & ~a550;
assign a556 = ~a554 & ~a534;
assign a558 = a554 & a534;
assign a560 = ~a558 & ~a556;
assign a562 = a560 & a506;
assign a564 = ~a506 & l142;
assign a566 = ~a564 & ~a562;
assign a568 = ~l384 & l320;
assign a570 = ~l320 & i126;
assign a572 = ~a570 & ~a568;
assign a574 = ~a572 & a506;
assign a576 = ~a506 & l144;
assign a578 = ~a576 & ~a574;
assign a580 = ~l382 & l320;
assign a582 = ~l320 & i124;
assign a584 = ~a582 & ~a580;
assign a586 = ~a584 & a506;
assign a588 = ~a506 & l146;
assign a590 = ~a588 & ~a586;
assign a592 = ~l380 & l320;
assign a594 = ~l320 & i122;
assign a596 = ~a594 & ~a592;
assign a598 = ~a596 & a506;
assign a600 = ~a506 & l148;
assign a602 = ~a600 & ~a598;
assign a604 = ~l378 & l320;
assign a606 = ~l320 & ~i120;
assign a608 = ~a606 & ~a604;
assign a610 = a608 & a506;
assign a612 = ~a506 & l150;
assign a614 = ~a612 & ~a610;
assign a616 = ~l172 & l152;
assign a618 = ~l172 & ~i14;
assign a620 = l172 & ~i12;
assign a622 = ~a620 & ~a618;
assign a624 = ~a622 & ~i118;
assign a626 = i118 & ~i10;
assign a628 = ~l374 & l172;
assign a630 = a628 & ~a626;
assign a632 = a630 & ~a624;
assign a634 = ~a632 & ~a616;
assign a636 = ~a634 & ~l376;
assign a638 = a634 & l376;
assign a640 = ~a638 & ~a636;
assign a642 = ~a640 & a506;
assign a644 = ~a506 & l152;
assign a646 = ~a644 & ~a642;
assign a648 = ~l372 & l320;
assign a650 = ~l320 & i116;
assign a652 = ~a650 & ~a648;
assign a654 = ~a652 & a506;
assign a656 = ~a506 & l154;
assign a658 = ~a656 & ~a654;
assign a660 = ~l370 & l320;
assign a662 = ~l320 & ~i114;
assign a664 = ~a662 & ~a660;
assign a666 = a664 & a506;
assign a668 = ~a506 & l156;
assign a670 = ~a668 & ~a666;
assign a672 = a510 & l158;
assign a674 = a514 & l160;
assign a676 = ~a674 & ~a672;
assign a678 = a522 & l164;
assign a680 = a526 & l162;
assign a682 = ~a680 & ~a678;
assign a684 = a682 & a676;
assign a686 = ~a552 & ~a534;
assign a688 = ~a686 & ~a550;
assign a690 = ~a688 & l356;
assign a692 = a688 & ~l356;
assign a694 = ~a692 & ~a690;
assign a696 = a694 & ~a684;
assign a698 = ~a694 & a684;
assign a700 = ~a698 & ~a696;
assign a702 = ~a700 & a506;
assign a704 = ~a506 & l158;
assign a706 = ~a704 & ~a702;
assign a708 = a506 & l344;
assign a710 = ~a506 & l160;
assign a712 = ~a710 & ~a708;
assign a714 = a506 & l342;
assign a716 = ~a506 & l162;
assign a718 = ~a716 & ~a714;
assign a720 = a506 & ~i96;
assign a722 = ~a506 & l164;
assign a724 = ~a722 & ~a720;
assign a726 = l202 & ~l200;
assign a728 = a726 & ~l196;
assign a730 = a728 & ~l220;
assign a732 = ~l218 & l198;
assign a734 = ~l186 & ~l184;
assign a736 = a734 & l192;
assign a738 = l212 & l210;
assign a740 = ~l226 & ~l214;
assign a742 = l208 & l206;
assign a744 = a742 & l204;
assign a746 = a744 & a740;
assign a748 = a746 & a738;
assign a750 = a748 & a736;
assign a752 = a750 & a732;
assign a754 = a752 & ~l216;
assign a756 = ~l224 & ~l222;
assign a758 = a756 & l190;
assign a760 = a758 & a754;
assign a762 = a760 & ~l178;
assign a764 = a762 & ~l188;
assign a766 = a764 & ~l194;
assign a768 = a766 & a730;
assign a770 = a768 & l182;
assign a772 = a752 & ~l188;
assign a774 = a772 & a726;
assign a776 = a774 & a758;
assign a778 = a776 & ~l220;
assign a780 = a778 & ~l196;
assign a782 = a780 & ~l194;
assign a784 = a782 & l216;
assign a786 = a784 & ~l180;
assign a788 = a756 & ~l226;
assign a790 = a732 & ~l180;
assign a792 = a790 & ~l216;
assign a794 = a726 & ~l182;
assign a796 = a794 & ~l228;
assign a798 = a796 & l192;
assign a800 = a738 & ~l214;
assign a802 = a744 & ~l196;
assign a804 = a802 & a800;
assign a806 = a804 & a798;
assign a808 = a806 & a792;
assign a810 = ~l220 & ~l194;
assign a812 = a810 & l190;
assign a814 = a812 & l186;
assign a816 = a814 & a808;
assign a818 = a816 & a788;
assign a820 = ~a818 & ~a786;
assign a822 = ~a820 & ~l178;
assign a824 = ~a822 & ~a770;
assign a826 = ~l206 & ~l204;
assign a828 = a726 & l182;
assign a830 = ~l188 & ~l186;
assign a832 = a830 & ~l184;
assign a834 = a832 & a788;
assign a836 = a834 & l208;
assign a838 = a836 & a800;
assign a840 = a838 & ~l178;
assign a842 = a840 & ~l216;
assign a844 = a842 & a828;
assign a846 = ~l220 & l196;
assign a848 = ~l198 & ~l192;
assign a850 = ~l218 & l180;
assign a852 = a850 & a848;
assign a854 = a852 & ~l194;
assign a856 = a854 & a846;
assign a858 = a856 & a844;
assign a860 = a858 & a826;
assign a862 = a818 & l178;
assign a864 = ~a862 & ~a860;
assign a866 = a754 & a726;
assign a868 = a866 & ~l182;
assign a870 = l194 & ~l180;
assign a872 = a870 & ~l190;
assign a874 = a872 & a868;
assign a876 = a874 & ~l188;
assign a878 = a876 & ~l228;
assign a880 = a878 & ~l196;
assign a882 = a880 & l224;
assign a884 = a808 & ~l190;
assign a886 = a884 & l194;
assign a888 = a886 & l226;
assign a890 = a886 & l186;
assign a892 = a792 & ~l190;
assign a894 = l194 & l192;
assign a896 = a894 & a800;
assign a898 = a802 & a726;
assign a900 = a898 & a896;
assign a902 = a900 & a892;
assign a904 = a902 & a788;
assign a906 = a904 & ~l186;
assign a908 = a906 & l188;
assign a910 = ~a908 & ~a890;
assign a912 = a910 & ~a888;
assign a914 = a912 & ~a882;
assign a916 = a738 & ~l194;
assign a918 = a916 & l230;
assign a920 = a918 & ~l208;
assign a922 = a920 & ~l206;
assign a924 = ~l214 & ~l204;
assign a926 = a924 & a922;
assign a928 = a872 & a774;
assign a930 = a928 & ~l196;
assign a932 = a930 & ~l216;
assign a934 = ~a932 & ~a926;
assign a936 = ~a934 & l182;
assign a938 = a930 & l216;
assign a940 = a938 & a756;
assign a942 = ~l216 & l180;
assign a944 = a746 & l218;
assign a946 = a944 & a942;
assign a948 = a946 & a756;
assign a950 = ~l198 & l178;
assign a952 = a730 & l192;
assign a954 = a952 & a950;
assign a956 = a954 & a948;
assign a958 = ~l228 & ~l194;
assign a960 = a738 & ~l182;
assign a962 = a960 & a958;
assign a964 = a962 & a956;
assign a966 = a964 & a830;
assign a968 = l196 & l178;
assign a970 = a968 & ~l228;
assign a972 = a970 & a788;
assign a974 = l206 & l204;
assign a976 = a974 & ~l216;
assign a978 = ~l214 & l208;
assign a980 = a978 & a976;
assign a982 = a980 & a960;
assign a984 = a982 & a854;
assign a986 = a984 & a726;
assign a988 = a986 & a972;
assign a990 = ~a988 & ~a966;
assign a992 = a990 & ~a940;
assign a994 = a992 & ~a936;
assign a996 = a994 & a914;
assign a998 = a996 & a864;
assign a1000 = a998 & a824;
assign a1002 = a926 & l216;
assign a1004 = a852 & a840;
assign a1006 = a1004 & ~l220;
assign a1008 = a1006 & a726;
assign a1010 = a1008 & l196;
assign a1012 = a1010 & ~l194;
assign a1014 = a1012 & a826;
assign a1016 = a1014 & l216;
assign a1018 = ~a1016 & ~a1002;
assign a1020 = a902 & l228;
assign a1022 = a1014 & ~l216;
assign a1024 = a1022 & ~l182;
assign a1026 = a922 & ~l182;
assign a1028 = a1026 & a924;
assign a1030 = ~a1028 & ~a1024;
assign a1032 = ~a1030 & l228;
assign a1034 = ~a1032 & ~a1020;
assign a1036 = a1034 & a1018;
assign a1038 = ~l228 & ~l216;
assign a1040 = a1038 & a1026;
assign a1042 = a1040 & a924;
assign a1044 = a868 & a756;
assign a1046 = a870 & ~l188;
assign a1048 = a1046 & a1044;
assign a1050 = ~a1048 & ~a1024;
assign a1052 = ~a1050 & ~l228;
assign a1054 = ~a1052 & ~a1042;
assign a1056 = a948 & a738;
assign a1058 = a1056 & a832;
assign a1060 = l194 & ~l178;
assign a1062 = a1060 & a1058;
assign a1064 = a1062 & ~l198;
assign a1066 = a1064 & a846;
assign a1068 = a1066 & ~l192;
assign a1070 = a1068 & a796;
assign a1072 = ~a1070 & a1054;
assign a1074 = l194 & l180;
assign a1076 = a1074 & l196;
assign a1078 = a1076 & a764;
assign a1080 = ~a1078 & ~a1068;
assign a1082 = ~a1080 & a828;
assign a1084 = ~l198 & l196;
assign a1086 = a894 & l190;
assign a1088 = a1086 & a844;
assign a1090 = a1088 & a974;
assign a1092 = a1090 & l218;
assign a1094 = a1092 & a1084;
assign a1096 = a1094 & ~l220;
assign a1098 = ~l202 & l200;
assign a1100 = l198 & ~l194;
assign a1102 = l218 & ~l180;
assign a1104 = a800 & l208;
assign a1106 = a1104 & a788;
assign a1108 = a736 & ~l188;
assign a1110 = a976 & l190;
assign a1112 = a1110 & a1108;
assign a1114 = a1112 & a1106;
assign a1116 = a1114 & a1102;
assign a1118 = a1116 & a1100;
assign a1120 = a1118 & a1098;
assign a1122 = a1120 & l178;
assign a1124 = a1122 & ~l228;
assign a1126 = a1124 & l182;
assign a1128 = ~a1126 & ~a1096;
assign a1130 = l196 & ~l180;
assign a1132 = a1098 & l182;
assign a1134 = a1132 & a1130;
assign a1136 = a1134 & a766;
assign a1138 = l212 & ~l204;
assign a1140 = a1038 & a836;
assign a1142 = a1140 & l214;
assign a1144 = a1142 & l190;
assign a1146 = ~l206 & l182;
assign a1148 = a1146 & a1144;
assign a1150 = a1148 & a1138;
assign a1152 = a1116 & ~l178;
assign a1154 = a1152 & a1084;
assign a1156 = a1132 & a810;
assign a1158 = a1156 & a1154;
assign a1160 = ~a1158 & ~a1150;
assign a1162 = a1160 & ~a1136;
assign a1164 = a1162 & a1128;
assign a1166 = a1164 & ~a1082;
assign a1168 = a1166 & a1072;
assign a1170 = a1168 & a1036;
assign a1172 = a1170 & a1000;
assign a1174 = a1104 & a974;
assign a1176 = a1174 & a726;
assign a1178 = ~l218 & ~l216;
assign a1180 = a1178 & a1176;
assign a1182 = a1180 & ~l198;
assign a1184 = a1182 & ~l196;
assign a1186 = a1184 & a1086;
assign a1188 = a1186 & a832;
assign a1190 = a1188 & l182;
assign a1192 = a1190 & l180;
assign a1194 = l192 & l190;
assign a1196 = a1194 & a728;
assign a1198 = a1196 & a1058;
assign a1200 = a1198 & a1100;
assign a1202 = a1200 & ~l220;
assign a1204 = a1202 & l182;
assign a1206 = l204 & l182;
assign a1208 = a1206 & a742;
assign a1210 = ~l198 & l190;
assign a1212 = a1210 & a896;
assign a1214 = a1212 & a1208;
assign a1216 = a1214 & a728;
assign a1218 = a942 & ~l228;
assign a1220 = a1218 & a1216;
assign a1222 = a1220 & l218;
assign a1224 = ~a1222 & ~a1204;
assign a1226 = a1224 & ~a1192;
assign a1228 = ~a1226 & l178;
assign a1230 = a762 & ~l182;
assign a1232 = a726 & l194;
assign a1234 = a1232 & l228;
assign a1236 = a1234 & a1230;
assign a1238 = a1236 & ~l180;
assign a1240 = a1238 & ~l188;
assign a1242 = a1240 & ~l196;
assign a1244 = ~a1242 & ~a1228;
assign a1246 = a880 & ~l224;
assign a1248 = a1246 & l222;
assign a1250 = a1202 & ~l228;
assign a1252 = a1250 & l182;
assign a1254 = a1252 & ~l178;
assign a1256 = a788 & ~l180;
assign a1258 = l182 & l178;
assign a1260 = a1258 & a1186;
assign a1262 = a1260 & a1256;
assign a1264 = a906 & l184;
assign a1266 = l220 & l178;
assign a1268 = a1266 & a1264;
assign a1270 = a830 & a788;
assign a1272 = l184 & l178;
assign a1274 = a1272 & a1270;
assign a1276 = a1274 & a884;
assign a1278 = a1276 & ~l220;
assign a1280 = l180 & ~l178;
assign a1282 = a1280 & a730;
assign a1284 = a1270 & a1214;
assign a1286 = a1284 & a1282;
assign a1288 = a1286 & a1038;
assign a1290 = ~a1288 & ~a1278;
assign a1292 = a1290 & ~a1268;
assign a1294 = a1292 & ~a1262;
assign a1296 = a1294 & ~a1254;
assign a1298 = a1296 & ~a1248;
assign a1300 = a1298 & a1244;
assign a1302 = a782 & ~l216;
assign a1304 = a1302 & l228;
assign a1306 = a1142 & ~l210;
assign a1308 = a1306 & l190;
assign a1310 = a1308 & ~l230;
assign a1312 = a1310 & a1146;
assign a1314 = l212 & l194;
assign a1316 = a1314 & a1312;
assign a1318 = ~l340 & ~l228;
assign a1320 = ~l196 & l194;
assign a1322 = a1320 & a976;
assign a1324 = a1322 & a1318;
assign a1326 = a1324 & a1008;
assign a1328 = a1148 & l204;
assign a1330 = a1328 & ~a1314;
assign a1332 = a1330 & ~l210;
assign a1334 = ~a1332 & ~a1326;
assign a1336 = a1334 & ~a1316;
assign a1338 = a1336 & ~a1304;
assign a1340 = a1188 & ~l228;
assign a1342 = a1340 & ~l178;
assign a1344 = a1342 & a788;
assign a1346 = ~l220 & ~l180;
assign a1348 = a1346 & l182;
assign a1350 = a1348 & a1344;
assign a1352 = l188 & ~l180;
assign a1354 = a1230 & a958;
assign a1356 = a1354 & a730;
assign a1358 = a1356 & a1352;
assign a1360 = a970 & a760;
assign a1362 = a1360 & ~l188;
assign a1364 = a1362 & a1074;
assign a1366 = a1364 & a726;
assign a1368 = a1366 & l182;
assign a1370 = ~a1368 & ~a1358;
assign a1372 = a1370 & ~a1350;
assign a1374 = a1372 & a1338;
assign a1376 = a1374 & a1300;
assign a1378 = a1376 & a1172;
assign a1380 = a768 & ~l228;
assign a1382 = ~a1380 & ~a1366;
assign a1384 = ~a1382 & ~l182;
assign a1386 = ~l210 & ~l194;
assign a1388 = a1142 & ~l182;
assign a1390 = a1388 & l190;
assign a1392 = a1390 & l212;
assign a1394 = a1392 & a1386;
assign a1396 = a1394 & ~l206;
assign a1398 = a1396 & l204;
assign a1400 = a1392 & l206;
assign a1402 = a1400 & ~l204;
assign a1404 = l206 & l182;
assign a1406 = a1138 & l210;
assign a1408 = a1406 & a1144;
assign a1410 = a1408 & a1404;
assign a1412 = l214 & l190;
assign a1414 = a1040 & l204;
assign a1416 = a1414 & a1412;
assign a1418 = ~a1416 & ~a1410;
assign a1420 = a1418 & ~a1402;
assign a1422 = ~l228 & ~l182;
assign a1424 = a1422 & ~l178;
assign a1426 = a1424 & a1264;
assign a1428 = a956 & a918;
assign a1430 = a1428 & l182;
assign a1432 = a1412 & ~l212;
assign a1434 = a1432 & ~l182;
assign a1436 = a1434 & ~l208;
assign a1438 = a1436 & l206;
assign a1440 = a1434 & ~l206;
assign a1442 = a1440 & ~l208;
assign a1444 = a1442 & ~l204;
assign a1446 = ~a1444 & ~a1438;
assign a1448 = a1440 & a834;
assign a1450 = a1448 & l204;
assign a1452 = l210 & ~l206;
assign a1454 = a1452 & a1432;
assign a1456 = a1454 & a1206;
assign a1458 = ~a1456 & ~a1450;
assign a1460 = a1458 & a1446;
assign a1462 = a1460 & ~a1430;
assign a1464 = a1462 & ~a1426;
assign a1466 = a1464 & a1420;
assign a1468 = a1466 & ~a1398;
assign a1470 = a1468 & ~a1384;
assign a1472 = l220 & l196;
assign a1474 = a1472 & a1240;
assign a1476 = a1090 & a790;
assign a1478 = a1476 & l220;
assign a1480 = a794 & l228;
assign a1482 = a1480 & l196;
assign a1484 = ~a1482 & ~a828;
assign a1486 = ~a1484 & l194;
assign a1488 = a1486 & a1346;
assign a1490 = a1488 & a764;
assign a1492 = a1108 & l198;
assign a1494 = a980 & a788;
assign a1496 = a1494 & a916;
assign a1498 = a1496 & l190;
assign a1500 = a1498 & a1422;
assign a1502 = a1500 & a1492;
assign a1504 = ~a968 & ~l218;
assign a1506 = ~a1504 & a1502;
assign a1508 = a1506 & ~l180;
assign a1510 = a1508 & a1098;
assign a1512 = ~a1510 & ~a1490;
assign a1514 = a1512 & ~a1478;
assign a1516 = a1514 & ~a1474;
assign a1518 = a1044 & a812;
assign a1520 = a1518 & ~l196;
assign a1522 = a1520 & ~l228;
assign a1524 = a1522 & ~l188;
assign a1526 = a1524 & l178;
assign a1528 = ~a1526 & a1516;
assign a1530 = a1528 & a1470;
assign a1532 = a786 & l178;
assign a1534 = a1098 & ~l194;
assign a1536 = a1534 & a1362;
assign a1538 = a1536 & ~l180;
assign a1540 = a1538 & l182;
assign a1542 = a1318 & a1184;
assign a1544 = a1542 & ~l192;
assign a1546 = a1544 & ~l220;
assign a1548 = a1546 & a834;
assign a1550 = ~l180 & l178;
assign a1552 = a1550 & ~l194;
assign a1554 = a1552 & a1548;
assign a1556 = ~a1554 & ~a1540;
assign a1558 = a1556 & ~a1532;
assign a1560 = a1522 & a1352;
assign a1562 = a1560 & l178;
assign a1564 = a1302 & a1258;
assign a1566 = l194 & ~l182;
assign a1568 = a1566 & a950;
assign a1570 = a1568 & a1198;
assign a1572 = a1570 & ~l228;
assign a1574 = a1046 & a866;
assign a1576 = a1574 & a758;
assign a1578 = a1576 & l182;
assign a1580 = a1578 & l178;
assign a1582 = ~a1580 & ~a1572;
assign a1584 = a1582 & ~a1564;
assign a1586 = a1584 & ~a1562;
assign a1588 = a1586 & a1558;
assign a1590 = a1120 & ~l178;
assign a1592 = a1590 & l182;
assign a1594 = a798 & l190;
assign a1596 = a1594 & a1064;
assign a1598 = ~a1596 & ~a1592;
assign a1600 = l212 & l204;
assign a1602 = a1600 & a1310;
assign a1604 = a1602 & ~l182;
assign a1606 = a1604 & l194;
assign a1608 = a1606 & ~l206;
assign a1610 = a1078 & a796;
assign a1612 = a1502 & a1282;
assign a1614 = a1390 & ~l206;
assign a1616 = a1614 & a1138;
assign a1618 = ~a1616 & ~a1612;
assign a1620 = a1422 & a1154;
assign a1622 = a1534 & ~l220;
assign a1624 = ~a1622 & ~a1232;
assign a1626 = ~a1624 & a1620;
assign a1628 = ~a1626 & a1618;
assign a1630 = a1628 & ~a1610;
assign a1632 = a1630 & ~a1608;
assign a1634 = a1354 & a1130;
assign a1636 = a1634 & ~l188;
assign a1638 = a1636 & a1098;
assign a1640 = a1344 & ~l182;
assign a1642 = ~a1640 & ~a1638;
assign a1644 = a1642 & a1632;
assign a1646 = a1644 & a1598;
assign a1648 = a1388 & ~l212;
assign a1650 = a1648 & a974;
assign a1652 = a1208 & l214;
assign a1654 = l230 & l194;
assign a1656 = a1654 & ~l210;
assign a1658 = ~a1656 & l212;
assign a1660 = ~a1658 & a1652;
assign a1662 = ~a1660 & ~a1650;
assign a1664 = a1600 & a1306;
assign a1666 = a1664 & a1654;
assign a1668 = a1666 & ~a1404;
assign a1670 = ~a1668 & a1662;
assign a1672 = ~a1340 & ~a1250;
assign a1674 = ~a1672 & l178;
assign a1676 = a1674 & ~l182;
assign a1678 = ~a1676 & a1670;
assign a1680 = a846 & l228;
assign a1682 = a1680 & a876;
assign a1684 = a1682 & a756;
assign a1686 = a756 & ~l216;
assign a1688 = l228 & l220;
assign a1690 = ~a1688 & ~l182;
assign a1692 = ~a1690 & l196;
assign a1694 = a1692 & a1686;
assign a1696 = a1694 & a928;
assign a1698 = ~a1696 & ~a1684;
assign a1700 = a1454 & ~l208;
assign a1702 = a1700 & l182;
assign a1704 = a1394 & a974;
assign a1706 = ~a1704 & ~a1702;
assign a1708 = a1706 & a1698;
assign a1710 = a1708 & a1678;
assign a1712 = a1710 & a1646;
assign a1714 = a1712 & a1588;
assign a1716 = a1714 & a1530;
assign a1718 = a1716 & a1378;
assign a1720 = ~a1718 & a506;
assign a1722 = ~a506 & l166;
assign a1724 = ~a1722 & ~a1720;
assign a1726 = a1588 & a1072;
assign a1728 = a1094 & l220;
assign a1730 = a1112 & ~l178;
assign a1732 = a1730 & a1104;
assign a1734 = ~a1102 & l220;
assign a1736 = a1734 & a1320;
assign a1738 = a1736 & a1732;
assign a1740 = a1738 & ~l198;
assign a1742 = a1740 & a828;
assign a1744 = ~a1742 & ~a1438;
assign a1746 = a1744 & ~a1326;
assign a1748 = a1746 & ~a1704;
assign a1750 = a1748 & ~a1728;
assign a1752 = a1750 & a996;
assign a1754 = a1752 & ~a1676;
assign a1756 = a1754 & a1034;
assign a1758 = a1756 & a1726;
assign a1760 = ~a1758 & a506;
assign a1762 = ~a506 & l168;
assign a1764 = ~a1762 & ~a1760;
assign a1766 = ~a1378 & a506;
assign a1768 = ~a506 & l170;
assign a1770 = ~a1768 & ~a1766;
assign a1772 = ~a1264 & ~a1246;
assign a1774 = a1520 & ~l188;
assign a1776 = a1774 & l228;
assign a1778 = a1776 & ~l180;
assign a1780 = ~a1778 & a1772;
assign a1782 = a1776 & l180;
assign a1784 = ~a1782 & ~a1564;
assign a1786 = a1784 & a1780;
assign a1788 = a1312 & l204;
assign a1790 = a1124 & ~l182;
assign a1792 = ~a1790 & ~a1788;
assign a1794 = a1428 & ~l228;
assign a1796 = a1794 & a832;
assign a1798 = a1386 & a1328;
assign a1800 = ~a1798 & ~a1796;
assign a1802 = a1800 & ~a1572;
assign a1804 = a1802 & a1792;
assign a1806 = a1804 & ~a1524;
assign a1808 = ~l212 & l204;
assign a1810 = a1808 & a1614;
assign a1812 = a1810 & ~l210;
assign a1814 = a1450 & l210;
assign a1816 = ~a1814 & ~a1396;
assign a1818 = a1816 & ~a1812;
assign a1820 = a1818 & ~a1538;
assign a1822 = a1328 & ~l212;
assign a1824 = ~a1822 & ~a1220;
assign a1826 = a1824 & ~a1204;
assign a1828 = a1590 & a1422;
assign a1830 = ~a1828 & ~a1190;
assign a1832 = a1830 & ~a1366;
assign a1834 = a1832 & a1826;
assign a1836 = a1834 & a1820;
assign a1838 = a1836 & a1806;
assign a1840 = a1838 & a1646;
assign a1842 = ~a1446 & ~l210;
assign a1844 = a1442 & l204;
assign a1846 = ~a1844 & ~a1842;
assign a1848 = a1846 & a1420;
assign a1850 = a1848 & ~a1240;
assign a1852 = a1850 & ~a1560;
assign a1854 = a1852 & ~a1532;
assign a1856 = a1854 & a1840;
assign a1858 = a1856 & a1786;
assign a1860 = a1858 & a1172;
assign a1862 = a1566 & a1280;
assign a1864 = ~a1862 & ~a1552;
assign a1866 = ~a1864 & a1548;
assign a1868 = a1326 & l182;
assign a1870 = ~a1868 & ~a1866;
assign a1872 = a1870 & ~a1728;
assign a1874 = a1436 & l210;
assign a1876 = ~a1874 & ~a1578;
assign a1878 = a1876 & a1872;
assign a1880 = a1878 & a1710;
assign a1882 = a1880 & a1860;
assign a1884 = ~a1882 & a506;
assign a1886 = ~a506 & l172;
assign a1888 = ~a1886 & ~a1884;
assign a1890 = l228 & l190;
assign a1892 = a1890 & l178;
assign a1894 = a1892 & a1048;
assign a1896 = ~a1894 & a824;
assign a1898 = a1128 & ~a1002;
assign a1900 = a1898 & a1896;
assign a1902 = a1900 & a1300;
assign a1904 = ~a1902 & a506;
assign a1906 = ~a506 & l174;
assign a1908 = ~a1906 & ~a1904;
assign a1910 = ~a392 & ~l232;
assign a1912 = l244 & i20;
assign a1914 = l246 & i22;
assign a1916 = l248 & i24;
assign a1918 = l250 & i26;
assign a1920 = ~a1918 & ~a1916;
assign a1922 = a1920 & ~a1914;
assign a1924 = a1922 & ~a1912;
assign a1926 = a1924 & l234;
assign a1928 = a1926 & a1910;
assign a1930 = a406 & a392;
assign a1932 = ~a1930 & ~a1928;
assign a1934 = a1910 & l234;
assign a1936 = a1934 & ~l236;
assign a1938 = a1936 & l284;
assign a1940 = a504 & ~l234;
assign a1942 = ~a1940 & ~a392;
assign a1944 = l240 & l138;
assign a1946 = ~a1944 & ~l236;
assign a1948 = a1946 & a1942;
assign a1950 = ~a1948 & l178;
assign a1952 = ~a1950 & ~a1938;
assign a1954 = a1936 & l266;
assign a1956 = ~a1948 & l180;
assign a1958 = ~a1956 & ~a1954;
assign a1960 = ~a1946 & a1942;
assign a1962 = ~a1700 & ~a1408;
assign a1964 = a1962 & a1872;
assign a1966 = a1964 & a1678;
assign a1968 = a1840 & a1168;
assign a1970 = a1968 & a1966;
assign a1972 = ~a1970 & a1960;
assign a1974 = ~a1942 & l182;
assign a1976 = ~a1974 & ~a1972;
assign a1978 = a1960 & a882;
assign a1980 = ~a1942 & l184;
assign a1982 = ~a1980 & ~a1978;
assign a1984 = ~a940 & ~a786;
assign a1986 = ~a1984 & a1960;
assign a1988 = ~a1942 & l186;
assign a1990 = ~a1988 & ~a1986;
assign a1992 = ~a890 & ~a818;
assign a1994 = a1992 & ~a1560;
assign a1996 = ~a1994 & a1960;
assign a1998 = ~a1942 & l188;
assign a2000 = ~a1998 & ~a1996;
assign a2002 = a1936 & l286;
assign a2004 = ~a1936 & l190;
assign a2006 = ~a2004 & ~a2002;
assign a2008 = a1936 & l270;
assign a2010 = ~a1948 & l192;
assign a2012 = ~a2010 & ~a2008;
assign a2014 = a1936 & l276;
assign a2016 = ~a1948 & l194;
assign a2018 = ~a2016 & ~a2014;
assign a2020 = a1936 & l274;
assign a2022 = ~a1948 & l196;
assign a2024 = ~a2022 & ~a2020;
assign a2026 = a1936 & l278;
assign a2028 = ~a1948 & l198;
assign a2030 = ~a2028 & ~a2026;
assign a2032 = a1936 & l280;
assign a2034 = ~a1948 & l200;
assign a2036 = ~a2034 & ~a2032;
assign a2038 = a1936 & l282;
assign a2040 = ~a1948 & l202;
assign a2042 = ~a2040 & ~a2038;
assign a2044 = a1936 & l262;
assign a2046 = ~a1948 & l204;
assign a2048 = ~a2046 & ~a2044;
assign a2050 = a1936 & l254;
assign a2052 = ~a1948 & l206;
assign a2054 = ~a2052 & ~a2050;
assign a2056 = a1936 & l256;
assign a2058 = ~a1948 & l208;
assign a2060 = ~a2058 & ~a2056;
assign a2062 = a1936 & l252;
assign a2064 = ~a1948 & l210;
assign a2066 = ~a2064 & ~a2062;
assign a2068 = a1936 & l258;
assign a2070 = ~a1948 & l212;
assign a2072 = ~a2070 & ~a2068;
assign a2074 = a1936 & l260;
assign a2076 = ~a1948 & l214;
assign a2078 = ~a2076 & ~a2074;
assign a2080 = ~a1778 & a1036;
assign a2082 = ~a2080 & a1960;
assign a2084 = ~a1942 & l216;
assign a2086 = ~a2084 & ~a2082;
assign a2088 = a1936 & l268;
assign a2090 = ~a1948 & l218;
assign a2092 = ~a2090 & ~a2088;
assign a2094 = a1936 & l272;
assign a2096 = ~a1948 & l220;
assign a2098 = ~a2096 & ~a2094;
assign a2100 = ~a1264 & ~a1248;
assign a2102 = ~a2100 & a1960;
assign a2104 = ~a1942 & l222;
assign a2106 = ~a2104 & ~a2102;
assign a2108 = a1960 & a888;
assign a2110 = ~a1942 & l224;
assign a2112 = ~a2110 & ~a2108;
assign a2114 = a1960 & a908;
assign a2116 = ~a1942 & l226;
assign a2118 = ~a2116 & ~a2114;
assign a2120 = ~a1240 & ~a936;
assign a2122 = ~a1578 & ~a860;
assign a2124 = a2122 & ~a1894;
assign a2126 = a2124 & a1698;
assign a2128 = a2126 & a2120;
assign a2130 = a2128 & ~a770;
assign a2132 = a2130 & a1784;
assign a2134 = ~a2132 & a1960;
assign a2136 = ~a1942 & l228;
assign a2138 = ~a2136 & ~a2134;
assign a2140 = a1936 & l238;
assign a2142 = ~a1948 & l230;
assign a2144 = ~a2142 & ~a2140;
assign a2146 = l242 & i16;
assign a2148 = a1910 & l290;
assign a2150 = a2148 & ~i24;
assign a2152 = a1910 & l288;
assign a2154 = a2152 & ~i26;
assign a2156 = ~a2154 & ~a2150;
assign a2158 = a1910 & l294;
assign a2160 = a2158 & ~i20;
assign a2162 = a1910 & l292;
assign a2164 = a2162 & ~i22;
assign a2166 = ~a2164 & ~a2160;
assign a2168 = a2166 & a2156;
assign a2170 = ~a2168 & a2146;
assign a2172 = l296 & ~i24;
assign a2174 = l298 & ~i26;
assign a2176 = ~a2174 & ~a2172;
assign a2178 = l300 & ~i20;
assign a2180 = l302 & ~i22;
assign a2182 = ~a2180 & ~a2178;
assign a2184 = a2182 & a2176;
assign a2186 = ~a2184 & ~a1910;
assign a2188 = a2186 & l304;
assign a2190 = ~a2188 & ~a2170;
assign a2192 = l264 & l262;
assign a2194 = a2192 & l260;
assign a2196 = a2194 & ~l258;
assign a2198 = a2196 & ~l256;
assign a2200 = a2198 & ~l254;
assign a2202 = a2200 & ~l252;
assign a2204 = l268 & l266;
assign a2206 = ~l274 & ~l272;
assign a2208 = ~l276 & l252;
assign a2210 = a2208 & l262;
assign a2212 = l282 & ~l280;
assign a2214 = a2212 & ~l278;
assign a2216 = l258 & l256;
assign a2218 = a2216 & l254;
assign a2220 = a2218 & l284;
assign a2222 = a2220 & a2214;
assign a2224 = a2222 & a2210;
assign a2226 = a2224 & ~l260;
assign a2228 = a2226 & a2206;
assign a2230 = a2228 & l270;
assign a2232 = a2230 & a2204;
assign a2234 = a2232 & ~l238;
assign a2236 = l264 & l260;
assign a2238 = a2236 & ~l262;
assign a2240 = a2238 & l254;
assign a2242 = a2240 & a2216;
assign a2244 = a2242 & ~l252;
assign a2246 = ~a2244 & ~a2234;
assign a2248 = a2246 & ~a2202;
assign a2250 = ~l270 & l266;
assign a2252 = a2250 & l274;
assign a2254 = a2252 & ~l268;
assign a2256 = a2254 & a2226;
assign a2258 = a2198 & l254;
assign a2260 = ~l256 & ~l254;
assign a2262 = l258 & l238;
assign a2264 = a2262 & a2236;
assign a2266 = a2264 & a2210;
assign a2268 = a2266 & a2260;
assign a2270 = ~l258 & ~l256;
assign a2272 = a2270 & a2240;
assign a2274 = a2272 & l252;
assign a2276 = l260 & ~l252;
assign a2278 = a2218 & a2192;
assign a2280 = a2278 & ~l276;
assign a2282 = a2280 & a2276;
assign a2284 = ~a2282 & ~a2274;
assign a2286 = a2284 & ~a2268;
assign a2288 = a2286 & ~a2258;
assign a2290 = a2288 & ~a2256;
assign a2292 = a2236 & ~l254;
assign a2294 = a2292 & ~l262;
assign a2296 = a2294 & a2270;
assign a2298 = a2296 & ~l252;
assign a2300 = a2272 & ~l252;
assign a2302 = ~a2300 & ~a2298;
assign a2304 = a2302 & a2290;
assign a2306 = a2304 & a2248;
assign a2308 = a2306 & a1934;
assign a2310 = ~a2308 & ~l306;
assign a2312 = ~a2310 & ~a392;
assign a2314 = a392 & l308;
assign a2316 = ~a2314 & ~a2312;
assign a2318 = ~a2316 & ~a2190;
assign a2320 = l290 & ~i24;
assign a2322 = l292 & ~i22;
assign a2324 = a2158 & i20;
assign a2326 = a2162 & ~l294;
assign a2328 = ~a2326 & ~a2324;
assign a2330 = ~a2328 & ~a2322;
assign a2332 = a1910 & ~l292;
assign a2334 = a2332 & ~l294;
assign a2336 = a2334 & l290;
assign a2338 = ~a2336 & ~a2330;
assign a2340 = ~a2338 & ~a2320;
assign a2342 = l288 & ~i26;
assign a2344 = a2342 & a2340;
assign a2346 = l288 & i26;
assign a2348 = l290 & i24;
assign a2350 = l292 & i22;
assign a2352 = ~a2326 & ~a2160;
assign a2354 = ~a2352 & ~a2350;
assign a2356 = ~a2354 & ~a2336;
assign a2358 = ~a2356 & ~a2348;
assign a2360 = a2358 & a2346;
assign a2362 = ~a2360 & ~a2344;
assign a2364 = a2354 & a2348;
assign a2366 = a2330 & a2320;
assign a2368 = a2324 & a2322;
assign a2370 = a2350 & a2160;
assign a2372 = ~a2370 & ~a2368;
assign a2374 = a2372 & ~a2366;
assign a2376 = a2374 & ~a2364;
assign a2378 = a2376 & a2362;
assign a2380 = l242 & ~i16;
assign a2382 = a2380 & ~a2378;
assign a2384 = a2382 & a1942;
assign a2386 = a2334 & ~l290;
assign a2388 = a2386 & l288;
assign a2390 = ~a2388 & ~a2358;
assign a2392 = ~a2390 & ~a2346;
assign a2394 = a2392 & a2380;
assign a2396 = a2394 & a1942;
assign a2398 = ~a2396 & ~i68;
assign a2400 = a2398 & ~a2384;
assign a2402 = a2400 & ~a2318;
assign a2404 = a2146 & a1910;
assign a2406 = l294 & i20;
assign a2408 = ~a2348 & ~a2346;
assign a2410 = a2408 & ~a2350;
assign a2412 = a2410 & ~a2406;
assign a2414 = a2412 & a2404;
assign a2416 = a1926 & ~a1910;
assign a2418 = ~a2416 & ~a2414;
assign a2420 = a2308 & a1924;
assign a2422 = l274 & ~l266;
assign a2424 = ~l260 & l252;
assign a2426 = a2424 & l270;
assign a2428 = a2426 & a2278;
assign a2430 = a2428 & ~l284;
assign a2432 = ~l282 & l280;
assign a2434 = a2432 & a2430;
assign a2436 = a2434 & a2422;
assign a2438 = a2436 & ~l276;
assign a2440 = a2438 & l278;
assign a2442 = a2440 & l268;
assign a2444 = a2212 & l276;
assign a2446 = a2444 & a2430;
assign a2448 = l278 & ~l268;
assign a2450 = a2448 & a2446;
assign a2452 = a2450 & l274;
assign a2454 = a2452 & ~l272;
assign a2456 = a2454 & l266;
assign a2458 = a2438 & ~l272;
assign a2460 = a2458 & a2448;
assign a2462 = ~a2460 & ~a2456;
assign a2464 = a2462 & ~a2442;
assign a2466 = a2430 & ~l274;
assign a2468 = a2466 & a2444;
assign a2470 = ~l268 & ~l266;
assign a2472 = a2470 & a2468;
assign a2474 = a2472 & l278;
assign a2476 = ~l272 & l268;
assign a2478 = l278 & ~l276;
assign a2480 = a2478 & a2476;
assign a2482 = a2480 & a2466;
assign a2484 = a2482 & l266;
assign a2486 = a2484 & a2212;
assign a2488 = l272 & ~l266;
assign a2490 = a2488 & a2450;
assign a2492 = ~a2490 & ~a2486;
assign a2494 = a2492 & ~a2474;
assign a2496 = a2454 & ~l266;
assign a2498 = a2428 & ~l274;
assign a2500 = a2498 & a2478;
assign a2502 = a2500 & ~l272;
assign a2504 = a2502 & a2212;
assign a2506 = a2504 & ~l268;
assign a2508 = a2498 & a2444;
assign a2510 = a2508 & ~l268;
assign a2512 = ~l278 & l266;
assign a2514 = a2512 & a2510;
assign a2516 = a2514 & l284;
assign a2518 = ~a2516 & ~a2506;
assign a2520 = a2518 & ~a2496;
assign a2522 = a2520 & a2494;
assign a2524 = a2292 & a2216;
assign a2526 = a2524 & l252;
assign a2528 = a2526 & ~l262;
assign a2530 = a2472 & ~l278;
assign a2532 = a2530 & ~l272;
assign a2534 = l272 & l266;
assign a2536 = a2534 & a2452;
assign a2538 = ~a2536 & ~a2532;
assign a2540 = a2538 & ~a2528;
assign a2542 = ~l278 & l268;
assign a2544 = a2542 & a2446;
assign a2546 = a2544 & a2534;
assign a2548 = a2524 & ~l252;
assign a2550 = a2548 & ~l276;
assign a2552 = ~a2550 & ~a2546;
assign a2554 = a2548 & ~l262;
assign a2556 = a2544 & a2422;
assign a2558 = a2556 & l272;
assign a2560 = a2200 & l252;
assign a2562 = ~a2560 & ~a2558;
assign a2564 = a2530 & l272;
assign a2566 = ~a2564 & a2562;
assign a2568 = a2566 & ~a2554;
assign a2570 = a2568 & a2552;
assign a2572 = a2570 & ~a2274;
assign a2574 = a2572 & a2540;
assign a2576 = a2574 & a2522;
assign a2578 = a2576 & a2464;
assign a2580 = a2196 & l256;
assign a2582 = a2580 & ~l254;
assign a2584 = ~a2582 & ~a2282;
assign a2586 = l284 & l266;
assign a2588 = a2586 & l268;
assign a2590 = a2588 & a2504;
assign a2592 = a2432 & l268;
assign a2594 = a2592 & a2488;
assign a2596 = a2594 & a2500;
assign a2598 = ~a2596 & ~a2590;
assign a2600 = a2242 & l252;
assign a2602 = a2432 & l270;
assign a2604 = a2424 & a2280;
assign a2606 = l278 & ~l266;
assign a2608 = a2606 & a2604;
assign a2610 = a2608 & a2602;
assign a2612 = a2610 & l284;
assign a2614 = a2612 & l274;
assign a2616 = a2614 & ~l268;
assign a2618 = ~a2616 & ~a2600;
assign a2620 = a2618 & ~a2244;
assign a2622 = a2620 & a2598;
assign a2624 = a2512 & a2468;
assign a2626 = ~a2624 & ~a2258;
assign a2628 = a2626 & a2622;
assign a2630 = a2628 & a2584;
assign a2632 = a2544 & ~l272;
assign a2634 = a2632 & l274;
assign a2636 = ~a2634 & ~a2268;
assign a2638 = l274 & l272;
assign a2640 = a2638 & a2610;
assign a2642 = l256 & ~l252;
assign a2644 = a2642 & a2194;
assign a2646 = a2644 & ~l254;
assign a2648 = a2646 & l258;
assign a2650 = a2648 & ~l238;
assign a2652 = ~a2650 & ~a2640;
assign a2654 = a2652 & ~a2300;
assign a2656 = a2654 & ~a2296;
assign a2658 = a2586 & a2508;
assign a2660 = a2658 & ~l278;
assign a2662 = a2660 & l268;
assign a2664 = a2444 & a2428;
assign a2666 = a2664 & a2448;
assign a2668 = a2666 & l284;
assign a2670 = a2668 & ~l266;
assign a2672 = ~a2670 & ~a2662;
assign a2674 = a2510 & l284;
assign a2676 = a2674 & ~l266;
assign a2678 = a2668 & l274;
assign a2680 = a2678 & l266;
assign a2682 = ~a2680 & ~a2676;
assign a2684 = a2542 & a2458;
assign a2686 = a2612 & l268;
assign a2688 = a2482 & a2432;
assign a2690 = a2688 & ~l266;
assign a2692 = ~a2690 & ~a2686;
assign a2694 = a2692 & ~a2684;
assign a2696 = a2694 & a2682;
assign a2698 = a2696 & a2672;
assign a2700 = ~a2202 & l286;
assign a2702 = a2700 & a2698;
assign a2704 = a2702 & a2656;
assign a2706 = a2704 & a2636;
assign a2708 = a2706 & a2630;
assign a2710 = a2708 & a2578;
assign a2712 = ~a2710 & a2420;
assign a2714 = l236 & i28;
assign a2716 = a2714 & a392;
assign a2718 = ~a2716 & ~a2712;
assign a2720 = a2404 & i18;
assign a2722 = ~a2404 & l238;
assign a2724 = ~a2722 & ~a2720;
assign a2726 = a2128 & a1984;
assign a2728 = a2726 & a1780;
assign a2730 = a780 & ~l180;
assign a2732 = a2730 & a1038;
assign a2734 = a1670 & ~a1020;
assign a2736 = a2734 & ~a2732;
assign a2738 = a2736 & ~a1524;
assign a2740 = a2738 & a914;
assign a2742 = a2740 & a1054;
assign a2744 = a2742 & a2728;
assign a2746 = ~a2744 & a506;
assign a2748 = ~a506 & l240;
assign a2750 = ~a2748 & ~a2746;
assign a2752 = ~a1910 & l244;
assign a2754 = ~a2752 & ~a2158;
assign a2756 = ~a1910 & l246;
assign a2758 = ~a2756 & ~a2162;
assign a2760 = ~a1910 & l248;
assign a2762 = ~a2760 & ~a2148;
assign a2764 = ~a1910 & l250;
assign a2766 = ~a2764 & ~a2152;
assign a2768 = a2404 & i62;
assign a2770 = ~a2404 & l252;
assign a2772 = ~a2770 & ~a2768;
assign a2774 = a2404 & i60;
assign a2776 = ~a2404 & l254;
assign a2778 = ~a2776 & ~a2774;
assign a2780 = a2404 & i58;
assign a2782 = ~a2404 & l256;
assign a2784 = ~a2782 & ~a2780;
assign a2786 = a2404 & i56;
assign a2788 = ~a2404 & l258;
assign a2790 = ~a2788 & ~a2786;
assign a2792 = a2404 & i54;
assign a2794 = ~a2404 & l260;
assign a2796 = ~a2794 & ~a2792;
assign a2798 = a2404 & i52;
assign a2800 = ~a2404 & l262;
assign a2802 = ~a2800 & ~a2798;
assign a2804 = a2404 & ~i30;
assign a2806 = ~a2404 & l264;
assign a2808 = ~a2806 & ~a2804;
assign a2810 = a2404 & i50;
assign a2812 = ~a2404 & l266;
assign a2814 = ~a2812 & ~a2810;
assign a2816 = a2404 & i48;
assign a2818 = ~a2404 & l268;
assign a2820 = ~a2818 & ~a2816;
assign a2822 = ~a2404 & l270;
assign a2824 = ~a2822 & ~i46;
assign a2826 = a2404 & i44;
assign a2828 = ~a2404 & l272;
assign a2830 = ~a2828 & ~a2826;
assign a2832 = a2404 & i42;
assign a2834 = ~a2404 & l274;
assign a2836 = ~a2834 & ~a2832;
assign a2838 = a2404 & i40;
assign a2840 = ~a2404 & l276;
assign a2842 = ~a2840 & ~a2838;
assign a2844 = a2404 & i38;
assign a2846 = ~a2404 & l278;
assign a2848 = ~a2846 & ~a2844;
assign a2850 = a2404 & i36;
assign a2852 = ~a2404 & l280;
assign a2854 = ~a2852 & ~a2850;
assign a2856 = ~a2404 & l282;
assign a2858 = ~a2856 & ~i34;
assign a2860 = a2404 & i32;
assign a2862 = ~a2404 & l284;
assign a2864 = ~a2862 & ~a2860;
assign a2866 = ~a1910 & l286;
assign a2868 = ~a2866 & ~a2804;
assign a2870 = i66 & i64;
assign a2872 = a2870 & a1910;
assign a2874 = ~a1910 & l288;
assign a2876 = ~a2874 & ~a2872;
assign a2878 = i66 & ~i64;
assign a2880 = a2878 & a1910;
assign a2882 = ~a1910 & l290;
assign a2884 = ~a2882 & ~a2880;
assign a2886 = ~i66 & i64;
assign a2888 = a2886 & a1910;
assign a2890 = ~a1910 & l292;
assign a2892 = ~a2890 & ~a2888;
assign a2894 = ~i66 & ~i64;
assign a2896 = a2894 & a1910;
assign a2898 = ~a1910 & l294;
assign a2900 = ~a2898 & ~a2896;
assign a2902 = ~a2168 & l290;
assign a2904 = a2186 & l296;
assign a2906 = ~a2904 & ~a2902;
assign a2908 = ~a2168 & l288;
assign a2910 = a2186 & l298;
assign a2912 = ~a2910 & ~a2908;
assign a2914 = ~a2168 & l294;
assign a2916 = a2186 & l300;
assign a2918 = ~a2916 & ~a2914;
assign a2920 = ~a2168 & l292;
assign a2922 = a2186 & l302;
assign a2924 = ~a2922 & ~a2920;
assign a2926 = ~a1924 & l234;
assign a2928 = a2926 & a504;
assign a2930 = l138 & ~i70;
assign a2932 = ~a2930 & ~l176;
assign a2934 = ~a2932 & ~a406;
assign a2936 = a2934 & ~l234;
assign a2938 = ~a2936 & ~a2928;
assign a2940 = a2938 & a392;
assign a2942 = a2940 & l306;
assign a2944 = l310 & l138;
assign a2946 = a2944 & ~l312;
assign a2948 = a2946 & i70;
assign a2950 = a2948 & i72;
assign a2952 = ~a2950 & ~a2714;
assign a2954 = a2952 & ~a2420;
assign a2956 = ~a2954 & ~a392;
assign a2958 = ~a2956 & ~a2942;
assign a2960 = l320 & ~l318;
assign a2962 = ~l320 & i76;
assign a2964 = ~a2962 & ~a2960;
assign a2966 = ~a2964 & a506;
assign a2968 = ~a506 & l310;
assign a2970 = ~a2968 & ~a2966;
assign a2972 = a412 & l316;
assign a2974 = a414 & l312;
assign a2976 = ~a2974 & ~a2972;
assign a2978 = a2940 & l314;
assign a2980 = a2948 & i74;
assign a2982 = ~a2980 & ~a2714;
assign a2984 = ~a2982 & ~a392;
assign a2986 = ~a2984 & ~a2978;
assign a2988 = ~l234 & ~l176;
assign a2990 = ~a2988 & ~a392;
assign a2992 = a2990 & l234;
assign a2994 = a2992 & a2710;
assign a2996 = ~a2990 & l316;
assign a2998 = ~a2996 & ~a2994;
assign a3000 = a2470 & a2228;
assign a3002 = a3000 & ~l322;
assign a3004 = a3002 & ~l270;
assign a3006 = a2424 & a2216;
assign a3008 = a3006 & ~l284;
assign a3010 = a3008 & a2212;
assign a3012 = l276 & l262;
assign a3014 = a3012 & l254;
assign a3016 = a3014 & a3010;
assign a3018 = a3016 & ~l268;
assign a3020 = a3018 & ~l274;
assign a3022 = ~l278 & ~l272;
assign a3024 = a3022 & a2250;
assign a3026 = a3024 & a3020;
assign a3028 = a3026 & ~l322;
assign a3030 = a3012 & a2216;
assign a3032 = a3030 & l238;
assign a3034 = a3032 & a2276;
assign a3036 = a3034 & ~l254;
assign a3038 = ~a3036 & ~a3028;
assign a3040 = a3038 & ~a3004;
assign a3042 = ~a2582 & ~a2202;
assign a3044 = a3042 & a2540;
assign a3046 = ~a2442 & ~a2256;
assign a3048 = a2636 & ~a2232;
assign a3050 = a3048 & a3046;
assign a3052 = a3050 & a2462;
assign a3054 = a3052 & ~a2686;
assign a3056 = a3054 & a3044;
assign a3058 = a2672 & a2494;
assign a3060 = ~l268 & l254;
assign a3062 = a3060 & a3030;
assign a3064 = a3062 & a2426;
assign a3066 = a3064 & a2606;
assign a3068 = a3066 & ~l264;
assign a3070 = a3068 & a2212;
assign a3072 = a3070 & l284;
assign a3074 = a3072 & l272;
assign a3076 = a2440 & l272;
assign a3078 = ~a3076 & ~a3074;
assign a3080 = a3072 & ~l272;
assign a3082 = a3080 & ~l274;
assign a3084 = a2296 & l252;
assign a3086 = ~a3084 & ~a3082;
assign a3088 = a2646 & l276;
assign a3090 = a2632 & l266;
assign a3092 = a2506 & ~l284;
assign a3094 = a3080 & l274;
assign a3096 = ~a3094 & ~a3092;
assign a3098 = a3096 & ~a3090;
assign a3100 = a3098 & ~a3088;
assign a3102 = a3100 & a3086;
assign a3104 = a3102 & a3078;
assign a3106 = a3104 & a3058;
assign a3108 = a3106 & a3056;
assign a3110 = a3108 & a3040;
assign a3112 = ~a3110 & a1936;
assign a3114 = ~a2944 & ~l236;
assign a3116 = ~l324 & l320;
assign a3118 = ~l320 & i78;
assign a3120 = ~a3118 & ~a3116;
assign a3122 = ~a3120 & ~a3114;
assign a3124 = ~a3122 & ~a3112;
assign a3126 = ~a3076 & ~a3004;
assign a3128 = a3126 & ~a2474;
assign a3130 = a3070 & ~l284;
assign a3132 = a3130 & ~l272;
assign a3134 = a3132 & l274;
assign a3136 = a2670 & l272;
assign a3138 = ~a3136 & ~a3134;
assign a3140 = a3138 & ~a3082;
assign a3142 = ~a2564 & ~a2496;
assign a3144 = a2642 & a2264;
assign a3146 = l262 & ~l254;
assign a3148 = a3146 & a3144;
assign a3150 = ~a3148 & ~a3092;
assign a3152 = a3150 & ~a2298;
assign a3154 = a3152 & a3142;
assign a3156 = l272 & l270;
assign a3158 = a3156 & a3020;
assign a3160 = a3158 & a2606;
assign a3162 = ~a3160 & ~a3028;
assign a3164 = a3162 & ~a3036;
assign a3166 = a2514 & l272;
assign a3168 = a2670 & l274;
assign a3170 = a2686 & ~l274;
assign a3172 = ~l262 & ~l254;
assign a3174 = a3022 & a2254;
assign a3176 = a3174 & a3010;
assign a3178 = a3176 & ~l276;
assign a3180 = a3178 & a3172;
assign a3182 = ~a3180 & ~a2556;
assign a3184 = a3182 & ~a2536;
assign a3186 = a3184 & ~a3170;
assign a3188 = a3186 & ~a3168;
assign a3190 = a3188 & ~a3166;
assign a3192 = a3190 & a3164;
assign a3194 = a3192 & a3154;
assign a3196 = a3194 & a2630;
assign a3198 = a3196 & a3046;
assign a3200 = a3198 & a3140;
assign a3202 = a3200 & a3128;
assign a3204 = ~a3202 & a1936;
assign a3206 = ~l326 & l320;
assign a3208 = ~l320 & i80;
assign a3210 = ~a3208 & ~a3206;
assign a3212 = ~a3210 & ~a3114;
assign a3214 = ~a3212 & ~a3204;
assign a3216 = a3034 & l254;
assign a3218 = ~a3216 & ~a2490;
assign a3220 = a2624 & ~l268;
assign a3222 = ~a3220 & ~a2590;
assign a3224 = a3222 & ~a2272;
assign a3226 = a3224 & a3040;
assign a3228 = a2262 & a2208;
assign a3230 = ~l262 & ~l260;
assign a3232 = a3230 & a3228;
assign a3234 = a3232 & a2260;
assign a3236 = ~a3234 & ~a3180;
assign a3238 = a2506 & ~l266;
assign a3240 = l254 & l252;
assign a3242 = a3240 & a2196;
assign a3244 = a3130 & a2638;
assign a3246 = a3074 & ~l274;
assign a3248 = ~a3246 & ~a3244;
assign a3250 = a3248 & ~a3242;
assign a3252 = a3250 & ~a3238;
assign a3254 = a3252 & a3236;
assign a3256 = a3144 & l254;
assign a3258 = a2256 & l272;
assign a3260 = l262 & l260;
assign a3262 = a3260 & ~l258;
assign a3264 = l256 & l254;
assign a3266 = a3264 & a3262;
assign a3268 = a2476 & ~l278;
assign a3270 = a3016 & a2252;
assign a3272 = a3270 & a3268;
assign a3274 = ~a3272 & ~a3266;
assign a3276 = a3274 & ~a3258;
assign a3278 = a3276 & ~a3256;
assign a3280 = a3278 & a3086;
assign a3282 = a3280 & a3254;
assign a3284 = a3282 & a2248;
assign a3286 = a3284 & a3226;
assign a3288 = a3286 & a3138;
assign a3290 = a3288 & a3218;
assign a3292 = ~a3290 & a1936;
assign a3294 = ~l328 & l320;
assign a3296 = ~l320 & i82;
assign a3298 = ~a3296 & ~a3294;
assign a3300 = ~a3298 & ~a3114;
assign a3302 = ~a3300 & ~a3292;
assign a3304 = a2522 & ~a2232;
assign a3306 = a3304 & a2698;
assign a3308 = a3306 & a2622;
assign a3310 = a3308 & a2290;
assign a3312 = ~a3310 & a1936;
assign a3314 = ~l330 & l320;
assign a3316 = ~l320 & i84;
assign a3318 = ~a3316 & ~a3314;
assign a3320 = ~a3318 & ~a3114;
assign a3322 = ~a3320 & ~a3312;
assign a3324 = ~a3244 & ~a3004;
assign a3326 = a3324 & ~a3216;
assign a3328 = a3326 & a3078;
assign a3330 = a3328 & a2578;
assign a3332 = a3330 & a3162;
assign a3334 = ~a3332 & a1936;
assign a3336 = ~l332 & l320;
assign a3338 = ~l320 & i86;
assign a3340 = ~a3338 & ~a3336;
assign a3342 = ~a3340 & ~a3114;
assign a3344 = ~a3342 & ~a3334;
assign a3346 = ~a2680 & a2618;
assign a3348 = ~a3272 & ~a2244;
assign a3350 = ~a2624 & a2570;
assign a3352 = a3350 & a2656;
assign a3354 = a3352 & a3056;
assign a3356 = a3354 & a3236;
assign a3358 = a3356 & a3348;
assign a3360 = a3358 & a3346;
assign a3362 = ~a3360 & a1936;
assign a3364 = ~l334 & l320;
assign a3366 = ~l320 & i88;
assign a3368 = ~a3366 & ~a3364;
assign a3370 = ~a3368 & ~a3114;
assign a3372 = ~a3370 & ~a3362;
assign a3374 = ~a2554 & ~a2516;
assign a3376 = ~a2616 & ~a2258;
assign a3378 = a3376 & a3154;
assign a3380 = a3132 & ~l274;
assign a3382 = a2582 & l252;
assign a3384 = ~a2650 & ~a2486;
assign a3386 = a3384 & ~a3382;
assign a3388 = a3386 & ~a3380;
assign a3390 = a3388 & a2682;
assign a3392 = a3390 & a3052;
assign a3394 = a3392 & a3226;
assign a3396 = a3394 & a3378;
assign a3398 = a3396 & a3374;
assign a3400 = ~a3398 & a1936;
assign a3402 = ~l336 & l320;
assign a3404 = ~l320 & i90;
assign a3406 = ~a3404 & ~a3402;
assign a3408 = ~a3406 & ~a3114;
assign a3410 = ~a3408 & ~a3400;
assign a3412 = ~a2690 & ~a2496;
assign a3414 = a2654 & a2566;
assign a3416 = ~a2528 & ~a2486;
assign a3418 = a3254 & ~a2202;
assign a3420 = a3164 & ~a2600;
assign a3422 = a3420 & a2584;
assign a3424 = a2660 & ~l272;
assign a3426 = a3266 & l252;
assign a3428 = ~a2686 & ~a2678;
assign a3430 = ~a3428 & l272;
assign a3432 = a2232 & l238;
assign a3434 = ~a3432 & ~a3094;
assign a3436 = a3434 & ~a2460;
assign a3438 = a3436 & ~a3430;
assign a3440 = ~a2676 & ~a2514;
assign a3442 = ~a3440 & ~l272;
assign a3444 = ~a3442 & a3438;
assign a3446 = a3444 & ~a3426;
assign a3448 = a3446 & ~a3424;
assign a3450 = a3448 & a3422;
assign a3452 = a3450 & a3418;
assign a3454 = a3452 & a3416;
assign a3456 = a3454 & a3414;
assign a3458 = a3456 & a3412;
assign a3460 = ~a3458 & a1936;
assign a3462 = ~l338 & l320;
assign a3464 = ~l320 & i92;
assign a3466 = ~a3464 & ~a3462;
assign a3468 = ~a3466 & ~a3114;
assign a3470 = ~a3468 & ~a3460;
assign a3472 = a3470 & ~a3410;
assign a3474 = a3472 & a1942;
assign a3476 = a3474 & a3372;
assign a3478 = a3476 & a3344;
assign a3480 = a3478 & a3322;
assign a3482 = a3480 & a3302;
assign a3484 = a3482 & a3214;
assign a3486 = a3484 & ~a3124;
assign a3488 = ~a3470 & a1942;
assign a3490 = a3488 & a3344;
assign a3492 = a3490 & ~a3322;
assign a3494 = a3492 & a3372;
assign a3496 = a3494 & a3302;
assign a3498 = a3496 & a3214;
assign a3500 = a3498 & ~a3124;
assign a3502 = a3500 & ~a3410;
assign a3504 = ~a3502 & ~a3486;
assign a3506 = a3490 & a3322;
assign a3508 = a3506 & ~a3302;
assign a3510 = a3508 & a3372;
assign a3512 = a3510 & ~a3214;
assign a3514 = a3512 & a3124;
assign a3516 = a3514 & ~a3410;
assign a3518 = a3372 & a1942;
assign a3520 = a3470 & a3410;
assign a3522 = a3520 & a3518;
assign a3524 = a3522 & ~a3124;
assign a3526 = a3524 & a3344;
assign a3528 = a3526 & ~a3322;
assign a3530 = a3528 & a3302;
assign a3532 = a3530 & ~a3214;
assign a3534 = ~a3532 & ~a3516;
assign a3536 = a3534 & a3504;
assign a3538 = a3480 & ~a3302;
assign a3540 = a3538 & a3214;
assign a3542 = a3540 & ~a3124;
assign a3544 = a3510 & a3214;
assign a3546 = a3544 & ~a3124;
assign a3548 = a3546 & ~a3410;
assign a3550 = a3488 & a3372;
assign a3552 = a3344 & a3322;
assign a3554 = a3410 & ~a3124;
assign a3556 = a3554 & a3552;
assign a3558 = ~a3302 & ~a3214;
assign a3560 = a3558 & a3556;
assign a3562 = a3560 & a3550;
assign a3564 = ~a3562 & ~a3548;
assign a3566 = a3564 & ~a3542;
assign a3568 = a3526 & a3322;
assign a3570 = a3568 & ~a3302;
assign a3572 = a3570 & ~a3214;
assign a3574 = a3478 & ~a3322;
assign a3576 = a3574 & ~a3302;
assign a3578 = a3576 & ~a3214;
assign a3580 = a3578 & ~a3124;
assign a3582 = ~a3580 & ~a3572;
assign a3584 = ~a3214 & ~a3124;
assign a3586 = a3506 & a3302;
assign a3588 = a3586 & a3372;
assign a3590 = a3588 & a3584;
assign a3592 = a3590 & a3410;
assign a3594 = a3302 & a3214;
assign a3596 = a3594 & a3556;
assign a3598 = a3596 & a3550;
assign a3600 = a3372 & ~a3214;
assign a3602 = ~a3302 & ~a3124;
assign a3604 = a3602 & a3410;
assign a3606 = a3604 & a3492;
assign a3608 = a3606 & a3600;
assign a3610 = ~a3608 & ~a3598;
assign a3612 = a3610 & ~a3592;
assign a3614 = a3612 & a3582;
assign a3616 = a3614 & a3566;
assign a3618 = a3616 & a3536;
assign a3620 = ~a3214 & a3124;
assign a3622 = a3620 & a3522;
assign a3624 = a3622 & a3344;
assign a3626 = a3624 & a3322;
assign a3628 = a3626 & ~a3302;
assign a3630 = ~a3344 & a3322;
assign a3632 = a3630 & a3474;
assign a3634 = a3632 & ~a3302;
assign a3636 = a3634 & a3124;
assign a3638 = a3636 & a3600;
assign a3640 = a3538 & ~a3214;
assign a3642 = a3640 & a3124;
assign a3644 = ~a3642 & ~a3638;
assign a3646 = a3644 & ~a3628;
assign a3648 = a3630 & a1942;
assign a3650 = a3648 & ~a3470;
assign a3652 = a3650 & a3372;
assign a3654 = a3652 & a3302;
assign a3656 = a3654 & ~a3214;
assign a3658 = a3656 & ~a3124;
assign a3660 = a3658 & a3410;
assign a3662 = ~a3344 & ~a3214;
assign a3664 = a3662 & a3322;
assign a3666 = a3664 & a3524;
assign a3668 = a3666 & a3302;
assign a3670 = ~a3344 & ~a3322;
assign a3672 = a3670 & a3524;
assign a3674 = a3672 & a3302;
assign a3676 = a3674 & ~a3214;
assign a3678 = ~a3676 & ~a3668;
assign a3680 = a3678 & ~a3660;
assign a3682 = ~a3344 & a3214;
assign a3684 = a3682 & a3322;
assign a3686 = a3550 & ~a3302;
assign a3688 = a3686 & a3124;
assign a3690 = a3688 & a3410;
assign a3692 = a3690 & a3684;
assign a3694 = a3652 & ~a3302;
assign a3696 = a3694 & a3214;
assign a3698 = a3696 & ~a3410;
assign a3700 = a3698 & a3124;
assign a3702 = ~a3700 & ~a3692;
assign a3704 = a3666 & ~a3302;
assign a3706 = a3656 & a3124;
assign a3708 = a3706 & a3410;
assign a3710 = ~a3708 & ~a3704;
assign a3712 = a3710 & a3702;
assign a3714 = a3712 & a3680;
assign a3716 = a3714 & a3646;
assign a3718 = a3716 & a3618;
assign a3720 = a3484 & a3124;
assign a3722 = a3632 & a3372;
assign a3724 = a3722 & a3302;
assign a3726 = a3724 & a3214;
assign a3728 = a3726 & a3124;
assign a3730 = ~a3728 & ~a3720;
assign a3732 = a3482 & ~a3214;
assign a3734 = ~a3410 & a3214;
assign a3736 = a3734 & a3588;
assign a3738 = a3654 & a3214;
assign a3740 = a3738 & ~a3410;
assign a3742 = ~a3740 & ~a3736;
assign a3744 = a3742 & ~a3732;
assign a3746 = a3744 & a3730;
assign a3748 = a3540 & a3124;
assign a3750 = a3722 & ~a3302;
assign a3752 = a3750 & a3214;
assign a3754 = a3752 & a3124;
assign a3756 = ~a3754 & ~a3748;
assign a3758 = a3650 & a3124;
assign a3760 = a3410 & ~a3302;
assign a3762 = a3760 & a3600;
assign a3764 = a3762 & a3758;
assign a3766 = ~a3372 & a1942;
assign a3768 = a3766 & a3344;
assign a3770 = a3768 & a3322;
assign a3772 = a3770 & ~a3302;
assign a3774 = a3772 & ~a3214;
assign a3776 = a3774 & a3124;
assign a3778 = a3776 & a3410;
assign a3780 = a3778 & ~a3470;
assign a3782 = ~a3780 & ~a3764;
assign a3784 = a3724 & ~a3214;
assign a3786 = a3784 & a3124;
assign a3788 = a3550 & a3302;
assign a3790 = a3662 & ~a3322;
assign a3792 = a3790 & a3788;
assign a3794 = a3792 & a3124;
assign a3796 = a3794 & ~a3410;
assign a3798 = ~a3796 & ~a3786;
assign a3800 = a3798 & a3782;
assign a3802 = a3800 & a3756;
assign a3804 = a3802 & a3746;
assign a3806 = a3648 & a3470;
assign a3808 = a3410 & a3302;
assign a3810 = a3808 & a3214;
assign a3812 = a3810 & a3372;
assign a3814 = a3812 & ~a3124;
assign a3816 = a3814 & a3806;
assign a3818 = a3726 & ~a3124;
assign a3820 = ~a3818 & ~a3816;
assign a3822 = a3772 & a3214;
assign a3824 = a3822 & a3124;
assign a3826 = a3824 & a3410;
assign a3828 = a3826 & ~a3470;
assign a3830 = a3770 & a3302;
assign a3832 = a3830 & ~a3214;
assign a3834 = a3832 & a3470;
assign a3836 = a3834 & a3124;
assign a3838 = a3836 & a3410;
assign a3840 = ~a3838 & ~a3828;
assign a3842 = a3586 & a3124;
assign a3844 = a3842 & ~a3410;
assign a3846 = a3844 & a3600;
assign a3848 = ~a3846 & a3840;
assign a3850 = a3848 & a3820;
assign a3852 = a3696 & a3554;
assign a3854 = a3544 & a3124;
assign a3856 = a3854 & ~a3410;
assign a3858 = ~a3856 & ~a3852;
assign a3860 = a3672 & ~a3302;
assign a3862 = a3860 & a3214;
assign a3864 = a3650 & a3604;
assign a3866 = a3864 & a3600;
assign a3868 = ~a3866 & ~a3862;
assign a3870 = a3752 & ~a3124;
assign a3872 = a3686 & a3670;
assign a3874 = a3872 & a3584;
assign a3876 = a3874 & a3410;
assign a3878 = ~a3876 & ~a3870;
assign a3880 = a3878 & a3868;
assign a3882 = a3880 & a3858;
assign a3884 = a3882 & a3850;
assign a3886 = a3884 & a3804;
assign a3888 = a3886 & a3718;
assign a3890 = a3522 & ~a3302;
assign a3892 = a3214 & a3124;
assign a3894 = a3892 & a3890;
assign a3896 = a3788 & a3214;
assign a3898 = a3896 & a3124;
assign a3900 = a3898 & a3410;
assign a3902 = ~a3900 & ~a3894;
assign a3904 = ~a3902 & a3552;
assign a3906 = a3738 & a3124;
assign a3908 = a3906 & a3410;
assign a3910 = a3894 & a3630;
assign a3912 = ~a3910 & ~a3908;
assign a3914 = a3604 & a3214;
assign a3916 = a3914 & a3372;
assign a3918 = a3916 & a3806;
assign a3920 = a3738 & ~a3124;
assign a3922 = a3920 & a3410;
assign a3924 = ~a3922 & ~a3918;
assign a3926 = a3924 & a3912;
assign a3928 = a3926 & ~a3904;
assign a3930 = a3842 & a3410;
assign a3932 = a3930 & a3600;
assign a3934 = a3514 & a3410;
assign a3936 = ~a3934 & ~a3932;
assign a3938 = a3936 & a3928;
assign a3940 = a3854 & a3410;
assign a3942 = a3626 & a3302;
assign a3944 = ~a3942 & ~a3940;
assign a3946 = a3546 & a3410;
assign a3948 = a3568 & a3302;
assign a3950 = a3948 & ~a3214;
assign a3952 = ~a3950 & ~a3946;
assign a3954 = a3952 & a3944;
assign a3956 = ~a3410 & ~a3124;
assign a3958 = a3956 & a3512;
assign a3960 = a3810 & a3124;
assign a3962 = a3960 & a3806;
assign a3964 = a3962 & a3372;
assign a3966 = ~a3964 & ~a3958;
assign a3968 = a3622 & ~a3344;
assign a3970 = a3968 & a3322;
assign a3972 = a3768 & ~a3322;
assign a3974 = a3972 & a3302;
assign a3976 = a3974 & a3214;
assign a3978 = a3976 & a3124;
assign a3980 = a3978 & a3410;
assign a3982 = ~a3980 & ~a3970;
assign a3984 = a3982 & a3966;
assign a3986 = a3984 & a3954;
assign a3988 = a3986 & a3938;
assign a3990 = a3688 & ~a3410;
assign a3992 = a3990 & a3664;
assign a3994 = a3570 & a3214;
assign a3996 = ~a3994 & ~a3992;
assign a3998 = ~a3784 & ~a3698;
assign a4000 = ~a3998 & ~a3124;
assign a4002 = a3670 & a3476;
assign a4004 = a4002 & ~a3302;
assign a4006 = a4004 & a3214;
assign a4008 = a4006 & ~a3124;
assign a4010 = a3792 & ~a3124;
assign a4012 = a4010 & a3410;
assign a4014 = ~a4012 & ~a4008;
assign a4016 = a4014 & ~a4000;
assign a4018 = a4016 & a3996;
assign a4020 = a3948 & a3214;
assign a4022 = a3860 & ~a3214;
assign a4024 = a3990 & a3790;
assign a4026 = a3674 & a3214;
assign a4028 = ~a4026 & ~a4024;
assign a4030 = a4028 & ~a4022;
assign a4032 = a4002 & a3302;
assign a4034 = a4032 & a3214;
assign a4036 = a4034 & ~a3124;
assign a4038 = a3670 & a3488;
assign a4040 = ~a3916 & ~a3814;
assign a4042 = ~a4040 & a4038;
assign a4044 = ~a4042 & ~a4036;
assign a4046 = a4044 & a4030;
assign a4048 = a4046 & ~a4020;
assign a4050 = a4048 & a4018;
assign a4052 = a4050 & a3988;
assign a4054 = a3640 & ~a3124;
assign a4056 = a3590 & ~a3410;
assign a4058 = ~a4056 & ~a4054;
assign a4060 = a3496 & ~a3214;
assign a4062 = a4060 & ~a3124;
assign a4064 = a4062 & a3410;
assign a4066 = a3528 & ~a3302;
assign a4068 = a4066 & ~a3214;
assign a4070 = a3968 & ~a3322;
assign a4072 = a4070 & ~a3302;
assign a4074 = ~a4072 & ~a4068;
assign a4076 = a4074 & ~a4064;
assign a4078 = a4076 & a4058;
assign a4080 = a3574 & a3302;
assign a4082 = a4080 & ~a3214;
assign a4084 = a4082 & ~a3124;
assign a4086 = ~a3410 & ~a3214;
assign a4088 = a3602 & a3494;
assign a4090 = a4088 & a4086;
assign a4092 = a3576 & a3214;
assign a4094 = a4092 & ~a3124;
assign a4096 = ~a4094 & ~a4090;
assign a4098 = a4096 & ~a4084;
assign a4100 = a4098 & a4078;
assign a4102 = a4080 & a3214;
assign a4104 = a4102 & ~a3124;
assign a4106 = a4062 & ~a3410;
assign a4108 = a4088 & a3214;
assign a4110 = a4108 & ~a3410;
assign a4112 = ~a4110 & ~a4106;
assign a4114 = a4112 & ~a4104;
assign a4116 = a4032 & ~a3214;
assign a4118 = a4116 & ~a3124;
assign a4120 = a3874 & ~a3410;
assign a4122 = ~a4120 & ~a4118;
assign a4124 = a3830 & a3214;
assign a4126 = a4124 & a3470;
assign a4128 = a4126 & a3124;
assign a4130 = a4128 & ~a3410;
assign a4132 = a3972 & ~a3302;
assign a4134 = a4132 & a3214;
assign a4136 = a4134 & a3124;
assign a4138 = a4136 & a3410;
assign a4140 = a4138 & a3470;
assign a4142 = ~a4140 & ~a4130;
assign a4144 = a4142 & a4122;
assign a4146 = a3872 & a3214;
assign a4148 = a4146 & a3124;
assign a4150 = a4148 & a3410;
assign a4152 = a3518 & ~a3322;
assign a4154 = a3808 & a3470;
assign a4156 = a4154 & a3682;
assign a4158 = a4156 & a4152;
assign a4160 = a4158 & a3124;
assign a4162 = ~a4160 & ~a4150;
assign a4164 = a3794 & a3410;
assign a4166 = a4070 & a3302;
assign a4168 = ~a4166 & ~a4164;
assign a4170 = a3706 & ~a3410;
assign a4172 = ~a2964 & ~a1942;
assign a4174 = ~a4172 & ~a4170;
assign a4176 = a4174 & a4168;
assign a4178 = a4176 & a4162;
assign a4180 = a4178 & a4144;
assign a4182 = a4180 & a4114;
assign a4184 = a4182 & a4100;
assign a4186 = a4184 & a4052;
assign a4190 = a2404 & i94;
assign a4192 = ~a2404 & l322;
assign a4194 = ~a4192 & ~a4190;
assign a4196 = a3530 & a3214;
assign a4198 = ~a4196 & ~a4068;
assign a4200 = a4198 & a4114;
assign a4202 = a3500 & a3410;
assign a4204 = ~a4202 & a4200;
assign a4206 = ~a3470 & ~a3124;
assign a4208 = a4206 & a4124;
assign a4210 = a4208 & ~a3410;
assign a4212 = a3956 & a3834;
assign a4214 = ~a4212 & ~a4210;
assign a4216 = a4214 & a4058;
assign a4218 = a4216 & a3952;
assign a4220 = a3832 & ~a3124;
assign a4222 = ~a3470 & ~a3410;
assign a4224 = a4222 & a4220;
assign a4226 = a3822 & a3554;
assign a4228 = a4226 & a3470;
assign a4230 = ~a4228 & ~a4224;
assign a4232 = a4220 & a3410;
assign a4234 = a4232 & ~a3470;
assign a4236 = a3776 & ~a3410;
assign a4238 = a4236 & ~a3470;
assign a4240 = ~a4238 & ~a4234;
assign a4242 = a4240 & a4230;
assign a4244 = ~a4020 & ~a3994;
assign a4246 = a4244 & a4242;
assign a4248 = a3976 & ~a3124;
assign a4250 = a4248 & ~a3410;
assign a4252 = a4250 & ~a3470;
assign a4254 = a4248 & a3410;
assign a4256 = a4254 & ~a3470;
assign a4258 = ~a4256 & ~a4252;
assign a4260 = a3974 & ~a3214;
assign a4262 = a4260 & a3554;
assign a4264 = a4262 & ~a3470;
assign a4266 = ~a3120 & ~a1942;
assign a4268 = ~a4266 & ~a4264;
assign a4270 = a4268 & a4258;
assign a4272 = a4262 & a3470;
assign a4274 = a4254 & a3470;
assign a4276 = ~a4274 & ~a4272;
assign a4278 = a4126 & a3956;
assign a4280 = a4232 & a3470;
assign a4282 = ~a4280 & ~a4278;
assign a4284 = a4282 & a4276;
assign a4286 = a4284 & a4270;
assign a4288 = a4286 & a4246;
assign a4290 = a4288 & a4218;
assign a4292 = a4290 & a4204;
assign a4294 = a3670 & ~a3410;
assign a4296 = a4294 & ~a3124;
assign a4298 = a4296 & a3896;
assign a4300 = ~a4298 & ~a4042;
assign a4302 = a3766 & a3630;
assign a4304 = a4302 & a3302;
assign a4306 = a4304 & a3214;
assign a4308 = a4306 & ~a3124;
assign a4310 = ~a4308 & a4300;
assign a4312 = ~a4036 & ~a4008;
assign a4314 = a4312 & a3820;
assign a4316 = a4314 & a4310;
assign a4318 = a4316 & a3880;
assign a4320 = a4304 & ~a3214;
assign a4322 = a4320 & ~a3124;
assign a4324 = a4322 & ~a3410;
assign a4326 = ~a4324 & ~a4118;
assign a4328 = a4322 & a3410;
assign a4330 = ~a4328 & a3680;
assign a4332 = a4330 & a4326;
assign a4334 = a4028 & a3924;
assign a4336 = a4334 & a4332;
assign a4338 = ~a4012 & ~a3704;
assign a4340 = a4004 & a3584;
assign a4342 = a3750 & a3584;
assign a4344 = ~a4342 & ~a4340;
assign a4346 = a4344 & ~a4022;
assign a4348 = a4346 & a4338;
assign a4350 = a3920 & ~a3410;
assign a4352 = ~a4350 & ~a3852;
assign a4354 = a4352 & ~a4000;
assign a4356 = a4354 & a4348;
assign a4358 = a4356 & a4336;
assign a4360 = a4358 & a4318;
assign a4362 = a4098 & ~a4064;
assign a4364 = ~a3736 & ~a3732;
assign a4366 = ~a4364 & ~a3124;
assign a4368 = ~a4366 & a4362;
assign a4370 = a4368 & a3618;
assign a4372 = a4370 & a4360;
assign a4376 = ~a4150 & a3702;
assign a4378 = a4376 & ~a4000;
assign a4380 = a4138 & ~a3470;
assign a4382 = ~a4380 & ~a3828;
assign a4384 = ~a3210 & ~a1942;
assign a4386 = ~a4384 & a4382;
assign a4388 = a4386 & ~a3548;
assign a4390 = a4388 & a4378;
assign a4392 = ~a4110 & ~a4084;
assign a4394 = a4392 & a3858;
assign a4396 = a4394 & a3954;
assign a4398 = a4396 & a4390;
assign a4400 = a3578 & a3124;
assign a4402 = a4236 & a3470;
assign a4404 = a3778 & a3470;
assign a4406 = ~a4404 & ~a4402;
assign a4408 = a4406 & ~a4400;
assign a4410 = a4408 & a3582;
assign a4412 = a4348 & a3646;
assign a4414 = a4412 & a4078;
assign a4416 = a4414 & a4410;
assign a4418 = a4320 & a3124;
assign a4420 = a4418 & ~a3410;
assign a4422 = a4420 & ~a3470;
assign a4424 = ~a4422 & ~a4170;
assign a4426 = a4424 & ~a3992;
assign a4428 = a4426 & ~a3708;
assign a4430 = a4116 & a3124;
assign a4432 = ~a4430 & a4428;
assign a4434 = a4420 & a3470;
assign a4436 = ~a4434 & ~a3970;
assign a4438 = a4436 & a4168;
assign a4440 = a4438 & a3798;
assign a4442 = a4440 & a4432;
assign a4444 = a3624 & ~a3322;
assign a4446 = a4444 & a3302;
assign a4448 = ~a4446 & ~a3532;
assign a4450 = a4448 & ~a3732;
assign a4452 = a4450 & a4442;
assign a4454 = a4260 & a3124;
assign a4456 = a4454 & ~a3410;
assign a4458 = a4456 & ~a3470;
assign a4460 = ~a4458 & ~a3846;
assign a4462 = ~a4224 & ~a4090;
assign a4464 = a4462 & ~a4106;
assign a4466 = a4464 & a4460;
assign a4468 = a4418 & a3410;
assign a4470 = a4468 & ~a3470;
assign a4472 = ~a4470 & ~a4234;
assign a4474 = a4454 & a3410;
assign a4476 = a4474 & ~a3470;
assign a4478 = ~a4476 & ~a4264;
assign a4480 = a4478 & ~a3592;
assign a4482 = a4480 & a4472;
assign a4484 = a4482 & a3936;
assign a4486 = a4484 & a4466;
assign a4488 = a4468 & a3470;
assign a4490 = ~a4488 & ~a4212;
assign a4492 = a4490 & ~a4280;
assign a4494 = a4456 & a3470;
assign a4496 = ~a4272 & ~a3838;
assign a4498 = a4496 & ~a4494;
assign a4500 = a4498 & a4492;
assign a4502 = a4500 & a4332;
assign a4504 = a4502 & a4486;
assign a4506 = a4504 & a4452;
assign a4508 = a4506 & a4416;
assign a4512 = a3978 & ~a3410;
assign a4514 = ~a4278 & ~a4130;
assign a4516 = a4514 & ~a4512;
assign a4518 = a4516 & ~a4104;
assign a4520 = a4102 & a3124;
assign a4522 = ~a4520 & ~a4094;
assign a4524 = a4522 & a3504;
assign a4526 = a4524 & a4518;
assign a4528 = a3976 & a3520;
assign a4530 = a4306 & a3124;
assign a4532 = ~a4530 & ~a4160;
assign a4534 = a4152 & a3344;
assign a4536 = a4534 & a3470;
assign a4538 = a4536 & a3960;
assign a4540 = ~a3298 & ~a1942;
assign a4542 = ~a4540 & ~a4538;
assign a4544 = a4542 & a4532;
assign a4546 = a4544 & ~a4528;
assign a4548 = a4546 & a4244;
assign a4550 = a4548 & a4316;
assign a4552 = a4550 & a4526;
assign a4554 = a3498 & a3124;
assign a4556 = a4554 & a3410;
assign a4558 = a3980 & ~a3470;
assign a4560 = ~a4558 & ~a4210;
assign a4562 = a4560 & a4258;
assign a4564 = a4562 & ~a4556;
assign a4566 = a4554 & ~a3410;
assign a4568 = a4294 & a3898;
assign a4570 = ~a4568 & ~a4566;
assign a4572 = a3742 & ~a3598;
assign a4574 = a4572 & a4570;
assign a4576 = a4574 & a4564;
assign a4578 = ~a4202 & ~a4196;
assign a4580 = a4578 & a3730;
assign a4582 = a4580 & a4576;
assign a4584 = a4582 & a4506;
assign a4588 = ~a4380 & ~a4340;
assign a4590 = a4588 & a4362;
assign a4592 = ~a4538 & a4122;
assign a4594 = a4592 & a4590;
assign a4596 = ~a4556 & a4162;
assign a4598 = a4512 & a3470;
assign a4600 = ~a4598 & ~a4458;
assign a4602 = a4600 & a4478;
assign a4604 = a4276 & ~a4256;
assign a4606 = a4604 & a4602;
assign a4608 = a4606 & a4596;
assign a4610 = a4608 & a4200;
assign a4612 = a4610 & a4594;
assign a4614 = ~a4430 & ~a4400;
assign a4616 = a4614 & a4570;
assign a4618 = ~a4494 & ~a4252;
assign a4620 = a4618 & a4312;
assign a4622 = a3790 & a3690;
assign a4624 = ~a3876 & ~a3608;
assign a4626 = a4624 & ~a4622;
assign a4628 = a4626 & ~a3580;
assign a4630 = a4628 & a4620;
assign a4632 = a4630 & a4616;
assign a4634 = a4512 & ~a3470;
assign a4636 = ~a4634 & ~a4140;
assign a4638 = a3894 & a3670;
assign a4640 = ~a4638 & ~a3794;
assign a4642 = a4640 & a4636;
assign a4644 = a4300 & ~a3862;
assign a4646 = a4644 & ~a3500;
assign a4648 = a4646 & a4642;
assign a4650 = a4648 & ~a4520;
assign a4652 = ~a4166 & ~a3980;
assign a4654 = a4652 & a4448;
assign a4656 = ~a3318 & ~a1942;
assign a4658 = ~a4656 & ~a3676;
assign a4660 = ~a4072 & ~a4012;
assign a4662 = a4660 & a4658;
assign a4664 = a4662 & a4030;
assign a4666 = a4664 & a4654;
assign a4668 = a4666 & a4650;
assign a4670 = a4668 & a4632;
assign a4674 = ~a4568 & ~a3638;
assign a4676 = a4674 & a4376;
assign a4678 = ~a3754 & ~a3728;
assign a4680 = a4678 & a3966;
assign a4682 = a4680 & a4676;
assign a4684 = ~a3340 & ~a1942;
assign a4686 = ~a4684 & ~a3764;
assign a4688 = a4686 & ~a4468;
assign a4690 = a4688 & ~a4638;
assign a4692 = a4690 & a3912;
assign a4694 = ~a4622 & ~a4072;
assign a4696 = a3906 & ~a3410;
assign a4698 = ~a4696 & a4532;
assign a4700 = a4698 & a4694;
assign a4702 = a4700 & a4692;
assign a4704 = a4702 & a4442;
assign a4706 = a4704 & a4682;
assign a4710 = a4530 & a3520;
assign a4712 = ~a4710 & a4242;
assign a4714 = a4308 & ~a3410;
assign a4716 = ~a4714 & ~a4434;
assign a4718 = a4716 & ~a4402;
assign a4720 = a4718 & a4500;
assign a4722 = a4720 & a4712;
assign a4724 = a4636 & a4562;
assign a4726 = a3826 & a3470;
assign a4728 = ~a4726 & ~a4404;
assign a4730 = a3824 & a3472;
assign a4732 = a3694 & ~a3124;
assign a4734 = a4732 & a4086;
assign a4736 = ~a4734 & ~a4730;
assign a4738 = a4736 & a4728;
assign a4740 = ~a4530 & ~a4322;
assign a4742 = ~a4740 & a4222;
assign a4744 = ~a4742 & ~a3780;
assign a4746 = a4744 & a4514;
assign a4748 = a4746 & a4738;
assign a4750 = a4748 & a4724;
assign a4752 = a4308 & a3520;
assign a4754 = ~a4752 & ~a4470;
assign a4756 = a4306 & ~a3470;
assign a4758 = a4756 & a3410;
assign a4760 = ~a4758 & ~a4328;
assign a4762 = a4760 & a4754;
assign a4764 = ~a4740 & a3472;
assign a4766 = ~a4764 & a4382;
assign a4768 = a4766 & a4762;
assign a4770 = ~a3368 & ~a1942;
assign a4772 = ~a4770 & ~a4422;
assign a4774 = a4772 & ~a4120;
assign a4776 = a4774 & ~a4528;
assign a4778 = a4776 & a4602;
assign a4780 = a4778 & a4768;
assign a4782 = a4780 & a4750;
assign a4786 = a4530 & ~a3410;
assign a4788 = ~a4786 & ~a4298;
assign a4790 = a4788 & a4718;
assign a4792 = a4790 & a4426;
assign a4794 = a4216 & ~a4000;
assign a4796 = a4794 & a4792;
assign a4798 = a4344 & ~a3818;
assign a4800 = a4798 & a4392;
assign a4802 = a4800 & a3804;
assign a4804 = a4802 & a4796;
assign a4806 = ~a3406 & ~a1942;
assign a4808 = ~a4806 & ~a3866;
assign a4810 = a4808 & ~a3700;
assign a4812 = a4810 & a4326;
assign a4814 = a4812 & a4466;
assign a4816 = a4814 & a4632;
assign a4818 = ~a4730 & ~a3870;
assign a4820 = a4818 & ~a3856;
assign a4822 = a4820 & a3644;
assign a4824 = a4822 & a3566;
assign a4826 = a4824 & a4526;
assign a4828 = a4826 & a4816;
assign a4832 = a4648 & ~a3542;
assign a4834 = a4832 & a4576;
assign a4836 = a4834 & a4486;
assign a4838 = ~a4714 & ~a4328;
assign a4840 = ~a4838 & ~a3470;
assign a4842 = ~a4840 & ~a3660;
assign a4844 = a4842 & a4428;
assign a4846 = a4844 & a3756;
assign a4848 = ~a4742 & ~a4726;
assign a4850 = ~a3466 & ~a1942;
assign a4852 = ~a4850 & ~a4228;
assign a4854 = a4852 & ~a4758;
assign a4856 = a4854 & a4848;
assign a4858 = a4856 & a4818;
assign a4860 = a4858 & a3928;
assign a4862 = a4860 & a4846;
assign a4864 = a4862 & a4416;
assign a4868 = a1936 & l322;
assign a4870 = ~a1948 & l340;
assign a4872 = ~a4870 & ~a4868;
assign a4874 = l314 & l138;
assign a4876 = ~a4874 & ~l236;
assign a4878 = a4876 & a2990;
assign a4880 = a4878 & i98;
assign a4882 = ~a4878 & l342;
assign a4884 = ~a4882 & ~a4880;
assign a4886 = a4878 & i100;
assign a4888 = ~a4878 & l344;
assign a4890 = ~a4888 & ~a4886;
assign a4892 = ~l368 & l320;
assign a4894 = ~l320 & i112;
assign a4896 = ~a4894 & ~a4892;
assign a4898 = ~a4896 & a506;
assign a4900 = ~a506 & l346;
assign a4902 = ~a4900 & ~a4898;
assign a4904 = ~l366 & l320;
assign a4906 = ~l320 & i110;
assign a4908 = ~a4906 & ~a4904;
assign a4910 = ~a4908 & a506;
assign a4912 = ~a506 & l348;
assign a4914 = ~a4912 & ~a4910;
assign a4916 = ~l364 & l320;
assign a4918 = ~l320 & i108;
assign a4920 = ~a4918 & ~a4916;
assign a4922 = ~a4920 & a506;
assign a4924 = ~a506 & l350;
assign a4926 = ~a4924 & ~a4922;
assign a4928 = ~l362 & l320;
assign a4930 = ~l320 & i106;
assign a4932 = ~a4930 & ~a4928;
assign a4934 = ~a4932 & a506;
assign a4936 = ~a506 & l352;
assign a4938 = ~a4936 & ~a4934;
assign a4940 = ~l360 & l320;
assign a4942 = ~l320 & i104;
assign a4944 = ~a4942 & ~a4940;
assign a4946 = ~a4944 & a506;
assign a4948 = ~a506 & l354;
assign a4950 = ~a4948 & ~a4946;
assign a4952 = ~l358 & l320;
assign a4954 = ~l320 & ~i102;
assign a4956 = ~a4954 & ~a4952;
assign a4958 = a4956 & a506;
assign a4960 = ~a506 & l356;
assign a4962 = ~a4960 & ~a4958;
assign a4966 = a4226 & ~a3470;
assign a4968 = ~a4966 & a4762;
assign a4970 = ~a4944 & ~a1942;
assign a4972 = ~a4970 & ~a3980;
assign a4974 = a4972 & a4968;
assign a4976 = a4060 & a3124;
assign a4978 = a4976 & a3410;
assign a4980 = ~a4978 & a4246;
assign a4982 = a4980 & a4974;
assign a4984 = a4796 & a4594;
assign a4988 = ~a4932 & ~a1942;
assign a4990 = ~a4988 & a4014;
assign a4994 = a4092 & a3124;
assign a4996 = a4108 & a3410;
assign a4998 = a4148 & ~a3410;
assign a5000 = ~a4998 & ~a4996;
assign a5002 = a5000 & ~a4994;
assign a5004 = ~a3372 & ~a3214;
assign a5006 = ~a3930 & ~a3606;
assign a5008 = ~a5006 & a5004;
assign a5010 = a4976 & ~a3410;
assign a5012 = ~a5010 & ~a5008;
assign a5014 = a4066 & a3214;
assign a5016 = a3344 & ~a3322;
assign a5018 = a5016 & a3214;
assign a5020 = a5018 & a3990;
assign a5022 = a4146 & a3956;
assign a5024 = ~a5022 & ~a5020;
assign a5026 = a5024 & ~a5014;
assign a5028 = a3772 & a3472;
assign a5030 = a3972 & ~a3214;
assign a5032 = a5030 & a3470;
assign a5034 = a5032 & a3760;
assign a5036 = ~a5034 & ~a5028;
assign a5038 = ~a5036 & ~a3124;
assign a5040 = ~a3372 & a3214;
assign a5042 = a5040 & a3606;
assign a5044 = ~a5042 & ~a5038;
assign a5046 = a4134 & ~a3124;
assign a5048 = a5046 & a3470;
assign a5050 = a5048 & a3410;
assign a5052 = a3476 & a3124;
assign a5054 = a3790 & ~a3302;
assign a5056 = a5054 & a5052;
assign a5058 = a3766 & a3470;
assign a5060 = ~a3596 & ~a3560;
assign a5062 = ~a5060 & a5058;
assign a5064 = ~a5062 & ~a5056;
assign a5066 = a5064 & ~a5050;
assign a5068 = a5066 & a5044;
assign a5070 = a5068 & a5026;
assign a5072 = a5070 & a5012;
assign a5074 = a5072 & a5002;
assign a5076 = a4058 & a4018;
assign a5078 = a5076 & a5074;
assign a5080 = a4302 & ~a3302;
assign a5082 = a5080 & a3520;
assign a5084 = a5082 & ~a3124;
assign a5086 = ~a5084 & ~a4130;
assign a5088 = a4474 & a3470;
assign a5090 = a4206 & a3774;
assign a5092 = a5090 & a3410;
assign a5094 = a5004 & a3864;
assign a5096 = a5080 & a3214;
assign a5098 = a5096 & a4222;
assign a5100 = ~a5098 & ~a5094;
assign a5102 = a5100 & ~a5092;
assign a5104 = a5102 & ~a5088;
assign a5106 = a5104 & a5086;
assign a5108 = a5004 & a3636;
assign a5110 = a4136 & ~a3410;
assign a5112 = a5110 & ~a3470;
assign a5114 = ~a5112 & ~a5108;
assign a5116 = a5114 & a4694;
assign a5118 = a5116 & a5106;
assign a5120 = a3900 & a3670;
assign a5122 = a4010 & ~a3410;
assign a5124 = a5110 & a3470;
assign a5126 = ~a5124 & ~a5122;
assign a5128 = a5126 & ~a5120;
assign a5130 = ~a3864 & ~a3634;
assign a5132 = a3956 & a3508;
assign a5134 = ~a5132 & ~a3842;
assign a5136 = a5134 & a5130;
assign a5138 = ~a5136 & a5040;
assign a5140 = ~a5138 & a5128;
assign a5142 = a5140 & a5118;
assign a5144 = a5016 & a3894;
assign a5146 = ~a5144 & ~a4140;
assign a5148 = a5146 & a4588;
assign a5150 = a5148 & a5142;
assign a5152 = a5150 & a5078;
assign a5154 = a4128 & a3410;
assign a5156 = a5032 & a3956;
assign a5158 = ~a5156 & ~a5154;
assign a5160 = a5048 & ~a3410;
assign a5162 = ~a5160 & ~a4252;
assign a5164 = a5162 & a4738;
assign a5166 = a5164 & a3888;
assign a5168 = a5166 & a5158;
assign a5170 = a5168 & ~a3980;
assign a5172 = a5170 & a5152;
assign a5174 = a4444 & ~a3302;
assign a5176 = ~a5174 & a4214;
assign a5178 = a5176 & a4592;
assign a5180 = a5178 & a4712;
assign a5182 = a5180 & a4048;
assign a5184 = a4208 & a3410;
assign a5186 = a5046 & a4222;
assign a5188 = ~a5186 & ~a5184;
assign a5190 = a4132 & a3620;
assign a5192 = a5190 & a3410;
assign a5194 = a5192 & a3470;
assign a5196 = a5096 & a3124;
assign a5198 = a5196 & a3410;
assign a5200 = a5198 & ~a3470;
assign a5202 = ~a5200 & ~a5194;
assign a5204 = a5202 & a5188;
assign a5206 = ~a4634 & ~a4494;
assign a5208 = a5206 & a5204;
assign a5210 = a5132 & a5004;
assign a5212 = a4250 & a3470;
assign a5214 = ~a5212 & ~a5210;
assign a5216 = a5192 & ~a3470;
assign a5218 = ~a5216 & ~a4324;
assign a5220 = a5218 & ~a4446;
assign a5222 = a5220 & a5214;
assign a5224 = a5222 & a5208;
assign a5226 = a5224 & a4608;
assign a5228 = a5018 & a3690;
assign a5230 = a3836 & ~a3410;
assign a5232 = ~a5230 & ~a5228;
assign a5234 = a5232 & a4424;
assign a5236 = a5234 & a4790;
assign a5238 = a3634 & ~a3124;
assign a5240 = a5238 & a5004;
assign a5242 = a5080 & ~a3214;
assign a5244 = a5242 & ~a3124;
assign a5246 = a5244 & a4222;
assign a5248 = ~a5246 & ~a4488;
assign a5250 = a5248 & ~a5240;
assign a5252 = a5250 & a4282;
assign a5254 = a5252 & a4968;
assign a5256 = a5254 & a5236;
assign a5258 = a5256 & a5226;
assign a5260 = a5258 & a5182;
assign a5262 = ~a4978 & a4578;
assign a5264 = a4034 & a3124;
assign a5266 = ~a5190 & ~a3824;
assign a5268 = ~a5266 & a4222;
assign a5270 = ~a5268 & ~a5264;
assign a5272 = a4082 & a3124;
assign a5274 = a5190 & a3472;
assign a5276 = ~a5274 & ~a4638;
assign a5278 = a5276 & a4168;
assign a5280 = a5278 & ~a5272;
assign a5282 = a5280 & a5270;
assign a5284 = ~a4920 & ~a1942;
assign a5286 = a5004 & a3844;
assign a5288 = a5242 & a3124;
assign a5290 = ~a4222 & ~a3520;
assign a5292 = ~a5290 & a5288;
assign a5294 = ~a5292 & ~a5286;
assign a5296 = a5294 & ~a5284;
assign a5298 = a5296 & a5282;
assign a5300 = a5298 & a5262;
assign a5302 = a5300 & a5260;
assign a5306 = a3658 & ~a3410;
assign a5308 = ~a5306 & ~a4342;
assign a5310 = a5308 & a5282;
assign a5312 = a5310 & a4204;
assign a5314 = a5288 & a3410;
assign a5316 = a5314 & ~a3470;
assign a5318 = a5198 & a3470;
assign a5320 = ~a5318 & ~a5316;
assign a5322 = a5320 & a5294;
assign a5324 = ~a4908 & ~a1942;
assign a5326 = ~a5324 & a5322;
assign a5328 = a5326 & a5312;
assign a5330 = a5328 & a5074;
assign a5332 = a5226 & a5142;
assign a5334 = a5332 & a5166;
assign a5338 = a5016 & ~a3214;
assign a5340 = a5338 & a3688;
assign a5342 = a4006 & a3124;
assign a5344 = ~a5342 & ~a5340;
assign a5346 = ~a4978 & ~a4520;
assign a5348 = a5346 & a5344;
assign a5350 = a5348 & a4616;
assign a5352 = a5350 & a5312;
assign a5354 = a5352 & a5168;
assign a5356 = a5354 & a5322;
assign a5358 = ~a4896 & ~a1942;
assign a5360 = a5260 & a3988;
assign a5362 = a5360 & a5152;
assign a5364 = a5362 & ~a5358;
assign a5370 = ~a1942 & ~a652;
assign a5372 = ~a5370 & ~a3980;
assign a5374 = a5372 & a4590;
assign a5378 = a1604 & ~l194;
assign a5380 = ~a1700 & ~a1326;
assign a5382 = a5380 & ~a1476;
assign a5384 = a5382 & ~a5378;
assign a5386 = a5384 & a1860;
assign a5388 = ~a5386 & a506;
assign a5390 = ~a506 & l374;
assign a5392 = ~a5390 & ~a5388;
assign a5394 = a1874 & ~l206;
assign a5396 = ~a5394 & ~a1844;
assign a5398 = a5396 & ~a5378;
assign a5400 = a1356 & ~l188;
assign a5402 = ~a5400 & a1818;
assign a5404 = a5402 & a5398;
assign a5406 = a5404 & a2100;
assign a5408 = a1896 & a1644;
assign a5410 = a5408 & a5406;
assign a5412 = ~a5410 & a506;
assign a5414 = ~a506 & l376;
assign a5416 = ~a5414 & ~a5412;
assign a5420 = ~a1942 & ~a596;
assign a5424 = ~a1942 & ~a584;
assign a5426 = ~a5424 & a5354;
assign a5430 = ~a1942 & ~a572;
assign a5434 = a398 & i132;
assign a5436 = ~a398 & i134;
assign a5438 = ~a5436 & ~a5434;
assign a5440 = a5438 & l386;
assign a5442 = ~a5440 & ~a1910;
assign a5444 = i134 & ~i132;
assign a5446 = ~a5444 & ~a2346;
assign a5448 = a5446 & ~a2350;
assign a5450 = a5448 & ~a2406;
assign a5452 = a5450 & a2380;
assign a5454 = a5452 & ~a2348;
assign a5456 = ~a5454 & a1910;
assign a5460 = a2392 & ~a2380;
assign a5462 = a5460 & a1942;
assign a5464 = ~a5462 & i132;
assign a5466 = a5462 & a2400;
assign a5468 = ~a2388 & ~a2340;
assign a5470 = ~a5468 & ~a2342;
assign a5472 = ~a1910 & ~a398;
assign a5474 = ~a5472 & ~a5470;
assign a5476 = a2380 & ~a1940;
assign a5478 = ~a5476 & ~a2378;
assign a5480 = ~a5478 & a5474;
assign a5482 = a5480 & ~a2384;
assign a5484 = a5482 & ~a5466;
assign a5488 = l390 & i130;
assign a5490 = a5488 & a392;
assign a5492 = a420 & i70;
assign a5494 = ~a5492 & ~a5490;
assign a5496 = ~l170 & l168;
assign a5498 = a5496 & l166;
assign a5500 = a5498 & l162;
assign a5502 = ~l172 & l158;
assign a5504 = ~a5502 & ~a5500;
assign a5506 = ~l170 & ~l168;
assign a5508 = a5506 & l166;
assign a5510 = a5508 & l160;
assign a5512 = a5496 & ~l166;
assign a5514 = a5512 & l164;
assign a5516 = ~a5514 & ~a5510;
assign a5518 = a5516 & a5504;
assign a5520 = a5508 & i10;
assign a5522 = ~a5520 & ~a616;
assign a5524 = a5498 & i12;
assign a5526 = a5512 & i14;
assign a5528 = ~a5526 & ~a5524;
assign a5530 = a5528 & a5522;
assign a5532 = ~a5530 & l174;
assign a5534 = a5498 & i6;
assign a5536 = ~l172 & l142;
assign a5538 = ~a5536 & ~a5534;
assign a5540 = a5508 & i4;
assign a5542 = a5512 & i8;
assign a5544 = ~a5542 & ~a5540;
assign a5546 = a5544 & a5538;
assign a5548 = ~a5546 & a5532;
assign a5550 = ~a5548 & ~a5518;
assign a5552 = a5548 & a5518;
assign a5554 = ~a5552 & ~a5550;
assign a5556 = ~a5554 & a420;
assign a5558 = a5556 & a502;
assign a5560 = a5554 & a500;
assign a5562 = ~a5560 & ~a5558;
assign p0 = ~a5562;

assert property (~p0);

endmodule
