module m6s1 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474,i476,i478,i480,
i482,i484,i486,i488,i490,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474,i476,i478,i480,
i482,i484,i486,i488,i490;

output p0;

wire a6662,a6682,a6690,a6696,a6702,a6708,na6710,a6712,a6074,a6920,a7152,a7352,a7590,a7812,a7852,
a7864,a7900,a7930,a7942,a7954,a7966,a7978,a7990,a8002,a8020,a16268,a16274,a16280,a16286,a16292,
a16298,a16304,a16310,a16660,a16800,a16936,a17072,a17208,a17342,a17476,a17610,a17742,a17872,a15370,a15474,
a15578,a15682,a15786,a15884,a15982,na2430,a17882,na2432,na2436,a17900,a17916,na2434,na5594,na5596,na5600,
na5598,a6592,a6476,a6548,a6512,na17918,na17920,na17922,na17924,a15314,a6522,a6566,a6608,a6494,a18026,
na18028,na6410,na6404,a6424,a6448,a18098,z0,a19208,a19248,a19262,a19274,a19282,a19292,a19300,a19308,
a19318,a19326,a19334,a19342,a19348,a19354,a19360,a19336,na16352,na19362,a6346,a19364,a19924,a19912,a19834,
a19808,a19770,a19732,a19698,a19664,a19630,a19926,a19938,a19944,a19950,a19956,a19962,a19968,a19974,a19980,
a19986,a19992,a16070,a20004,a20010,a20016,a20022,a20028,a20034,a20040,a20046,a20052,a20058,a20060,a20072,
a20078,a20084,a20090,a20096,a20102,a20108,a20114,a20120,a20126,a20128,a20140,a20146,a20152,a20158,a20164,
a20170,a20176,a20182,a20188,a20194,a20196,a20208,a20214,a20220,a20226,a20232,a20238,a20244,a20250,a20256,
a20262,a20264,a20276,a20282,a20288,a20294,a20300,a20306,a20312,a20318,a20324,a20330,a20332,a20344,a20350,
a20356,a20362,a20368,a20374,a20380,a20386,a20392,a20398,a8042,a20412,a20418,a20424,a20430,a20436,a20442,
a20448,a20454,a20460,a20466,a20564,a20636,a20666,a20716,a20762,a20800,a20816,a20836,a20854,a20870,na20872,
na20874,na20876,na20878,a6384,a6372,a6362,a6394,a19886,a19494,a20898,na21812,a22630,na6674,z1,a22638,
a22656,a22664,a22668,a22670,a22676,z2,na11396,z3,z4,z5,z6,a15296,a22688,a22696,a22706,
a22712,a22686,a24442,a24660,a26604,a26614,a26616,a26622,a10920,a10962,a10816,a10876,a27060,a11278,a22600,
a15956,a22172,a27108,a15858,a22230,a27156,a15760,a22288,a27204,a15656,a22346,a27252,a15552,a22404,a27300,
a15448,a22462,a27348,a27382,a11380,a22520,a27398,a27414,a27430,a11040,a27454,a27460,a27466,a27472,a27478,
a27484,a27490,a27498,a28230,a28254,a28004,a28082,a28278,a28302,a27902,a27890,a27802,a27790,a27698,a27684,
a27588,a27572,a28314,a28320,a28326,a28332,a28338,a28344,a28350,a28356,a28362,a28368,a24820,a24812,a24792,
a24784,a24772,a24764,a24748,a24740,a24728,a24720,na26802,a28380,a28386,a28392,a28398,a28404,a28410,a28416,
a28422,a28428,a28434,a25690,a25682,a25662,a25654,a25642,a25634,a25618,a25610,a25598,a25590,na26780,a28446,
a28452,a28458,a28464,a28470,a28476,a28482,a28488,a28494,a28500,a25566,a25558,a25538,a25530,a25518,a25510,
a25494,a25486,a25474,a25466,na26752,a28512,a28518,a28524,a28530,a28536,a28542,a28548,a28554,a28560,a28566,
a25442,a25434,a25414,a25406,a25394,a25386,a25370,a25362,a25350,a25342,na26724,a28578,a28584,a28590,a28596,
a28602,a28608,a28614,a28620,a28626,a28632,a25318,a25310,a25290,a25282,a25270,a25262,a25246,a25238,a25226,
a25218,na26696,a28644,a28650,a28656,a28662,a28668,a28674,a28680,a28686,a28692,a28698,a25194,a25186,a25166,
a25158,a25146,a25138,a25122,a25114,a25102,a25094,na26668,a28710,a28716,a28722,a28728,a28734,a28740,a28746,
a28752,a28758,a28764,a25070,a25062,a25042,a25034,a25022,a25014,a24998,a24990,a24978,a24970,a26636,a28776,
a28782,a28788,a28794,a28800,a28806,a28812,a28818,a28824,a28830,a24946,a24938,a24918,a24910,a24898,a24890,
a24874,a24866,a24854,a24846,a22946,a22778,a22806,a22834,a22862,a22890,a22918,a22750,a28834,na28842,na28854,
a28866,a28878,z7,a28882,a28888,a28894,a28900,a28906,a28912,a28918,a28924,a21698,na24508,na1690,z8,
a28938,a28942,a28972,a17616,a29058,a29072,a29084,a29096,a17748,a17488,a17350,a17216,a17082,a16950,a16808,
a16674,a16356,a29102,a29108,a29114,a29120,a28072,a29122,a27972,a27938,a27872,a27838,a27768,a27734,a27664,
a27630,a29132,a27452,na27436,a29144,a29154,a29160,a19484,a19474,a19510,a19518,a19526,a19534,a29170,a29180,
a29190,a29200,a29210,a29220,a29230,a29240,na29242,a29340,z9,a29390,a29408,a29426,a29440,a30318,a30352,
na30354,na30356,na30358,a30366,na2330,na2332,na2336,a30384,na30386,a30392,na2334,a30410,a30416,a30428,a30434,
a30468,a30482,a30490,a30496,a30506,a32028,a32548,na32550,a29254,na32552,a29248,na32554,a29262,na32556,a29270,
na32562,na15294,a32564,c1,a1688,a1690,a1692,a1694,a1696,a1698,a1700,a1702,a1704,a1706,a1708,
a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,a1732,a1734,a1736,a1738,
a1740,a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,a1758,a1760,a1762,a1764,a1766,a1768,
a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,a1790,a1792,a1794,a1796,a1798,
a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,a1822,a1824,a1826,a1828,
a1830,a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,a1848,a1850,a1852,a1854,a1856,a1858,
a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,a1882,a1884,a1886,a1888,
a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,a1910,a1912,a1914,a1916,a1918,
a1920,a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,a1938,a1940,a1942,a1944,a1946,a1948,
a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,a1972,a1974,a1976,a1978,
a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,a1998,a2000,a2002,a2004,a2006,a2008,
a2010,a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,a2030,a2032,a2034,a2036,a2038,
a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,a2058,a2060,a2062,a2064,a2066,a2068,
a2070,a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,a2090,a2092,a2094,a2096,a2098,
a2100,a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,a2120,a2122,a2124,a2126,a2128,
a2130,a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,a2152,a2154,a2156,a2158,
a2160,a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,a2178,a2180,a2182,a2184,a2186,a2188,
a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,a2208,a2210,a2212,a2214,a2216,a2218,
a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,a2238,a2240,a2242,a2244,a2246,a2248,
a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,a2268,a2270,a2272,a2274,a2276,a2278,
a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,a2298,a2300,a2302,a2304,a2306,a2308,
a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,a2328,a2330,a2332,a2334,a2336,a2338,
a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,a2358,a2360,a2362,a2364,a2366,a2368,
a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,a2388,a2390,a2392,a2394,a2396,a2398,
a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,a2420,a2422,a2424,a2426,a2428,
a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,a2448,a2450,a2452,a2454,a2456,a2458,
a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,a2478,a2480,a2482,a2484,a2486,a2488,
a2490,a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,a2508,a2510,a2512,a2514,a2516,a2518,
a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,a2540,a2542,a2544,a2546,a2548,
a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,a2572,a2574,a2576,a2578,
a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,a2602,a2604,a2606,a2608,
a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,a2630,a2632,a2634,a2636,a2638,
a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,a2662,a2664,a2666,a2668,
a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,a2692,a2694,a2696,a2698,
a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,a2718,a2720,a2722,a2724,a2726,a2728,
a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,a2752,a2754,a2756,a2758,
a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,a2782,a2784,a2786,a2788,
a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,a2810,a2812,a2814,a2816,a2818,
a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,a2840,a2842,a2844,a2846,a2848,
a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,a2870,a2872,a2874,a2876,a2878,
a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,a2900,a2902,a2904,a2906,a2908,
a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2930,a2932,a2934,a2936,a2938,
a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,a2960,a2962,a2964,a2966,a2968,
a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,a2988,a2990,a2992,a2994,a2996,a2998,
a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,a3022,a3024,a3026,a3028,
a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,a3048,a3050,a3052,a3054,a3056,a3058,
a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,a3078,a3080,a3082,a3084,a3086,a3088,
a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,a3112,a3114,a3116,a3118,
a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,a3142,a3144,a3146,a3148,
a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,a3172,a3174,a3176,a3178,
a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3200,a3202,a3204,a3206,a3208,
a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,a3228,a3230,a3232,a3234,a3236,a3238,
a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,a3262,a3264,a3266,a3268,
a3270,a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,a3288,a3290,a3292,a3294,a3296,a3298,
a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,a3324,a3326,a3328,
a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,a3354,a3356,a3358,
a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3382,a3384,a3386,a3388,
a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,a3408,a3410,a3412,a3414,a3416,a3418,
a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,a3438,a3440,a3442,a3444,a3446,a3448,
a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,a3468,a3470,a3472,a3474,a3476,a3478,
a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,a3498,a3500,a3502,a3504,a3506,a3508,
a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,a3528,a3530,a3532,a3534,a3536,a3538,
a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,a3558,a3560,a3562,a3564,a3566,a3568,
a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,a3588,a3590,a3592,a3594,a3596,a3598,
a3600,a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,a3618,a3620,a3622,a3624,a3626,a3628,
a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3648,a3650,a3652,a3654,a3656,a3658,
a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,a3678,a3680,a3682,a3684,a3686,a3688,
a3690,a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,a3712,a3714,a3716,a3718,
a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,a3738,a3740,a3742,a3744,a3746,a3748,
a3750,a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,a3768,a3770,a3772,a3774,a3776,a3778,
a3780,a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,a3798,a3800,a3802,a3804,a3806,a3808,
a3810,a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,a3828,a3830,a3832,a3834,a3836,a3838,
a3840,a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,a3858,a3860,a3862,a3864,a3866,a3868,
a3870,a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,a3888,a3890,a3892,a3894,a3896,a3898,
a3900,a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,a3918,a3920,a3922,a3924,a3926,a3928,
a3930,a3932,a3934,a3936,a3938,a3940,a3942,a3944,a3946,a3948,a3950,a3952,a3954,a3956,a3958,
a3960,a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,a3978,a3980,a3982,a3984,a3986,a3988,
a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,a4008,a4010,a4012,a4014,a4016,a4018,
a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,a4038,a4040,a4042,a4044,a4046,a4048,
a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,a4068,a4070,a4072,a4074,a4076,a4078,
a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,a4096,a4098,a4100,a4102,a4104,a4106,a4108,
a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4124,a4126,a4128,a4130,a4132,a4134,a4136,a4138,
a4140,a4142,a4144,a4146,a4148,a4150,a4152,a4154,a4156,a4158,a4160,a4162,a4164,a4166,a4168,
a4170,a4172,a4174,a4176,a4178,a4180,a4182,a4184,a4186,a4188,a4190,a4192,a4194,a4196,a4198,
a4200,a4202,a4204,a4206,a4208,a4210,a4212,a4214,a4216,a4218,a4220,a4222,a4224,a4226,a4228,
a4230,a4232,a4234,a4236,a4238,a4240,a4242,a4244,a4246,a4248,a4250,a4252,a4254,a4256,a4258,
a4260,a4262,a4264,a4266,a4268,a4270,a4272,a4274,a4276,a4278,a4280,a4282,a4284,a4286,a4288,
a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,a4306,a4308,a4310,a4312,a4314,a4316,a4318,
a4320,a4322,a4324,a4326,a4328,a4330,a4332,a4334,a4336,a4338,a4340,a4342,a4344,a4346,a4348,
a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,a4368,a4370,a4372,a4374,a4376,a4378,
a4380,a4382,a4384,a4386,a4388,a4390,a4392,a4394,a4396,a4398,a4400,a4402,a4404,a4406,a4408,
a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,a4432,a4434,a4436,a4438,
a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,a4458,a4460,a4462,a4464,a4466,a4468,
a4470,a4472,a4474,a4476,a4478,a4480,a4482,a4484,a4486,a4488,a4490,a4492,a4494,a4496,a4498,
a4500,a4502,a4504,a4506,a4508,a4510,a4512,a4514,a4516,a4518,a4520,a4522,a4524,a4526,a4528,
a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,a4554,a4556,a4558,
a4560,a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,a4578,a4580,a4582,a4584,a4586,a4588,
a4590,a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,a4612,a4614,a4616,a4618,
a4620,a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,a4642,a4644,a4646,a4648,
a4650,a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,a4672,a4674,a4676,a4678,
a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,a4696,a4698,a4700,a4702,a4704,a4706,a4708,
a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,a4726,a4728,a4730,a4732,a4734,a4736,a4738,
a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,a4756,a4758,a4760,a4762,a4764,a4766,a4768,
a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4784,a4786,a4788,a4790,a4792,a4794,a4796,a4798,
a4800,a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,a4818,a4820,a4822,a4824,a4826,a4828,
a4830,a4832,a4834,a4836,a4838,a4840,a4842,a4844,a4846,a4848,a4850,a4852,a4854,a4856,a4858,
a4860,a4862,a4864,a4866,a4868,a4870,a4872,a4874,a4876,a4878,a4880,a4882,a4884,a4886,a4888,
a4890,a4892,a4894,a4896,a4898,a4900,a4902,a4904,a4906,a4908,a4910,a4912,a4914,a4916,a4918,
a4920,a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,a4938,a4940,a4942,a4944,a4946,a4948,
a4950,a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,a4968,a4970,a4972,a4974,a4976,a4978,
a4980,a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,a4998,a5000,a5002,a5004,a5006,a5008,
a5010,a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,a5028,a5030,a5032,a5034,a5036,a5038,
a5040,a5042,a5044,a5046,a5048,a5050,a5052,a5054,a5056,a5058,a5060,a5062,a5064,a5066,a5068,
a5070,a5072,a5074,a5076,a5078,a5080,a5082,a5084,a5086,a5088,a5090,a5092,a5094,a5096,a5098,
a5100,a5102,a5104,a5106,a5108,a5110,a5112,a5114,a5116,a5118,a5120,a5122,a5124,a5126,a5128,
a5130,a5132,a5134,a5136,a5138,a5140,a5142,a5144,a5146,a5148,a5150,a5152,a5154,a5156,a5158,
a5160,a5162,a5164,a5166,a5168,a5170,a5172,a5174,a5176,a5178,a5180,a5182,a5184,a5186,a5188,
a5190,a5192,a5194,a5196,a5198,a5200,a5202,a5204,a5206,a5208,a5210,a5212,a5214,a5216,a5218,
a5220,a5222,a5224,a5226,a5228,a5230,a5232,a5234,a5236,a5238,a5240,a5242,a5244,a5246,a5248,
a5250,a5252,a5254,a5256,a5258,a5260,a5262,a5264,a5266,a5268,a5270,a5272,a5274,a5276,a5278,
a5280,a5282,a5284,a5286,a5288,a5290,a5292,a5294,a5296,a5298,a5300,a5302,a5304,a5306,a5308,
a5310,a5312,a5314,a5316,a5318,a5320,a5322,a5324,a5326,a5328,a5330,a5332,a5334,a5336,a5338,
a5340,a5342,a5344,a5346,a5348,a5350,a5352,a5354,a5356,a5358,a5360,a5362,a5364,a5366,a5368,
a5370,a5372,a5374,a5376,a5378,a5380,a5382,a5384,a5386,a5388,a5390,a5392,a5394,a5396,a5398,
a5400,a5402,a5404,a5406,a5408,a5410,a5412,a5414,a5416,a5418,a5420,a5422,a5424,a5426,a5428,
a5430,a5432,a5434,a5436,a5438,a5440,a5442,a5444,a5446,a5448,a5450,a5452,a5454,a5456,a5458,
a5460,a5462,a5464,a5466,a5468,a5470,a5472,a5474,a5476,a5478,a5480,a5482,a5484,a5486,a5488,
a5490,a5492,a5494,a5496,a5498,a5500,a5502,a5504,a5506,a5508,a5510,a5512,a5514,a5516,a5518,
a5520,a5522,a5524,a5526,a5528,a5530,a5532,a5534,a5536,a5538,a5540,a5542,a5544,a5546,a5548,
a5550,a5552,a5554,a5556,a5558,a5560,a5562,a5564,a5566,a5568,a5570,a5572,a5574,a5576,a5578,
a5580,a5582,a5584,a5586,a5588,a5590,a5592,a5594,a5596,a5598,a5600,a5602,a5604,a5606,a5608,
a5610,a5612,a5614,a5616,a5618,a5620,a5622,a5624,a5626,a5628,a5630,a5632,a5634,a5636,a5638,
a5640,a5642,a5644,a5646,a5648,a5650,a5652,a5654,a5656,a5658,a5660,a5662,a5664,a5666,a5668,
a5670,a5672,a5674,a5676,a5678,a5680,a5682,a5684,a5686,a5688,a5690,a5692,a5694,a5696,a5698,
a5700,a5702,a5704,a5706,a5708,a5710,a5712,a5714,a5716,a5718,a5720,a5722,a5724,a5726,a5728,
a5730,a5732,a5734,a5736,a5738,a5740,a5742,a5744,a5746,a5748,a5750,a5752,a5754,a5756,a5758,
a5760,a5762,a5764,a5766,a5768,a5770,a5772,a5774,a5776,a5778,a5780,a5782,a5784,a5786,a5788,
a5790,a5792,a5794,a5796,a5798,a5800,a5802,a5804,a5806,a5808,a5810,a5812,a5814,a5816,a5818,
a5820,a5822,a5824,a5826,a5828,a5830,a5832,a5834,a5836,a5838,a5840,a5842,a5844,a5846,a5848,
a5850,a5852,a5854,a5856,a5858,a5860,a5862,a5864,a5866,a5868,a5870,a5872,a5874,a5876,a5878,
a5880,a5882,a5884,a5886,a5888,a5890,a5892,a5894,a5896,a5898,a5900,a5902,a5904,a5906,a5908,
a5910,a5912,a5914,a5916,a5918,a5920,a5922,a5924,a5926,a5928,a5930,a5932,a5934,a5936,a5938,
a5940,a5942,a5944,a5946,a5948,a5950,a5952,a5954,a5956,a5958,a5960,a5962,a5964,a5966,a5968,
a5970,a5972,a5974,a5976,a5978,a5980,a5982,a5984,a5986,a5988,a5990,a5992,a5994,a5996,a5998,
a6000,a6002,a6004,a6006,a6008,a6010,a6012,a6014,a6016,a6018,a6020,a6022,a6024,a6026,a6028,
a6030,a6032,a6034,a6036,a6038,a6040,a6042,a6044,a6046,a6048,a6050,a6052,a6054,a6056,a6058,
a6060,a6062,a6064,a6066,a6068,a6070,a6072,a6076,a6078,a6080,a6082,a6084,a6086,a6088,a6090,
a6092,a6094,a6096,a6098,a6100,a6102,a6104,a6106,a6108,a6110,a6112,a6114,a6116,a6118,a6120,
a6122,a6124,a6126,a6128,a6130,a6132,a6134,a6136,a6138,a6140,a6142,a6144,a6146,a6148,a6150,
a6152,a6154,a6156,a6158,a6160,a6162,a6164,a6166,a6168,a6170,a6172,a6174,a6176,a6178,a6180,
a6182,a6184,a6186,a6188,a6190,a6192,a6194,a6196,a6198,a6200,a6202,a6204,a6206,a6208,a6210,
a6212,a6214,a6216,a6218,a6220,a6222,a6224,a6226,a6228,a6230,a6232,a6234,a6236,a6238,a6240,
a6242,a6244,a6246,a6248,a6250,a6252,a6254,a6256,a6258,a6260,a6262,a6264,a6266,a6268,a6270,
a6272,a6274,a6276,a6278,a6280,a6282,a6284,a6286,a6288,a6290,a6292,a6294,a6296,a6298,a6300,
a6302,a6304,a6306,a6308,a6310,a6312,a6314,a6316,a6318,a6320,a6322,a6324,a6326,a6328,a6330,
a6332,a6334,a6336,a6338,a6340,a6342,a6344,a6348,a6350,a6352,a6354,a6356,a6358,a6360,a6364,
a6366,a6368,a6370,a6374,a6376,a6378,a6380,a6382,a6386,a6388,a6390,a6392,a6396,a6398,a6400,
a6402,a6404,a6406,a6408,a6410,a6412,a6414,a6416,a6418,a6420,a6422,a6426,a6428,a6430,a6432,
a6434,a6436,a6438,a6440,a6442,a6444,a6446,a6450,a6452,a6454,a6456,a6458,a6460,a6462,a6464,
a6466,a6468,a6470,a6472,a6474,a6478,a6480,a6482,a6484,a6486,a6488,a6490,a6492,a6496,a6498,
a6500,a6502,a6504,a6506,a6508,a6510,a6514,a6516,a6518,a6520,a6524,a6526,a6528,a6530,a6532,
a6534,a6536,a6538,a6540,a6542,a6544,a6546,a6550,a6552,a6554,a6556,a6558,a6560,a6562,a6564,
a6568,a6570,a6572,a6574,a6576,a6578,a6580,a6582,a6584,a6586,a6588,a6590,a6594,a6596,a6598,
a6600,a6602,a6604,a6606,a6610,a6612,a6614,a6616,a6618,a6620,a6622,a6624,a6626,a6628,a6630,
a6632,a6634,a6636,a6638,a6640,a6642,a6644,a6646,a6648,a6650,a6652,a6654,a6656,a6658,a6660,
a6664,a6666,a6668,a6670,a6672,a6674,a6676,a6678,a6680,a6684,a6686,a6688,a6692,a6694,a6698,
a6700,a6704,a6706,a6710,a6714,a6716,a6718,a6720,a6722,a6724,a6726,a6728,a6730,a6732,a6734,
a6736,a6738,a6740,a6742,a6744,a6746,a6748,a6750,a6752,a6754,a6756,a6758,a6760,a6762,a6764,
a6766,a6768,a6770,a6772,a6774,a6776,a6778,a6780,a6782,a6784,a6786,a6788,a6790,a6792,a6794,
a6796,a6798,a6800,a6802,a6804,a6806,a6808,a6810,a6812,a6814,a6816,a6818,a6820,a6822,a6824,
a6826,a6828,a6830,a6832,a6834,a6836,a6838,a6840,a6842,a6844,a6846,a6848,a6850,a6852,a6854,
a6856,a6858,a6860,a6862,a6864,a6866,a6868,a6870,a6872,a6874,a6876,a6878,a6880,a6882,a6884,
a6886,a6888,a6890,a6892,a6894,a6896,a6898,a6900,a6902,a6904,a6906,a6908,a6910,a6912,a6914,
a6916,a6918,a6922,a6924,a6926,a6928,a6930,a6932,a6934,a6936,a6938,a6940,a6942,a6944,a6946,
a6948,a6950,a6952,a6954,a6956,a6958,a6960,a6962,a6964,a6966,a6968,a6970,a6972,a6974,a6976,
a6978,a6980,a6982,a6984,a6986,a6988,a6990,a6992,a6994,a6996,a6998,a7000,a7002,a7004,a7006,
a7008,a7010,a7012,a7014,a7016,a7018,a7020,a7022,a7024,a7026,a7028,a7030,a7032,a7034,a7036,
a7038,a7040,a7042,a7044,a7046,a7048,a7050,a7052,a7054,a7056,a7058,a7060,a7062,a7064,a7066,
a7068,a7070,a7072,a7074,a7076,a7078,a7080,a7082,a7084,a7086,a7088,a7090,a7092,a7094,a7096,
a7098,a7100,a7102,a7104,a7106,a7108,a7110,a7112,a7114,a7116,a7118,a7120,a7122,a7124,a7126,
a7128,a7130,a7132,a7134,a7136,a7138,a7140,a7142,a7144,a7146,a7148,a7150,a7154,a7156,a7158,
a7160,a7162,a7164,a7166,a7168,a7170,a7172,a7174,a7176,a7178,a7180,a7182,a7184,a7186,a7188,
a7190,a7192,a7194,a7196,a7198,a7200,a7202,a7204,a7206,a7208,a7210,a7212,a7214,a7216,a7218,
a7220,a7222,a7224,a7226,a7228,a7230,a7232,a7234,a7236,a7238,a7240,a7242,a7244,a7246,a7248,
a7250,a7252,a7254,a7256,a7258,a7260,a7262,a7264,a7266,a7268,a7270,a7272,a7274,a7276,a7278,
a7280,a7282,a7284,a7286,a7288,a7290,a7292,a7294,a7296,a7298,a7300,a7302,a7304,a7306,a7308,
a7310,a7312,a7314,a7316,a7318,a7320,a7322,a7324,a7326,a7328,a7330,a7332,a7334,a7336,a7338,
a7340,a7342,a7344,a7346,a7348,a7350,a7354,a7356,a7358,a7360,a7362,a7364,a7366,a7368,a7370,
a7372,a7374,a7376,a7378,a7380,a7382,a7384,a7386,a7388,a7390,a7392,a7394,a7396,a7398,a7400,
a7402,a7404,a7406,a7408,a7410,a7412,a7414,a7416,a7418,a7420,a7422,a7424,a7426,a7428,a7430,
a7432,a7434,a7436,a7438,a7440,a7442,a7444,a7446,a7448,a7450,a7452,a7454,a7456,a7458,a7460,
a7462,a7464,a7466,a7468,a7470,a7472,a7474,a7476,a7478,a7480,a7482,a7484,a7486,a7488,a7490,
a7492,a7494,a7496,a7498,a7500,a7502,a7504,a7506,a7508,a7510,a7512,a7514,a7516,a7518,a7520,
a7522,a7524,a7526,a7528,a7530,a7532,a7534,a7536,a7538,a7540,a7542,a7544,a7546,a7548,a7550,
a7552,a7554,a7556,a7558,a7560,a7562,a7564,a7566,a7568,a7570,a7572,a7574,a7576,a7578,a7580,
a7582,a7584,a7586,a7588,a7592,a7594,a7596,a7598,a7600,a7602,a7604,a7606,a7608,a7610,a7612,
a7614,a7616,a7618,a7620,a7622,a7624,a7626,a7628,a7630,a7632,a7634,a7636,a7638,a7640,a7642,
a7644,a7646,a7648,a7650,a7652,a7654,a7656,a7658,a7660,a7662,a7664,a7666,a7668,a7670,a7672,
a7674,a7676,a7678,a7680,a7682,a7684,a7686,a7688,a7690,a7692,a7694,a7696,a7698,a7700,a7702,
a7704,a7706,a7708,a7710,a7712,a7714,a7716,a7718,a7720,a7722,a7724,a7726,a7728,a7730,a7732,
a7734,a7736,a7738,a7740,a7742,a7744,a7746,a7748,a7750,a7752,a7754,a7756,a7758,a7760,a7762,
a7764,a7766,a7768,a7770,a7772,a7774,a7776,a7778,a7780,a7782,a7784,a7786,a7788,a7790,a7792,
a7794,a7796,a7798,a7800,a7802,a7804,a7806,a7808,a7810,a7814,a7816,a7818,a7820,a7822,a7824,
a7826,a7828,a7830,a7832,a7834,a7836,a7838,a7840,a7842,a7844,a7846,a7848,a7850,a7854,a7856,
a7858,a7860,a7862,a7866,a7868,a7870,a7872,a7874,a7876,a7878,a7880,a7882,a7884,a7886,a7888,
a7890,a7892,a7894,a7896,a7898,a7902,a7904,a7906,a7908,a7910,a7912,a7914,a7916,a7918,a7920,
a7922,a7924,a7926,a7928,a7932,a7934,a7936,a7938,a7940,a7944,a7946,a7948,a7950,a7952,a7956,
a7958,a7960,a7962,a7964,a7968,a7970,a7972,a7974,a7976,a7980,a7982,a7984,a7986,a7988,a7992,
a7994,a7996,a7998,a8000,a8004,a8006,a8008,a8010,a8012,a8014,a8016,a8018,a8022,a8024,a8026,
a8028,a8030,a8032,a8034,a8036,a8038,a8040,a8044,a8046,a8048,a8050,a8052,a8054,a8056,a8058,
a8060,a8062,a8064,a8066,a8068,a8070,a8072,a8074,a8076,a8078,a8080,a8082,a8084,a8086,a8088,
a8090,a8092,a8094,a8096,a8098,a8100,a8102,a8104,a8106,a8108,a8110,a8112,a8114,a8116,a8118,
a8120,a8122,a8124,a8126,a8128,a8130,a8132,a8134,a8136,a8138,a8140,a8142,a8144,a8146,a8148,
a8150,a8152,a8154,a8156,a8158,a8160,a8162,a8164,a8166,a8168,a8170,a8172,a8174,a8176,a8178,
a8180,a8182,a8184,a8186,a8188,a8190,a8192,a8194,a8196,a8198,a8200,a8202,a8204,a8206,a8208,
a8210,a8212,a8214,a8216,a8218,a8220,a8222,a8224,a8226,a8228,a8230,a8232,a8234,a8236,a8238,
a8240,a8242,a8244,a8246,a8248,a8250,a8252,a8254,a8256,a8258,a8260,a8262,a8264,a8266,a8268,
a8270,a8272,a8274,a8276,a8278,a8280,a8282,a8284,a8286,a8288,a8290,a8292,a8294,a8296,a8298,
a8300,a8302,a8304,a8306,a8308,a8310,a8312,a8314,a8316,a8318,a8320,a8322,a8324,a8326,a8328,
a8330,a8332,a8334,a8336,a8338,a8340,a8342,a8344,a8346,a8348,a8350,a8352,a8354,a8356,a8358,
a8360,a8362,a8364,a8366,a8368,a8370,a8372,a8374,a8376,a8378,a8380,a8382,a8384,a8386,a8388,
a8390,a8392,a8394,a8396,a8398,a8400,a8402,a8404,a8406,a8408,a8410,a8412,a8414,a8416,a8418,
a8420,a8422,a8424,a8426,a8428,a8430,a8432,a8434,a8436,a8438,a8440,a8442,a8444,a8446,a8448,
a8450,a8452,a8454,a8456,a8458,a8460,a8462,a8464,a8466,a8468,a8470,a8472,a8474,a8476,a8478,
a8480,a8482,a8484,a8486,a8488,a8490,a8492,a8494,a8496,a8498,a8500,a8502,a8504,a8506,a8508,
a8510,a8512,a8514,a8516,a8518,a8520,a8522,a8524,a8526,a8528,a8530,a8532,a8534,a8536,a8538,
a8540,a8542,a8544,a8546,a8548,a8550,a8552,a8554,a8556,a8558,a8560,a8562,a8564,a8566,a8568,
a8570,a8572,a8574,a8576,a8578,a8580,a8582,a8584,a8586,a8588,a8590,a8592,a8594,a8596,a8598,
a8600,a8602,a8604,a8606,a8608,a8610,a8612,a8614,a8616,a8618,a8620,a8622,a8624,a8626,a8628,
a8630,a8632,a8634,a8636,a8638,a8640,a8642,a8644,a8646,a8648,a8650,a8652,a8654,a8656,a8658,
a8660,a8662,a8664,a8666,a8668,a8670,a8672,a8674,a8676,a8678,a8680,a8682,a8684,a8686,a8688,
a8690,a8692,a8694,a8696,a8698,a8700,a8702,a8704,a8706,a8708,a8710,a8712,a8714,a8716,a8718,
a8720,a8722,a8724,a8726,a8728,a8730,a8732,a8734,a8736,a8738,a8740,a8742,a8744,a8746,a8748,
a8750,a8752,a8754,a8756,a8758,a8760,a8762,a8764,a8766,a8768,a8770,a8772,a8774,a8776,a8778,
a8780,a8782,a8784,a8786,a8788,a8790,a8792,a8794,a8796,a8798,a8800,a8802,a8804,a8806,a8808,
a8810,a8812,a8814,a8816,a8818,a8820,a8822,a8824,a8826,a8828,a8830,a8832,a8834,a8836,a8838,
a8840,a8842,a8844,a8846,a8848,a8850,a8852,a8854,a8856,a8858,a8860,a8862,a8864,a8866,a8868,
a8870,a8872,a8874,a8876,a8878,a8880,a8882,a8884,a8886,a8888,a8890,a8892,a8894,a8896,a8898,
a8900,a8902,a8904,a8906,a8908,a8910,a8912,a8914,a8916,a8918,a8920,a8922,a8924,a8926,a8928,
a8930,a8932,a8934,a8936,a8938,a8940,a8942,a8944,a8946,a8948,a8950,a8952,a8954,a8956,a8958,
a8960,a8962,a8964,a8966,a8968,a8970,a8972,a8974,a8976,a8978,a8980,a8982,a8984,a8986,a8988,
a8990,a8992,a8994,a8996,a8998,a9000,a9002,a9004,a9006,a9008,a9010,a9012,a9014,a9016,a9018,
a9020,a9022,a9024,a9026,a9028,a9030,a9032,a9034,a9036,a9038,a9040,a9042,a9044,a9046,a9048,
a9050,a9052,a9054,a9056,a9058,a9060,a9062,a9064,a9066,a9068,a9070,a9072,a9074,a9076,a9078,
a9080,a9082,a9084,a9086,a9088,a9090,a9092,a9094,a9096,a9098,a9100,a9102,a9104,a9106,a9108,
a9110,a9112,a9114,a9116,a9118,a9120,a9122,a9124,a9126,a9128,a9130,a9132,a9134,a9136,a9138,
a9140,a9142,a9144,a9146,a9148,a9150,a9152,a9154,a9156,a9158,a9160,a9162,a9164,a9166,a9168,
a9170,a9172,a9174,a9176,a9178,a9180,a9182,a9184,a9186,a9188,a9190,a9192,a9194,a9196,a9198,
a9200,a9202,a9204,a9206,a9208,a9210,a9212,a9214,a9216,a9218,a9220,a9222,a9224,a9226,a9228,
a9230,a9232,a9234,a9236,a9238,a9240,a9242,a9244,a9246,a9248,a9250,a9252,a9254,a9256,a9258,
a9260,a9262,a9264,a9266,a9268,a9270,a9272,a9274,a9276,a9278,a9280,a9282,a9284,a9286,a9288,
a9290,a9292,a9294,a9296,a9298,a9300,a9302,a9304,a9306,a9308,a9310,a9312,a9314,a9316,a9318,
a9320,a9322,a9324,a9326,a9328,a9330,a9332,a9334,a9336,a9338,a9340,a9342,a9344,a9346,a9348,
a9350,a9352,a9354,a9356,a9358,a9360,a9362,a9364,a9366,a9368,a9370,a9372,a9374,a9376,a9378,
a9380,a9382,a9384,a9386,a9388,a9390,a9392,a9394,a9396,a9398,a9400,a9402,a9404,a9406,a9408,
a9410,a9412,a9414,a9416,a9418,a9420,a9422,a9424,a9426,a9428,a9430,a9432,a9434,a9436,a9438,
a9440,a9442,a9444,a9446,a9448,a9450,a9452,a9454,a9456,a9458,a9460,a9462,a9464,a9466,a9468,
a9470,a9472,a9474,a9476,a9478,a9480,a9482,a9484,a9486,a9488,a9490,a9492,a9494,a9496,a9498,
a9500,a9502,a9504,a9506,a9508,a9510,a9512,a9514,a9516,a9518,a9520,a9522,a9524,a9526,a9528,
a9530,a9532,a9534,a9536,a9538,a9540,a9542,a9544,a9546,a9548,a9550,a9552,a9554,a9556,a9558,
a9560,a9562,a9564,a9566,a9568,a9570,a9572,a9574,a9576,a9578,a9580,a9582,a9584,a9586,a9588,
a9590,a9592,a9594,a9596,a9598,a9600,a9602,a9604,a9606,a9608,a9610,a9612,a9614,a9616,a9618,
a9620,a9622,a9624,a9626,a9628,a9630,a9632,a9634,a9636,a9638,a9640,a9642,a9644,a9646,a9648,
a9650,a9652,a9654,a9656,a9658,a9660,a9662,a9664,a9666,a9668,a9670,a9672,a9674,a9676,a9678,
a9680,a9682,a9684,a9686,a9688,a9690,a9692,a9694,a9696,a9698,a9700,a9702,a9704,a9706,a9708,
a9710,a9712,a9714,a9716,a9718,a9720,a9722,a9724,a9726,a9728,a9730,a9732,a9734,a9736,a9738,
a9740,a9742,a9744,a9746,a9748,a9750,a9752,a9754,a9756,a9758,a9760,a9762,a9764,a9766,a9768,
a9770,a9772,a9774,a9776,a9778,a9780,a9782,a9784,a9786,a9788,a9790,a9792,a9794,a9796,a9798,
a9800,a9802,a9804,a9806,a9808,a9810,a9812,a9814,a9816,a9818,a9820,a9822,a9824,a9826,a9828,
a9830,a9832,a9834,a9836,a9838,a9840,a9842,a9844,a9846,a9848,a9850,a9852,a9854,a9856,a9858,
a9860,a9862,a9864,a9866,a9868,a9870,a9872,a9874,a9876,a9878,a9880,a9882,a9884,a9886,a9888,
a9890,a9892,a9894,a9896,a9898,a9900,a9902,a9904,a9906,a9908,a9910,a9912,a9914,a9916,a9918,
a9920,a9922,a9924,a9926,a9928,a9930,a9932,a9934,a9936,a9938,a9940,a9942,a9944,a9946,a9948,
a9950,a9952,a9954,a9956,a9958,a9960,a9962,a9964,a9966,a9968,a9970,a9972,a9974,a9976,a9978,
a9980,a9982,a9984,a9986,a9988,a9990,a9992,a9994,a9996,a9998,a10000,a10002,a10004,a10006,a10008,
a10010,a10012,a10014,a10016,a10018,a10020,a10022,a10024,a10026,a10028,a10030,a10032,a10034,a10036,a10038,
a10040,a10042,a10044,a10046,a10048,a10050,a10052,a10054,a10056,a10058,a10060,a10062,a10064,a10066,a10068,
a10070,a10072,a10074,a10076,a10078,a10080,a10082,a10084,a10086,a10088,a10090,a10092,a10094,a10096,a10098,
a10100,a10102,a10104,a10106,a10108,a10110,a10112,a10114,a10116,a10118,a10120,a10122,a10124,a10126,a10128,
a10130,a10132,a10134,a10136,a10138,a10140,a10142,a10144,a10146,a10148,a10150,a10152,a10154,a10156,a10158,
a10160,a10162,a10164,a10166,a10168,a10170,a10172,a10174,a10176,a10178,a10180,a10182,a10184,a10186,a10188,
a10190,a10192,a10194,a10196,a10198,a10200,a10202,a10204,a10206,a10208,a10210,a10212,a10214,a10216,a10218,
a10220,a10222,a10224,a10226,a10228,a10230,a10232,a10234,a10236,a10238,a10240,a10242,a10244,a10246,a10248,
a10250,a10252,a10254,a10256,a10258,a10260,a10262,a10264,a10266,a10268,a10270,a10272,a10274,a10276,a10278,
a10280,a10282,a10284,a10286,a10288,a10290,a10292,a10294,a10296,a10298,a10300,a10302,a10304,a10306,a10308,
a10310,a10312,a10314,a10316,a10318,a10320,a10322,a10324,a10326,a10328,a10330,a10332,a10334,a10336,a10338,
a10340,a10342,a10344,a10346,a10348,a10350,a10352,a10354,a10356,a10358,a10360,a10362,a10364,a10366,a10368,
a10370,a10372,a10374,a10376,a10378,a10380,a10382,a10384,a10386,a10388,a10390,a10392,a10394,a10396,a10398,
a10400,a10402,a10404,a10406,a10408,a10410,a10412,a10414,a10416,a10418,a10420,a10422,a10424,a10426,a10428,
a10430,a10432,a10434,a10436,a10438,a10440,a10442,a10444,a10446,a10448,a10450,a10452,a10454,a10456,a10458,
a10460,a10462,a10464,a10466,a10468,a10470,a10472,a10474,a10476,a10478,a10480,a10482,a10484,a10486,a10488,
a10490,a10492,a10494,a10496,a10498,a10500,a10502,a10504,a10506,a10508,a10510,a10512,a10514,a10516,a10518,
a10520,a10522,a10524,a10526,a10528,a10530,a10532,a10534,a10536,a10538,a10540,a10542,a10544,a10546,a10548,
a10550,a10552,a10554,a10556,a10558,a10560,a10562,a10564,a10566,a10568,a10570,a10572,a10574,a10576,a10578,
a10580,a10582,a10584,a10586,a10588,a10590,a10592,a10594,a10596,a10598,a10600,a10602,a10604,a10606,a10608,
a10610,a10612,a10614,a10616,a10618,a10620,a10622,a10624,a10626,a10628,a10630,a10632,a10634,a10636,a10638,
a10640,a10642,a10644,a10646,a10648,a10650,a10652,a10654,a10656,a10658,a10660,a10662,a10664,a10666,a10668,
a10670,a10672,a10674,a10676,a10678,a10680,a10682,a10684,a10686,a10688,a10690,a10692,a10694,a10696,a10698,
a10700,a10702,a10704,a10706,a10708,a10710,a10712,a10714,a10716,a10718,a10720,a10722,a10724,a10726,a10728,
a10730,a10732,a10734,a10736,a10738,a10740,a10742,a10744,a10746,a10748,a10750,a10752,a10754,a10756,a10758,
a10760,a10762,a10764,a10766,a10768,a10770,a10772,a10774,a10776,a10778,a10780,a10782,a10784,a10786,a10788,
a10790,a10792,a10794,a10796,a10798,a10800,a10802,a10804,a10806,a10808,a10810,a10812,a10814,a10818,a10820,
a10822,a10824,a10826,a10828,a10830,a10832,a10834,a10836,a10838,a10840,a10842,a10844,a10846,a10848,a10850,
a10852,a10854,a10856,a10858,a10860,a10862,a10864,a10866,a10868,a10870,a10872,a10874,a10878,a10880,a10882,
a10884,a10886,a10888,a10890,a10892,a10894,a10896,a10898,a10900,a10902,a10904,a10906,a10908,a10910,a10912,
a10914,a10916,a10918,a10922,a10924,a10926,a10928,a10930,a10932,a10934,a10936,a10938,a10940,a10942,a10944,
a10946,a10948,a10950,a10952,a10954,a10956,a10958,a10960,a10964,a10966,a10968,a10970,a10972,a10974,a10976,
a10978,a10980,a10982,a10984,a10986,a10988,a10990,a10992,a10994,a10996,a10998,a11000,a11002,a11004,a11006,
a11008,a11010,a11012,a11014,a11016,a11018,a11020,a11022,a11024,a11026,a11028,a11030,a11032,a11034,a11036,
a11038,a11042,a11044,a11046,a11048,a11050,a11052,a11054,a11056,a11058,a11060,a11062,a11064,a11066,a11068,
a11070,a11072,a11074,a11076,a11078,a11080,a11082,a11084,a11086,a11088,a11090,a11092,a11094,a11096,a11098,
a11100,a11102,a11104,a11106,a11108,a11110,a11112,a11114,a11116,a11118,a11120,a11122,a11124,a11126,a11128,
a11130,a11132,a11134,a11136,a11138,a11140,a11142,a11144,a11146,a11148,a11150,a11152,a11154,a11156,a11158,
a11160,a11162,a11164,a11166,a11168,a11170,a11172,a11174,a11176,a11178,a11180,a11182,a11184,a11186,a11188,
a11190,a11192,a11194,a11196,a11198,a11200,a11202,a11204,a11206,a11208,a11210,a11212,a11214,a11216,a11218,
a11220,a11222,a11224,a11226,a11228,a11230,a11232,a11234,a11236,a11238,a11240,a11242,a11244,a11246,a11248,
a11250,a11252,a11254,a11256,a11258,a11260,a11262,a11264,a11266,a11268,a11270,a11272,a11274,a11276,a11280,
a11282,a11284,a11286,a11288,a11290,a11292,a11294,a11296,a11298,a11300,a11302,a11304,a11306,a11308,a11310,
a11312,a11314,a11316,a11318,a11320,a11322,a11324,a11326,a11328,a11330,a11332,a11334,a11336,a11338,a11340,
a11342,a11344,a11346,a11348,a11350,a11352,a11354,a11356,a11358,a11360,a11362,a11364,a11366,a11368,a11370,
a11372,a11374,a11376,a11378,a11382,a11384,a11386,a11388,a11390,a11392,a11394,a11396,a11398,a11400,a11402,
a11404,a11406,a11408,a11410,a11412,a11414,a11416,a11418,a11420,a11422,a11424,a11426,a11428,a11430,a11432,
a11434,a11436,a11438,a11440,a11442,a11444,a11446,a11448,a11450,a11452,a11454,a11456,a11458,a11460,a11462,
a11464,a11466,a11468,a11470,a11472,a11474,a11476,a11478,a11480,a11482,a11484,a11486,a11488,a11490,a11492,
a11494,a11496,a11498,a11500,a11502,a11504,a11506,a11508,a11510,a11512,a11514,a11516,a11518,a11520,a11522,
a11524,a11526,a11528,a11530,a11532,a11534,a11536,a11538,a11540,a11542,a11544,a11546,a11548,a11550,a11552,
a11554,a11556,a11558,a11560,a11562,a11564,a11566,a11568,a11570,a11572,a11574,a11576,a11578,a11580,a11582,
a11584,a11586,a11588,a11590,a11592,a11594,a11596,a11598,a11600,a11602,a11604,a11606,a11608,a11610,a11612,
a11614,a11616,a11618,a11620,a11622,a11624,a11626,a11628,a11630,a11632,a11634,a11636,a11638,a11640,a11642,
a11644,a11646,a11648,a11650,a11652,a11654,a11656,a11658,a11660,a11662,a11664,a11666,a11668,a11670,a11672,
a11674,a11676,a11678,a11680,a11682,a11684,a11686,a11688,a11690,a11692,a11694,a11696,a11698,a11700,a11702,
a11704,a11706,a11708,a11710,a11712,a11714,a11716,a11718,a11720,a11722,a11724,a11726,a11728,a11730,a11732,
a11734,a11736,a11738,a11740,a11742,a11744,a11746,a11748,a11750,a11752,a11754,a11756,a11758,a11760,a11762,
a11764,a11766,a11768,a11770,a11772,a11774,a11776,a11778,a11780,a11782,a11784,a11786,a11788,a11790,a11792,
a11794,a11796,a11798,a11800,a11802,a11804,a11806,a11808,a11810,a11812,a11814,a11816,a11818,a11820,a11822,
a11824,a11826,a11828,a11830,a11832,a11834,a11836,a11838,a11840,a11842,a11844,a11846,a11848,a11850,a11852,
a11854,a11856,a11858,a11860,a11862,a11864,a11866,a11868,a11870,a11872,a11874,a11876,a11878,a11880,a11882,
a11884,a11886,a11888,a11890,a11892,a11894,a11896,a11898,a11900,a11902,a11904,a11906,a11908,a11910,a11912,
a11914,a11916,a11918,a11920,a11922,a11924,a11926,a11928,a11930,a11932,a11934,a11936,a11938,a11940,a11942,
a11944,a11946,a11948,a11950,a11952,a11954,a11956,a11958,a11960,a11962,a11964,a11966,a11968,a11970,a11972,
a11974,a11976,a11978,a11980,a11982,a11984,a11986,a11988,a11990,a11992,a11994,a11996,a11998,a12000,a12002,
a12004,a12006,a12008,a12010,a12012,a12014,a12016,a12018,a12020,a12022,a12024,a12026,a12028,a12030,a12032,
a12034,a12036,a12038,a12040,a12042,a12044,a12046,a12048,a12050,a12052,a12054,a12056,a12058,a12060,a12062,
a12064,a12066,a12068,a12070,a12072,a12074,a12076,a12078,a12080,a12082,a12084,a12086,a12088,a12090,a12092,
a12094,a12096,a12098,a12100,a12102,a12104,a12106,a12108,a12110,a12112,a12114,a12116,a12118,a12120,a12122,
a12124,a12126,a12128,a12130,a12132,a12134,a12136,a12138,a12140,a12142,a12144,a12146,a12148,a12150,a12152,
a12154,a12156,a12158,a12160,a12162,a12164,a12166,a12168,a12170,a12172,a12174,a12176,a12178,a12180,a12182,
a12184,a12186,a12188,a12190,a12192,a12194,a12196,a12198,a12200,a12202,a12204,a12206,a12208,a12210,a12212,
a12214,a12216,a12218,a12220,a12222,a12224,a12226,a12228,a12230,a12232,a12234,a12236,a12238,a12240,a12242,
a12244,a12246,a12248,a12250,a12252,a12254,a12256,a12258,a12260,a12262,a12264,a12266,a12268,a12270,a12272,
a12274,a12276,a12278,a12280,a12282,a12284,a12286,a12288,a12290,a12292,a12294,a12296,a12298,a12300,a12302,
a12304,a12306,a12308,a12310,a12312,a12314,a12316,a12318,a12320,a12322,a12324,a12326,a12328,a12330,a12332,
a12334,a12336,a12338,a12340,a12342,a12344,a12346,a12348,a12350,a12352,a12354,a12356,a12358,a12360,a12362,
a12364,a12366,a12368,a12370,a12372,a12374,a12376,a12378,a12380,a12382,a12384,a12386,a12388,a12390,a12392,
a12394,a12396,a12398,a12400,a12402,a12404,a12406,a12408,a12410,a12412,a12414,a12416,a12418,a12420,a12422,
a12424,a12426,a12428,a12430,a12432,a12434,a12436,a12438,a12440,a12442,a12444,a12446,a12448,a12450,a12452,
a12454,a12456,a12458,a12460,a12462,a12464,a12466,a12468,a12470,a12472,a12474,a12476,a12478,a12480,a12482,
a12484,a12486,a12488,a12490,a12492,a12494,a12496,a12498,a12500,a12502,a12504,a12506,a12508,a12510,a12512,
a12514,a12516,a12518,a12520,a12522,a12524,a12526,a12528,a12530,a12532,a12534,a12536,a12538,a12540,a12542,
a12544,a12546,a12548,a12550,a12552,a12554,a12556,a12558,a12560,a12562,a12564,a12566,a12568,a12570,a12572,
a12574,a12576,a12578,a12580,a12582,a12584,a12586,a12588,a12590,a12592,a12594,a12596,a12598,a12600,a12602,
a12604,a12606,a12608,a12610,a12612,a12614,a12616,a12618,a12620,a12622,a12624,a12626,a12628,a12630,a12632,
a12634,a12636,a12638,a12640,a12642,a12644,a12646,a12648,a12650,a12652,a12654,a12656,a12658,a12660,a12662,
a12664,a12666,a12668,a12670,a12672,a12674,a12676,a12678,a12680,a12682,a12684,a12686,a12688,a12690,a12692,
a12694,a12696,a12698,a12700,a12702,a12704,a12706,a12708,a12710,a12712,a12714,a12716,a12718,a12720,a12722,
a12724,a12726,a12728,a12730,a12732,a12734,a12736,a12738,a12740,a12742,a12744,a12746,a12748,a12750,a12752,
a12754,a12756,a12758,a12760,a12762,a12764,a12766,a12768,a12770,a12772,a12774,a12776,a12778,a12780,a12782,
a12784,a12786,a12788,a12790,a12792,a12794,a12796,a12798,a12800,a12802,a12804,a12806,a12808,a12810,a12812,
a12814,a12816,a12818,a12820,a12822,a12824,a12826,a12828,a12830,a12832,a12834,a12836,a12838,a12840,a12842,
a12844,a12846,a12848,a12850,a12852,a12854,a12856,a12858,a12860,a12862,a12864,a12866,a12868,a12870,a12872,
a12874,a12876,a12878,a12880,a12882,a12884,a12886,a12888,a12890,a12892,a12894,a12896,a12898,a12900,a12902,
a12904,a12906,a12908,a12910,a12912,a12914,a12916,a12918,a12920,a12922,a12924,a12926,a12928,a12930,a12932,
a12934,a12936,a12938,a12940,a12942,a12944,a12946,a12948,a12950,a12952,a12954,a12956,a12958,a12960,a12962,
a12964,a12966,a12968,a12970,a12972,a12974,a12976,a12978,a12980,a12982,a12984,a12986,a12988,a12990,a12992,
a12994,a12996,a12998,a13000,a13002,a13004,a13006,a13008,a13010,a13012,a13014,a13016,a13018,a13020,a13022,
a13024,a13026,a13028,a13030,a13032,a13034,a13036,a13038,a13040,a13042,a13044,a13046,a13048,a13050,a13052,
a13054,a13056,a13058,a13060,a13062,a13064,a13066,a13068,a13070,a13072,a13074,a13076,a13078,a13080,a13082,
a13084,a13086,a13088,a13090,a13092,a13094,a13096,a13098,a13100,a13102,a13104,a13106,a13108,a13110,a13112,
a13114,a13116,a13118,a13120,a13122,a13124,a13126,a13128,a13130,a13132,a13134,a13136,a13138,a13140,a13142,
a13144,a13146,a13148,a13150,a13152,a13154,a13156,a13158,a13160,a13162,a13164,a13166,a13168,a13170,a13172,
a13174,a13176,a13178,a13180,a13182,a13184,a13186,a13188,a13190,a13192,a13194,a13196,a13198,a13200,a13202,
a13204,a13206,a13208,a13210,a13212,a13214,a13216,a13218,a13220,a13222,a13224,a13226,a13228,a13230,a13232,
a13234,a13236,a13238,a13240,a13242,a13244,a13246,a13248,a13250,a13252,a13254,a13256,a13258,a13260,a13262,
a13264,a13266,a13268,a13270,a13272,a13274,a13276,a13278,a13280,a13282,a13284,a13286,a13288,a13290,a13292,
a13294,a13296,a13298,a13300,a13302,a13304,a13306,a13308,a13310,a13312,a13314,a13316,a13318,a13320,a13322,
a13324,a13326,a13328,a13330,a13332,a13334,a13336,a13338,a13340,a13342,a13344,a13346,a13348,a13350,a13352,
a13354,a13356,a13358,a13360,a13362,a13364,a13366,a13368,a13370,a13372,a13374,a13376,a13378,a13380,a13382,
a13384,a13386,a13388,a13390,a13392,a13394,a13396,a13398,a13400,a13402,a13404,a13406,a13408,a13410,a13412,
a13414,a13416,a13418,a13420,a13422,a13424,a13426,a13428,a13430,a13432,a13434,a13436,a13438,a13440,a13442,
a13444,a13446,a13448,a13450,a13452,a13454,a13456,a13458,a13460,a13462,a13464,a13466,a13468,a13470,a13472,
a13474,a13476,a13478,a13480,a13482,a13484,a13486,a13488,a13490,a13492,a13494,a13496,a13498,a13500,a13502,
a13504,a13506,a13508,a13510,a13512,a13514,a13516,a13518,a13520,a13522,a13524,a13526,a13528,a13530,a13532,
a13534,a13536,a13538,a13540,a13542,a13544,a13546,a13548,a13550,a13552,a13554,a13556,a13558,a13560,a13562,
a13564,a13566,a13568,a13570,a13572,a13574,a13576,a13578,a13580,a13582,a13584,a13586,a13588,a13590,a13592,
a13594,a13596,a13598,a13600,a13602,a13604,a13606,a13608,a13610,a13612,a13614,a13616,a13618,a13620,a13622,
a13624,a13626,a13628,a13630,a13632,a13634,a13636,a13638,a13640,a13642,a13644,a13646,a13648,a13650,a13652,
a13654,a13656,a13658,a13660,a13662,a13664,a13666,a13668,a13670,a13672,a13674,a13676,a13678,a13680,a13682,
a13684,a13686,a13688,a13690,a13692,a13694,a13696,a13698,a13700,a13702,a13704,a13706,a13708,a13710,a13712,
a13714,a13716,a13718,a13720,a13722,a13724,a13726,a13728,a13730,a13732,a13734,a13736,a13738,a13740,a13742,
a13744,a13746,a13748,a13750,a13752,a13754,a13756,a13758,a13760,a13762,a13764,a13766,a13768,a13770,a13772,
a13774,a13776,a13778,a13780,a13782,a13784,a13786,a13788,a13790,a13792,a13794,a13796,a13798,a13800,a13802,
a13804,a13806,a13808,a13810,a13812,a13814,a13816,a13818,a13820,a13822,a13824,a13826,a13828,a13830,a13832,
a13834,a13836,a13838,a13840,a13842,a13844,a13846,a13848,a13850,a13852,a13854,a13856,a13858,a13860,a13862,
a13864,a13866,a13868,a13870,a13872,a13874,a13876,a13878,a13880,a13882,a13884,a13886,a13888,a13890,a13892,
a13894,a13896,a13898,a13900,a13902,a13904,a13906,a13908,a13910,a13912,a13914,a13916,a13918,a13920,a13922,
a13924,a13926,a13928,a13930,a13932,a13934,a13936,a13938,a13940,a13942,a13944,a13946,a13948,a13950,a13952,
a13954,a13956,a13958,a13960,a13962,a13964,a13966,a13968,a13970,a13972,a13974,a13976,a13978,a13980,a13982,
a13984,a13986,a13988,a13990,a13992,a13994,a13996,a13998,a14000,a14002,a14004,a14006,a14008,a14010,a14012,
a14014,a14016,a14018,a14020,a14022,a14024,a14026,a14028,a14030,a14032,a14034,a14036,a14038,a14040,a14042,
a14044,a14046,a14048,a14050,a14052,a14054,a14056,a14058,a14060,a14062,a14064,a14066,a14068,a14070,a14072,
a14074,a14076,a14078,a14080,a14082,a14084,a14086,a14088,a14090,a14092,a14094,a14096,a14098,a14100,a14102,
a14104,a14106,a14108,a14110,a14112,a14114,a14116,a14118,a14120,a14122,a14124,a14126,a14128,a14130,a14132,
a14134,a14136,a14138,a14140,a14142,a14144,a14146,a14148,a14150,a14152,a14154,a14156,a14158,a14160,a14162,
a14164,a14166,a14168,a14170,a14172,a14174,a14176,a14178,a14180,a14182,a14184,a14186,a14188,a14190,a14192,
a14194,a14196,a14198,a14200,a14202,a14204,a14206,a14208,a14210,a14212,a14214,a14216,a14218,a14220,a14222,
a14224,a14226,a14228,a14230,a14232,a14234,a14236,a14238,a14240,a14242,a14244,a14246,a14248,a14250,a14252,
a14254,a14256,a14258,a14260,a14262,a14264,a14266,a14268,a14270,a14272,a14274,a14276,a14278,a14280,a14282,
a14284,a14286,a14288,a14290,a14292,a14294,a14296,a14298,a14300,a14302,a14304,a14306,a14308,a14310,a14312,
a14314,a14316,a14318,a14320,a14322,a14324,a14326,a14328,a14330,a14332,a14334,a14336,a14338,a14340,a14342,
a14344,a14346,a14348,a14350,a14352,a14354,a14356,a14358,a14360,a14362,a14364,a14366,a14368,a14370,a14372,
a14374,a14376,a14378,a14380,a14382,a14384,a14386,a14388,a14390,a14392,a14394,a14396,a14398,a14400,a14402,
a14404,a14406,a14408,a14410,a14412,a14414,a14416,a14418,a14420,a14422,a14424,a14426,a14428,a14430,a14432,
a14434,a14436,a14438,a14440,a14442,a14444,a14446,a14448,a14450,a14452,a14454,a14456,a14458,a14460,a14462,
a14464,a14466,a14468,a14470,a14472,a14474,a14476,a14478,a14480,a14482,a14484,a14486,a14488,a14490,a14492,
a14494,a14496,a14498,a14500,a14502,a14504,a14506,a14508,a14510,a14512,a14514,a14516,a14518,a14520,a14522,
a14524,a14526,a14528,a14530,a14532,a14534,a14536,a14538,a14540,a14542,a14544,a14546,a14548,a14550,a14552,
a14554,a14556,a14558,a14560,a14562,a14564,a14566,a14568,a14570,a14572,a14574,a14576,a14578,a14580,a14582,
a14584,a14586,a14588,a14590,a14592,a14594,a14596,a14598,a14600,a14602,a14604,a14606,a14608,a14610,a14612,
a14614,a14616,a14618,a14620,a14622,a14624,a14626,a14628,a14630,a14632,a14634,a14636,a14638,a14640,a14642,
a14644,a14646,a14648,a14650,a14652,a14654,a14656,a14658,a14660,a14662,a14664,a14666,a14668,a14670,a14672,
a14674,a14676,a14678,a14680,a14682,a14684,a14686,a14688,a14690,a14692,a14694,a14696,a14698,a14700,a14702,
a14704,a14706,a14708,a14710,a14712,a14714,a14716,a14718,a14720,a14722,a14724,a14726,a14728,a14730,a14732,
a14734,a14736,a14738,a14740,a14742,a14744,a14746,a14748,a14750,a14752,a14754,a14756,a14758,a14760,a14762,
a14764,a14766,a14768,a14770,a14772,a14774,a14776,a14778,a14780,a14782,a14784,a14786,a14788,a14790,a14792,
a14794,a14796,a14798,a14800,a14802,a14804,a14806,a14808,a14810,a14812,a14814,a14816,a14818,a14820,a14822,
a14824,a14826,a14828,a14830,a14832,a14834,a14836,a14838,a14840,a14842,a14844,a14846,a14848,a14850,a14852,
a14854,a14856,a14858,a14860,a14862,a14864,a14866,a14868,a14870,a14872,a14874,a14876,a14878,a14880,a14882,
a14884,a14886,a14888,a14890,a14892,a14894,a14896,a14898,a14900,a14902,a14904,a14906,a14908,a14910,a14912,
a14914,a14916,a14918,a14920,a14922,a14924,a14926,a14928,a14930,a14932,a14934,a14936,a14938,a14940,a14942,
a14944,a14946,a14948,a14950,a14952,a14954,a14956,a14958,a14960,a14962,a14964,a14966,a14968,a14970,a14972,
a14974,a14976,a14978,a14980,a14982,a14984,a14986,a14988,a14990,a14992,a14994,a14996,a14998,a15000,a15002,
a15004,a15006,a15008,a15010,a15012,a15014,a15016,a15018,a15020,a15022,a15024,a15026,a15028,a15030,a15032,
a15034,a15036,a15038,a15040,a15042,a15044,a15046,a15048,a15050,a15052,a15054,a15056,a15058,a15060,a15062,
a15064,a15066,a15068,a15070,a15072,a15074,a15076,a15078,a15080,a15082,a15084,a15086,a15088,a15090,a15092,
a15094,a15096,a15098,a15100,a15102,a15104,a15106,a15108,a15110,a15112,a15114,a15116,a15118,a15120,a15122,
a15124,a15126,a15128,a15130,a15132,a15134,a15136,a15138,a15140,a15142,a15144,a15146,a15148,a15150,a15152,
a15154,a15156,a15158,a15160,a15162,a15164,a15166,a15168,a15170,a15172,a15174,a15176,a15178,a15180,a15182,
a15184,a15186,a15188,a15190,a15192,a15194,a15196,a15198,a15200,a15202,a15204,a15206,a15208,a15210,a15212,
a15214,a15216,a15218,a15220,a15222,a15224,a15226,a15228,a15230,a15232,a15234,a15236,a15238,a15240,a15242,
a15244,a15246,a15248,a15250,a15252,a15254,a15256,a15258,a15260,a15262,a15264,a15266,a15268,a15270,a15272,
a15274,a15276,a15278,a15280,a15282,a15284,a15286,a15288,a15290,a15292,a15294,a15298,a15300,a15302,a15304,
a15306,a15308,a15310,a15312,a15316,a15318,a15320,a15322,a15324,a15326,a15328,a15330,a15332,a15334,a15336,
a15338,a15340,a15342,a15344,a15346,a15348,a15350,a15352,a15354,a15356,a15358,a15360,a15362,a15364,a15366,
a15368,a15372,a15374,a15376,a15378,a15380,a15382,a15384,a15386,a15388,a15390,a15392,a15394,a15396,a15398,
a15400,a15402,a15404,a15406,a15408,a15410,a15412,a15414,a15416,a15418,a15420,a15422,a15424,a15426,a15428,
a15430,a15432,a15434,a15436,a15438,a15440,a15442,a15444,a15446,a15450,a15452,a15454,a15456,a15458,a15460,
a15462,a15464,a15466,a15468,a15470,a15472,a15476,a15478,a15480,a15482,a15484,a15486,a15488,a15490,a15492,
a15494,a15496,a15498,a15500,a15502,a15504,a15506,a15508,a15510,a15512,a15514,a15516,a15518,a15520,a15522,
a15524,a15526,a15528,a15530,a15532,a15534,a15536,a15538,a15540,a15542,a15544,a15546,a15548,a15550,a15554,
a15556,a15558,a15560,a15562,a15564,a15566,a15568,a15570,a15572,a15574,a15576,a15580,a15582,a15584,a15586,
a15588,a15590,a15592,a15594,a15596,a15598,a15600,a15602,a15604,a15606,a15608,a15610,a15612,a15614,a15616,
a15618,a15620,a15622,a15624,a15626,a15628,a15630,a15632,a15634,a15636,a15638,a15640,a15642,a15644,a15646,
a15648,a15650,a15652,a15654,a15658,a15660,a15662,a15664,a15666,a15668,a15670,a15672,a15674,a15676,a15678,
a15680,a15684,a15686,a15688,a15690,a15692,a15694,a15696,a15698,a15700,a15702,a15704,a15706,a15708,a15710,
a15712,a15714,a15716,a15718,a15720,a15722,a15724,a15726,a15728,a15730,a15732,a15734,a15736,a15738,a15740,
a15742,a15744,a15746,a15748,a15750,a15752,a15754,a15756,a15758,a15762,a15764,a15766,a15768,a15770,a15772,
a15774,a15776,a15778,a15780,a15782,a15784,a15788,a15790,a15792,a15794,a15796,a15798,a15800,a15802,a15804,
a15806,a15808,a15810,a15812,a15814,a15816,a15818,a15820,a15822,a15824,a15826,a15828,a15830,a15832,a15834,
a15836,a15838,a15840,a15842,a15844,a15846,a15848,a15850,a15852,a15854,a15856,a15860,a15862,a15864,a15866,
a15868,a15870,a15872,a15874,a15876,a15878,a15880,a15882,a15886,a15888,a15890,a15892,a15894,a15896,a15898,
a15900,a15902,a15904,a15906,a15908,a15910,a15912,a15914,a15916,a15918,a15920,a15922,a15924,a15926,a15928,
a15930,a15932,a15934,a15936,a15938,a15940,a15942,a15944,a15946,a15948,a15950,a15952,a15954,a15958,a15960,
a15962,a15964,a15966,a15968,a15970,a15972,a15974,a15976,a15978,a15980,a15984,a15986,a15988,a15990,a15992,
a15994,a15996,a15998,a16000,a16002,a16004,a16006,a16008,a16010,a16012,a16014,a16016,a16018,a16020,a16022,
a16024,a16026,a16028,a16030,a16032,a16034,a16036,a16038,a16040,a16042,a16044,a16046,a16048,a16050,a16052,
a16054,a16056,a16058,a16060,a16062,a16064,a16066,a16068,a16072,a16074,a16076,a16078,a16080,a16082,a16084,
a16086,a16088,a16090,a16092,a16094,a16096,a16098,a16100,a16102,a16104,a16106,a16108,a16110,a16112,a16114,
a16116,a16118,a16120,a16122,a16124,a16126,a16128,a16130,a16132,a16134,a16136,a16138,a16140,a16142,a16144,
a16146,a16148,a16150,a16152,a16154,a16156,a16158,a16160,a16162,a16164,a16166,a16168,a16170,a16172,a16174,
a16176,a16178,a16180,a16182,a16184,a16186,a16188,a16190,a16192,a16194,a16196,a16198,a16200,a16202,a16204,
a16206,a16208,a16210,a16212,a16214,a16216,a16218,a16220,a16222,a16224,a16226,a16228,a16230,a16232,a16234,
a16236,a16238,a16240,a16242,a16244,a16246,a16248,a16250,a16252,a16254,a16256,a16258,a16260,a16262,a16264,
a16266,a16270,a16272,a16276,a16278,a16282,a16284,a16288,a16290,a16294,a16296,a16300,a16302,a16306,a16308,
a16312,a16314,a16316,a16318,a16320,a16322,a16324,a16326,a16328,a16330,a16332,a16334,a16336,a16338,a16340,
a16342,a16344,a16346,a16348,a16350,a16352,a16354,a16358,a16360,a16362,a16364,a16366,a16368,a16370,a16372,
a16374,a16376,a16378,a16380,a16382,a16384,a16386,a16388,a16390,a16392,a16394,a16396,a16398,a16400,a16402,
a16404,a16406,a16408,a16410,a16412,a16414,a16416,a16418,a16420,a16422,a16424,a16426,a16428,a16430,a16432,
a16434,a16436,a16438,a16440,a16442,a16444,a16446,a16448,a16450,a16452,a16454,a16456,a16458,a16460,a16462,
a16464,a16466,a16468,a16470,a16472,a16474,a16476,a16478,a16480,a16482,a16484,a16486,a16488,a16490,a16492,
a16494,a16496,a16498,a16500,a16502,a16504,a16506,a16508,a16510,a16512,a16514,a16516,a16518,a16520,a16522,
a16524,a16526,a16528,a16530,a16532,a16534,a16536,a16538,a16540,a16542,a16544,a16546,a16548,a16550,a16552,
a16554,a16556,a16558,a16560,a16562,a16564,a16566,a16568,a16570,a16572,a16574,a16576,a16578,a16580,a16582,
a16584,a16586,a16588,a16590,a16592,a16594,a16596,a16598,a16600,a16602,a16604,a16606,a16608,a16610,a16612,
a16614,a16616,a16618,a16620,a16622,a16624,a16626,a16628,a16630,a16632,a16634,a16636,a16638,a16640,a16642,
a16644,a16646,a16648,a16650,a16652,a16654,a16656,a16658,a16662,a16664,a16666,a16668,a16670,a16672,a16676,
a16678,a16680,a16682,a16684,a16686,a16688,a16690,a16692,a16694,a16696,a16698,a16700,a16702,a16704,a16706,
a16708,a16710,a16712,a16714,a16716,a16718,a16720,a16722,a16724,a16726,a16728,a16730,a16732,a16734,a16736,
a16738,a16740,a16742,a16744,a16746,a16748,a16750,a16752,a16754,a16756,a16758,a16760,a16762,a16764,a16766,
a16768,a16770,a16772,a16774,a16776,a16778,a16780,a16782,a16784,a16786,a16788,a16790,a16792,a16794,a16796,
a16798,a16802,a16804,a16806,a16810,a16812,a16814,a16816,a16818,a16820,a16822,a16824,a16826,a16828,a16830,
a16832,a16834,a16836,a16838,a16840,a16842,a16844,a16846,a16848,a16850,a16852,a16854,a16856,a16858,a16860,
a16862,a16864,a16866,a16868,a16870,a16872,a16874,a16876,a16878,a16880,a16882,a16884,a16886,a16888,a16890,
a16892,a16894,a16896,a16898,a16900,a16902,a16904,a16906,a16908,a16910,a16912,a16914,a16916,a16918,a16920,
a16922,a16924,a16926,a16928,a16930,a16932,a16934,a16938,a16940,a16942,a16944,a16946,a16948,a16952,a16954,
a16956,a16958,a16960,a16962,a16964,a16966,a16968,a16970,a16972,a16974,a16976,a16978,a16980,a16982,a16984,
a16986,a16988,a16990,a16992,a16994,a16996,a16998,a17000,a17002,a17004,a17006,a17008,a17010,a17012,a17014,
a17016,a17018,a17020,a17022,a17024,a17026,a17028,a17030,a17032,a17034,a17036,a17038,a17040,a17042,a17044,
a17046,a17048,a17050,a17052,a17054,a17056,a17058,a17060,a17062,a17064,a17066,a17068,a17070,a17074,a17076,
a17078,a17080,a17084,a17086,a17088,a17090,a17092,a17094,a17096,a17098,a17100,a17102,a17104,a17106,a17108,
a17110,a17112,a17114,a17116,a17118,a17120,a17122,a17124,a17126,a17128,a17130,a17132,a17134,a17136,a17138,
a17140,a17142,a17144,a17146,a17148,a17150,a17152,a17154,a17156,a17158,a17160,a17162,a17164,a17166,a17168,
a17170,a17172,a17174,a17176,a17178,a17180,a17182,a17184,a17186,a17188,a17190,a17192,a17194,a17196,a17198,
a17200,a17202,a17204,a17206,a17210,a17212,a17214,a17218,a17220,a17222,a17224,a17226,a17228,a17230,a17232,
a17234,a17236,a17238,a17240,a17242,a17244,a17246,a17248,a17250,a17252,a17254,a17256,a17258,a17260,a17262,
a17264,a17266,a17268,a17270,a17272,a17274,a17276,a17278,a17280,a17282,a17284,a17286,a17288,a17290,a17292,
a17294,a17296,a17298,a17300,a17302,a17304,a17306,a17308,a17310,a17312,a17314,a17316,a17318,a17320,a17322,
a17324,a17326,a17328,a17330,a17332,a17334,a17336,a17338,a17340,a17344,a17346,a17348,a17352,a17354,a17356,
a17358,a17360,a17362,a17364,a17366,a17368,a17370,a17372,a17374,a17376,a17378,a17380,a17382,a17384,a17386,
a17388,a17390,a17392,a17394,a17396,a17398,a17400,a17402,a17404,a17406,a17408,a17410,a17412,a17414,a17416,
a17418,a17420,a17422,a17424,a17426,a17428,a17430,a17432,a17434,a17436,a17438,a17440,a17442,a17444,a17446,
a17448,a17450,a17452,a17454,a17456,a17458,a17460,a17462,a17464,a17466,a17468,a17470,a17472,a17474,a17478,
a17480,a17482,a17484,a17486,a17490,a17492,a17494,a17496,a17498,a17500,a17502,a17504,a17506,a17508,a17510,
a17512,a17514,a17516,a17518,a17520,a17522,a17524,a17526,a17528,a17530,a17532,a17534,a17536,a17538,a17540,
a17542,a17544,a17546,a17548,a17550,a17552,a17554,a17556,a17558,a17560,a17562,a17564,a17566,a17568,a17570,
a17572,a17574,a17576,a17578,a17580,a17582,a17584,a17586,a17588,a17590,a17592,a17594,a17596,a17598,a17600,
a17602,a17604,a17606,a17608,a17612,a17614,a17618,a17620,a17622,a17624,a17626,a17628,a17630,a17632,a17634,
a17636,a17638,a17640,a17642,a17644,a17646,a17648,a17650,a17652,a17654,a17656,a17658,a17660,a17662,a17664,
a17666,a17668,a17670,a17672,a17674,a17676,a17678,a17680,a17682,a17684,a17686,a17688,a17690,a17692,a17694,
a17696,a17698,a17700,a17702,a17704,a17706,a17708,a17710,a17712,a17714,a17716,a17718,a17720,a17722,a17724,
a17726,a17728,a17730,a17732,a17734,a17736,a17738,a17740,a17744,a17746,a17750,a17752,a17754,a17756,a17758,
a17760,a17762,a17764,a17766,a17768,a17770,a17772,a17774,a17776,a17778,a17780,a17782,a17784,a17786,a17788,
a17790,a17792,a17794,a17796,a17798,a17800,a17802,a17804,a17806,a17808,a17810,a17812,a17814,a17816,a17818,
a17820,a17822,a17824,a17826,a17828,a17830,a17832,a17834,a17836,a17838,a17840,a17842,a17844,a17846,a17848,
a17850,a17852,a17854,a17856,a17858,a17860,a17862,a17864,a17866,a17868,a17870,a17874,a17876,a17878,a17880,
a17884,a17886,a17888,a17890,a17892,a17894,a17896,a17898,a17902,a17904,a17906,a17908,a17910,a17912,a17914,
a17918,a17920,a17922,a17924,a17926,a17928,a17930,a17932,a17934,a17936,a17938,a17940,a17942,a17944,a17946,
a17948,a17950,a17952,a17954,a17956,a17958,a17960,a17962,a17964,a17966,a17968,a17970,a17972,a17974,a17976,
a17978,a17980,a17982,a17984,a17986,a17988,a17990,a17992,a17994,a17996,a17998,a18000,a18002,a18004,a18006,
a18008,a18010,a18012,a18014,a18016,a18018,a18020,a18022,a18024,a18028,a18030,a18032,a18034,a18036,a18038,
a18040,a18042,a18044,a18046,a18048,a18050,a18052,a18054,a18056,a18058,a18060,a18062,a18064,a18066,a18068,
a18070,a18072,a18074,a18076,a18078,a18080,a18082,a18084,a18086,a18088,a18090,a18092,a18094,a18096,a18100,
a18102,a18104,a18106,a18108,a18110,a18112,a18114,a18116,a18118,a18120,a18122,a18124,a18126,a18128,a18130,
a18132,a18134,a18136,a18138,a18140,a18142,a18144,a18146,a18148,a18150,a18152,a18154,a18156,a18158,a18160,
a18162,a18164,a18166,a18168,a18170,a18172,a18174,a18176,a18178,a18180,a18182,a18184,a18186,a18188,a18190,
a18192,a18194,a18196,a18198,a18200,a18202,a18204,a18206,a18208,a18210,a18212,a18214,a18216,a18218,a18220,
a18222,a18224,a18226,a18228,a18230,a18232,a18234,a18236,a18238,a18240,a18242,a18244,a18246,a18248,a18250,
a18252,a18254,a18256,a18258,a18260,a18262,a18264,a18266,a18268,a18270,a18272,a18274,a18276,a18278,a18280,
a18282,a18284,a18286,a18288,a18290,a18292,a18294,a18296,a18298,a18300,a18302,a18304,a18306,a18308,a18310,
a18312,a18314,a18316,a18318,a18320,a18322,a18324,a18326,a18328,a18330,a18332,a18334,a18336,a18338,a18340,
a18342,a18344,a18346,a18348,a18350,a18352,a18354,a18356,a18358,a18360,a18362,a18364,a18366,a18368,a18370,
a18372,a18374,a18376,a18378,a18380,a18382,a18384,a18386,a18388,a18390,a18392,a18394,a18396,a18398,a18400,
a18402,a18404,a18406,a18408,a18410,a18412,a18414,a18416,a18418,a18420,a18422,a18424,a18426,a18428,a18430,
a18432,a18434,a18436,a18438,a18440,a18442,a18444,a18446,a18448,a18450,a18452,a18454,a18456,a18458,a18460,
a18462,a18464,a18466,a18468,a18470,a18472,a18474,a18476,a18478,a18480,a18482,a18484,a18486,a18488,a18490,
a18492,a18494,a18496,a18498,a18500,a18502,a18504,a18506,a18508,a18510,a18512,a18514,a18516,a18518,a18520,
a18522,a18524,a18526,a18528,a18530,a18532,a18534,a18536,a18538,a18540,a18542,a18544,a18546,a18548,a18550,
a18552,a18554,a18556,a18558,a18560,a18562,a18564,a18566,a18568,a18570,a18572,a18574,a18576,a18578,a18580,
a18582,a18584,a18586,a18588,a18590,a18592,a18594,a18596,a18598,a18600,a18602,a18604,a18606,a18608,a18610,
a18612,a18614,a18616,a18618,a18620,a18622,a18624,a18626,a18628,a18630,a18632,a18634,a18636,a18638,a18640,
a18642,a18644,a18646,a18648,a18650,a18652,a18654,a18656,a18658,a18660,a18662,a18664,a18666,a18668,a18670,
a18672,a18674,a18676,a18678,a18680,a18682,a18684,a18686,a18688,a18690,a18692,a18694,a18696,a18698,a18700,
a18702,a18704,a18706,a18708,a18710,a18712,a18714,a18716,a18718,a18720,a18722,a18724,a18726,a18728,a18730,
a18732,a18734,a18736,a18738,a18740,a18742,a18744,a18746,a18748,a18750,a18752,a18754,a18756,a18758,a18760,
a18762,a18764,a18766,a18768,a18770,a18772,a18774,a18776,a18778,a18780,a18782,a18784,a18786,a18788,a18790,
a18792,a18794,a18796,a18798,a18800,a18802,a18804,a18806,a18808,a18810,a18812,a18814,a18816,a18818,a18820,
a18822,a18824,a18826,a18828,a18830,a18832,a18834,a18836,a18838,a18840,a18842,a18844,a18846,a18848,a18850,
a18852,a18854,a18856,a18858,a18860,a18862,a18864,a18866,a18868,a18870,a18872,a18874,a18876,a18878,a18880,
a18882,a18884,a18886,a18888,a18890,a18892,a18894,a18896,a18898,a18900,a18902,a18904,a18906,a18908,a18910,
a18912,a18914,a18916,a18918,a18920,a18922,a18924,a18926,a18928,a18930,a18932,a18934,a18936,a18938,a18940,
a18942,a18944,a18946,a18948,a18950,a18952,a18954,a18956,a18958,a18960,a18962,a18964,a18966,a18968,a18970,
a18972,a18974,a18976,a18978,a18980,a18982,a18984,a18986,a18988,a18990,a18992,a18994,a18996,a18998,a19000,
a19002,a19004,a19006,a19008,a19010,a19012,a19014,a19016,a19018,a19020,a19022,a19024,a19026,a19028,a19030,
a19032,a19034,a19036,a19038,a19040,a19042,a19044,a19046,a19048,a19050,a19052,a19054,a19056,a19058,a19060,
a19062,a19064,a19066,a19068,a19070,a19072,a19074,a19076,a19078,a19080,a19082,a19084,a19086,a19088,a19090,
a19092,a19094,a19096,a19098,a19100,a19102,a19104,a19106,a19108,a19110,a19112,a19114,a19116,a19118,a19120,
a19122,a19124,a19126,a19128,a19130,a19132,a19134,a19136,a19138,a19140,a19142,a19144,a19146,a19148,a19150,
a19152,a19154,a19156,a19158,a19160,a19162,a19164,a19166,a19168,a19170,a19172,a19174,a19176,a19178,a19180,
a19182,a19184,a19186,a19188,a19190,a19192,a19194,a19196,a19198,a19200,a19202,a19204,a19206,a19210,a19212,
a19214,a19216,a19218,a19220,a19222,a19224,a19226,a19228,a19230,a19232,a19234,a19236,a19238,a19240,a19242,
a19244,a19246,a19250,a19252,a19254,a19256,a19258,a19260,a19264,a19266,a19268,a19270,a19272,a19276,a19278,
a19280,a19284,a19286,a19288,a19290,a19294,a19296,a19298,a19302,a19304,a19306,a19310,a19312,a19314,a19316,
a19320,a19322,a19324,a19328,a19330,a19332,a19338,a19340,a19344,a19346,a19350,a19352,a19356,a19358,a19362,
a19366,a19368,a19370,a19372,a19374,a19376,a19378,a19380,a19382,a19384,a19386,a19388,a19390,a19392,a19394,
a19396,a19398,a19400,a19402,a19404,a19406,a19408,a19410,a19412,a19414,a19416,a19418,a19420,a19422,a19424,
a19426,a19428,a19430,a19432,a19434,a19436,a19438,a19440,a19442,a19444,a19446,a19448,a19450,a19452,a19454,
a19456,a19458,a19460,a19462,a19464,a19466,a19468,a19470,a19472,a19476,a19478,a19480,a19482,a19486,a19488,
a19490,a19492,a19496,a19498,a19500,a19502,a19504,a19506,a19508,a19512,a19514,a19516,a19520,a19522,a19524,
a19528,a19530,a19532,a19536,a19538,a19540,a19542,a19544,a19546,a19548,a19550,a19552,a19554,a19556,a19558,
a19560,a19562,a19564,a19566,a19568,a19570,a19572,a19574,a19576,a19578,a19580,a19582,a19584,a19586,a19588,
a19590,a19592,a19594,a19596,a19598,a19600,a19602,a19604,a19606,a19608,a19610,a19612,a19614,a19616,a19618,
a19620,a19622,a19624,a19626,a19628,a19632,a19634,a19636,a19638,a19640,a19642,a19644,a19646,a19648,a19650,
a19652,a19654,a19656,a19658,a19660,a19662,a19666,a19668,a19670,a19672,a19674,a19676,a19678,a19680,a19682,
a19684,a19686,a19688,a19690,a19692,a19694,a19696,a19700,a19702,a19704,a19706,a19708,a19710,a19712,a19714,
a19716,a19718,a19720,a19722,a19724,a19726,a19728,a19730,a19734,a19736,a19738,a19740,a19742,a19744,a19746,
a19748,a19750,a19752,a19754,a19756,a19758,a19760,a19762,a19764,a19766,a19768,a19772,a19774,a19776,a19778,
a19780,a19782,a19784,a19786,a19788,a19790,a19792,a19794,a19796,a19798,a19800,a19802,a19804,a19806,a19810,
a19812,a19814,a19816,a19818,a19820,a19822,a19824,a19826,a19828,a19830,a19832,a19836,a19838,a19840,a19842,
a19844,a19846,a19848,a19850,a19852,a19854,a19856,a19858,a19860,a19862,a19864,a19866,a19868,a19870,a19872,
a19874,a19876,a19878,a19880,a19882,a19884,a19888,a19890,a19892,a19894,a19896,a19898,a19900,a19902,a19904,
a19906,a19908,a19910,a19914,a19916,a19918,a19920,a19922,a19928,a19930,a19932,a19934,a19936,a19940,a19942,
a19946,a19948,a19952,a19954,a19958,a19960,a19964,a19966,a19970,a19972,a19976,a19978,a19982,a19984,a19988,
a19990,a19994,a19996,a19998,a20000,a20002,a20006,a20008,a20012,a20014,a20018,a20020,a20024,a20026,a20030,
a20032,a20036,a20038,a20042,a20044,a20048,a20050,a20054,a20056,a20062,a20064,a20066,a20068,a20070,a20074,
a20076,a20080,a20082,a20086,a20088,a20092,a20094,a20098,a20100,a20104,a20106,a20110,a20112,a20116,a20118,
a20122,a20124,a20130,a20132,a20134,a20136,a20138,a20142,a20144,a20148,a20150,a20154,a20156,a20160,a20162,
a20166,a20168,a20172,a20174,a20178,a20180,a20184,a20186,a20190,a20192,a20198,a20200,a20202,a20204,a20206,
a20210,a20212,a20216,a20218,a20222,a20224,a20228,a20230,a20234,a20236,a20240,a20242,a20246,a20248,a20252,
a20254,a20258,a20260,a20266,a20268,a20270,a20272,a20274,a20278,a20280,a20284,a20286,a20290,a20292,a20296,
a20298,a20302,a20304,a20308,a20310,a20314,a20316,a20320,a20322,a20326,a20328,a20334,a20336,a20338,a20340,
a20342,a20346,a20348,a20352,a20354,a20358,a20360,a20364,a20366,a20370,a20372,a20376,a20378,a20382,a20384,
a20388,a20390,a20394,a20396,a20400,a20402,a20404,a20406,a20408,a20410,a20414,a20416,a20420,a20422,a20426,
a20428,a20432,a20434,a20438,a20440,a20444,a20446,a20450,a20452,a20456,a20458,a20462,a20464,a20468,a20470,
a20472,a20474,a20476,a20478,a20480,a20482,a20484,a20486,a20488,a20490,a20492,a20494,a20496,a20498,a20500,
a20502,a20504,a20506,a20508,a20510,a20512,a20514,a20516,a20518,a20520,a20522,a20524,a20526,a20528,a20530,
a20532,a20534,a20536,a20538,a20540,a20542,a20544,a20546,a20548,a20550,a20552,a20554,a20556,a20558,a20560,
a20562,a20566,a20568,a20570,a20572,a20574,a20576,a20578,a20580,a20582,a20584,a20586,a20588,a20590,a20592,
a20594,a20596,a20598,a20600,a20602,a20604,a20606,a20608,a20610,a20612,a20614,a20616,a20618,a20620,a20622,
a20624,a20626,a20628,a20630,a20632,a20634,a20638,a20640,a20642,a20644,a20646,a20648,a20650,a20652,a20654,
a20656,a20658,a20660,a20662,a20664,a20668,a20670,a20672,a20674,a20676,a20678,a20680,a20682,a20684,a20686,
a20688,a20690,a20692,a20694,a20696,a20698,a20700,a20702,a20704,a20706,a20708,a20710,a20712,a20714,a20718,
a20720,a20722,a20724,a20726,a20728,a20730,a20732,a20734,a20736,a20738,a20740,a20742,a20744,a20746,a20748,
a20750,a20752,a20754,a20756,a20758,a20760,a20764,a20766,a20768,a20770,a20772,a20774,a20776,a20778,a20780,
a20782,a20784,a20786,a20788,a20790,a20792,a20794,a20796,a20798,a20802,a20804,a20806,a20808,a20810,a20812,
a20814,a20818,a20820,a20822,a20824,a20826,a20828,a20830,a20832,a20834,a20838,a20840,a20842,a20844,a20846,
a20848,a20850,a20852,a20856,a20858,a20860,a20862,a20864,a20866,a20868,a20872,a20874,a20876,a20878,a20880,
a20882,a20884,a20886,a20888,a20890,a20892,a20894,a20896,a20900,a20902,a20904,a20906,a20908,a20910,a20912,
a20914,a20916,a20918,a20920,a20922,a20924,a20926,a20928,a20930,a20932,a20934,a20936,a20938,a20940,a20942,
a20944,a20946,a20948,a20950,a20952,a20954,a20956,a20958,a20960,a20962,a20964,a20966,a20968,a20970,a20972,
a20974,a20976,a20978,a20980,a20982,a20984,a20986,a20988,a20990,a20992,a20994,a20996,a20998,a21000,a21002,
a21004,a21006,a21008,a21010,a21012,a21014,a21016,a21018,a21020,a21022,a21024,a21026,a21028,a21030,a21032,
a21034,a21036,a21038,a21040,a21042,a21044,a21046,a21048,a21050,a21052,a21054,a21056,a21058,a21060,a21062,
a21064,a21066,a21068,a21070,a21072,a21074,a21076,a21078,a21080,a21082,a21084,a21086,a21088,a21090,a21092,
a21094,a21096,a21098,a21100,a21102,a21104,a21106,a21108,a21110,a21112,a21114,a21116,a21118,a21120,a21122,
a21124,a21126,a21128,a21130,a21132,a21134,a21136,a21138,a21140,a21142,a21144,a21146,a21148,a21150,a21152,
a21154,a21156,a21158,a21160,a21162,a21164,a21166,a21168,a21170,a21172,a21174,a21176,a21178,a21180,a21182,
a21184,a21186,a21188,a21190,a21192,a21194,a21196,a21198,a21200,a21202,a21204,a21206,a21208,a21210,a21212,
a21214,a21216,a21218,a21220,a21222,a21224,a21226,a21228,a21230,a21232,a21234,a21236,a21238,a21240,a21242,
a21244,a21246,a21248,a21250,a21252,a21254,a21256,a21258,a21260,a21262,a21264,a21266,a21268,a21270,a21272,
a21274,a21276,a21278,a21280,a21282,a21284,a21286,a21288,a21290,a21292,a21294,a21296,a21298,a21300,a21302,
a21304,a21306,a21308,a21310,a21312,a21314,a21316,a21318,a21320,a21322,a21324,a21326,a21328,a21330,a21332,
a21334,a21336,a21338,a21340,a21342,a21344,a21346,a21348,a21350,a21352,a21354,a21356,a21358,a21360,a21362,
a21364,a21366,a21368,a21370,a21372,a21374,a21376,a21378,a21380,a21382,a21384,a21386,a21388,a21390,a21392,
a21394,a21396,a21398,a21400,a21402,a21404,a21406,a21408,a21410,a21412,a21414,a21416,a21418,a21420,a21422,
a21424,a21426,a21428,a21430,a21432,a21434,a21436,a21438,a21440,a21442,a21444,a21446,a21448,a21450,a21452,
a21454,a21456,a21458,a21460,a21462,a21464,a21466,a21468,a21470,a21472,a21474,a21476,a21478,a21480,a21482,
a21484,a21486,a21488,a21490,a21492,a21494,a21496,a21498,a21500,a21502,a21504,a21506,a21508,a21510,a21512,
a21514,a21516,a21518,a21520,a21522,a21524,a21526,a21528,a21530,a21532,a21534,a21536,a21538,a21540,a21542,
a21544,a21546,a21548,a21550,a21552,a21554,a21556,a21558,a21560,a21562,a21564,a21566,a21568,a21570,a21572,
a21574,a21576,a21578,a21580,a21582,a21584,a21586,a21588,a21590,a21592,a21594,a21596,a21598,a21600,a21602,
a21604,a21606,a21608,a21610,a21612,a21614,a21616,a21618,a21620,a21622,a21624,a21626,a21628,a21630,a21632,
a21634,a21636,a21638,a21640,a21642,a21644,a21646,a21648,a21650,a21652,a21654,a21656,a21658,a21660,a21662,
a21664,a21666,a21668,a21670,a21672,a21674,a21676,a21678,a21680,a21682,a21684,a21686,a21688,a21690,a21692,
a21694,a21696,a21700,a21702,a21704,a21706,a21708,a21710,a21712,a21714,a21716,a21718,a21720,a21722,a21724,
a21726,a21728,a21730,a21732,a21734,a21736,a21738,a21740,a21742,a21744,a21746,a21748,a21750,a21752,a21754,
a21756,a21758,a21760,a21762,a21764,a21766,a21768,a21770,a21772,a21774,a21776,a21778,a21780,a21782,a21784,
a21786,a21788,a21790,a21792,a21794,a21796,a21798,a21800,a21802,a21804,a21806,a21808,a21810,a21812,a21814,
a21816,a21818,a21820,a21822,a21824,a21826,a21828,a21830,a21832,a21834,a21836,a21838,a21840,a21842,a21844,
a21846,a21848,a21850,a21852,a21854,a21856,a21858,a21860,a21862,a21864,a21866,a21868,a21870,a21872,a21874,
a21876,a21878,a21880,a21882,a21884,a21886,a21888,a21890,a21892,a21894,a21896,a21898,a21900,a21902,a21904,
a21906,a21908,a21910,a21912,a21914,a21916,a21918,a21920,a21922,a21924,a21926,a21928,a21930,a21932,a21934,
a21936,a21938,a21940,a21942,a21944,a21946,a21948,a21950,a21952,a21954,a21956,a21958,a21960,a21962,a21964,
a21966,a21968,a21970,a21972,a21974,a21976,a21978,a21980,a21982,a21984,a21986,a21988,a21990,a21992,a21994,
a21996,a21998,a22000,a22002,a22004,a22006,a22008,a22010,a22012,a22014,a22016,a22018,a22020,a22022,a22024,
a22026,a22028,a22030,a22032,a22034,a22036,a22038,a22040,a22042,a22044,a22046,a22048,a22050,a22052,a22054,
a22056,a22058,a22060,a22062,a22064,a22066,a22068,a22070,a22072,a22074,a22076,a22078,a22080,a22082,a22084,
a22086,a22088,a22090,a22092,a22094,a22096,a22098,a22100,a22102,a22104,a22106,a22108,a22110,a22112,a22114,
a22116,a22118,a22120,a22122,a22124,a22126,a22128,a22130,a22132,a22134,a22136,a22138,a22140,a22142,a22144,
a22146,a22148,a22150,a22152,a22154,a22156,a22158,a22160,a22162,a22164,a22166,a22168,a22170,a22174,a22176,
a22178,a22180,a22182,a22184,a22186,a22188,a22190,a22192,a22194,a22196,a22198,a22200,a22202,a22204,a22206,
a22208,a22210,a22212,a22214,a22216,a22218,a22220,a22222,a22224,a22226,a22228,a22232,a22234,a22236,a22238,
a22240,a22242,a22244,a22246,a22248,a22250,a22252,a22254,a22256,a22258,a22260,a22262,a22264,a22266,a22268,
a22270,a22272,a22274,a22276,a22278,a22280,a22282,a22284,a22286,a22290,a22292,a22294,a22296,a22298,a22300,
a22302,a22304,a22306,a22308,a22310,a22312,a22314,a22316,a22318,a22320,a22322,a22324,a22326,a22328,a22330,
a22332,a22334,a22336,a22338,a22340,a22342,a22344,a22348,a22350,a22352,a22354,a22356,a22358,a22360,a22362,
a22364,a22366,a22368,a22370,a22372,a22374,a22376,a22378,a22380,a22382,a22384,a22386,a22388,a22390,a22392,
a22394,a22396,a22398,a22400,a22402,a22406,a22408,a22410,a22412,a22414,a22416,a22418,a22420,a22422,a22424,
a22426,a22428,a22430,a22432,a22434,a22436,a22438,a22440,a22442,a22444,a22446,a22448,a22450,a22452,a22454,
a22456,a22458,a22460,a22464,a22466,a22468,a22470,a22472,a22474,a22476,a22478,a22480,a22482,a22484,a22486,
a22488,a22490,a22492,a22494,a22496,a22498,a22500,a22502,a22504,a22506,a22508,a22510,a22512,a22514,a22516,
a22518,a22522,a22524,a22526,a22528,a22530,a22532,a22534,a22536,a22538,a22540,a22542,a22544,a22546,a22548,
a22550,a22552,a22554,a22556,a22558,a22560,a22562,a22564,a22566,a22568,a22570,a22572,a22574,a22576,a22578,
a22580,a22582,a22584,a22586,a22588,a22590,a22592,a22594,a22596,a22598,a22602,a22604,a22606,a22608,a22610,
a22612,a22614,a22616,a22618,a22620,a22622,a22624,a22626,a22628,a22632,a22634,a22636,a22640,a22642,a22644,
a22646,a22648,a22650,a22652,a22654,a22658,a22660,a22662,a22666,a22672,a22674,a22678,a22680,a22682,a22684,
a22690,a22692,a22694,a22698,a22700,a22702,a22704,a22708,a22710,a22714,a22716,a22718,a22720,a22722,a22724,
a22726,a22728,a22730,a22732,a22734,a22736,a22738,a22740,a22742,a22744,a22746,a22748,a22752,a22754,a22756,
a22758,a22760,a22762,a22764,a22766,a22768,a22770,a22772,a22774,a22776,a22780,a22782,a22784,a22786,a22788,
a22790,a22792,a22794,a22796,a22798,a22800,a22802,a22804,a22808,a22810,a22812,a22814,a22816,a22818,a22820,
a22822,a22824,a22826,a22828,a22830,a22832,a22836,a22838,a22840,a22842,a22844,a22846,a22848,a22850,a22852,
a22854,a22856,a22858,a22860,a22864,a22866,a22868,a22870,a22872,a22874,a22876,a22878,a22880,a22882,a22884,
a22886,a22888,a22892,a22894,a22896,a22898,a22900,a22902,a22904,a22906,a22908,a22910,a22912,a22914,a22916,
a22920,a22922,a22924,a22926,a22928,a22930,a22932,a22934,a22936,a22938,a22940,a22942,a22944,a22948,a22950,
a22952,a22954,a22956,a22958,a22960,a22962,a22964,a22966,a22968,a22970,a22972,a22974,a22976,a22978,a22980,
a22982,a22984,a22986,a22988,a22990,a22992,a22994,a22996,a22998,a23000,a23002,a23004,a23006,a23008,a23010,
a23012,a23014,a23016,a23018,a23020,a23022,a23024,a23026,a23028,a23030,a23032,a23034,a23036,a23038,a23040,
a23042,a23044,a23046,a23048,a23050,a23052,a23054,a23056,a23058,a23060,a23062,a23064,a23066,a23068,a23070,
a23072,a23074,a23076,a23078,a23080,a23082,a23084,a23086,a23088,a23090,a23092,a23094,a23096,a23098,a23100,
a23102,a23104,a23106,a23108,a23110,a23112,a23114,a23116,a23118,a23120,a23122,a23124,a23126,a23128,a23130,
a23132,a23134,a23136,a23138,a23140,a23142,a23144,a23146,a23148,a23150,a23152,a23154,a23156,a23158,a23160,
a23162,a23164,a23166,a23168,a23170,a23172,a23174,a23176,a23178,a23180,a23182,a23184,a23186,a23188,a23190,
a23192,a23194,a23196,a23198,a23200,a23202,a23204,a23206,a23208,a23210,a23212,a23214,a23216,a23218,a23220,
a23222,a23224,a23226,a23228,a23230,a23232,a23234,a23236,a23238,a23240,a23242,a23244,a23246,a23248,a23250,
a23252,a23254,a23256,a23258,a23260,a23262,a23264,a23266,a23268,a23270,a23272,a23274,a23276,a23278,a23280,
a23282,a23284,a23286,a23288,a23290,a23292,a23294,a23296,a23298,a23300,a23302,a23304,a23306,a23308,a23310,
a23312,a23314,a23316,a23318,a23320,a23322,a23324,a23326,a23328,a23330,a23332,a23334,a23336,a23338,a23340,
a23342,a23344,a23346,a23348,a23350,a23352,a23354,a23356,a23358,a23360,a23362,a23364,a23366,a23368,a23370,
a23372,a23374,a23376,a23378,a23380,a23382,a23384,a23386,a23388,a23390,a23392,a23394,a23396,a23398,a23400,
a23402,a23404,a23406,a23408,a23410,a23412,a23414,a23416,a23418,a23420,a23422,a23424,a23426,a23428,a23430,
a23432,a23434,a23436,a23438,a23440,a23442,a23444,a23446,a23448,a23450,a23452,a23454,a23456,a23458,a23460,
a23462,a23464,a23466,a23468,a23470,a23472,a23474,a23476,a23478,a23480,a23482,a23484,a23486,a23488,a23490,
a23492,a23494,a23496,a23498,a23500,a23502,a23504,a23506,a23508,a23510,a23512,a23514,a23516,a23518,a23520,
a23522,a23524,a23526,a23528,a23530,a23532,a23534,a23536,a23538,a23540,a23542,a23544,a23546,a23548,a23550,
a23552,a23554,a23556,a23558,a23560,a23562,a23564,a23566,a23568,a23570,a23572,a23574,a23576,a23578,a23580,
a23582,a23584,a23586,a23588,a23590,a23592,a23594,a23596,a23598,a23600,a23602,a23604,a23606,a23608,a23610,
a23612,a23614,a23616,a23618,a23620,a23622,a23624,a23626,a23628,a23630,a23632,a23634,a23636,a23638,a23640,
a23642,a23644,a23646,a23648,a23650,a23652,a23654,a23656,a23658,a23660,a23662,a23664,a23666,a23668,a23670,
a23672,a23674,a23676,a23678,a23680,a23682,a23684,a23686,a23688,a23690,a23692,a23694,a23696,a23698,a23700,
a23702,a23704,a23706,a23708,a23710,a23712,a23714,a23716,a23718,a23720,a23722,a23724,a23726,a23728,a23730,
a23732,a23734,a23736,a23738,a23740,a23742,a23744,a23746,a23748,a23750,a23752,a23754,a23756,a23758,a23760,
a23762,a23764,a23766,a23768,a23770,a23772,a23774,a23776,a23778,a23780,a23782,a23784,a23786,a23788,a23790,
a23792,a23794,a23796,a23798,a23800,a23802,a23804,a23806,a23808,a23810,a23812,a23814,a23816,a23818,a23820,
a23822,a23824,a23826,a23828,a23830,a23832,a23834,a23836,a23838,a23840,a23842,a23844,a23846,a23848,a23850,
a23852,a23854,a23856,a23858,a23860,a23862,a23864,a23866,a23868,a23870,a23872,a23874,a23876,a23878,a23880,
a23882,a23884,a23886,a23888,a23890,a23892,a23894,a23896,a23898,a23900,a23902,a23904,a23906,a23908,a23910,
a23912,a23914,a23916,a23918,a23920,a23922,a23924,a23926,a23928,a23930,a23932,a23934,a23936,a23938,a23940,
a23942,a23944,a23946,a23948,a23950,a23952,a23954,a23956,a23958,a23960,a23962,a23964,a23966,a23968,a23970,
a23972,a23974,a23976,a23978,a23980,a23982,a23984,a23986,a23988,a23990,a23992,a23994,a23996,a23998,a24000,
a24002,a24004,a24006,a24008,a24010,a24012,a24014,a24016,a24018,a24020,a24022,a24024,a24026,a24028,a24030,
a24032,a24034,a24036,a24038,a24040,a24042,a24044,a24046,a24048,a24050,a24052,a24054,a24056,a24058,a24060,
a24062,a24064,a24066,a24068,a24070,a24072,a24074,a24076,a24078,a24080,a24082,a24084,a24086,a24088,a24090,
a24092,a24094,a24096,a24098,a24100,a24102,a24104,a24106,a24108,a24110,a24112,a24114,a24116,a24118,a24120,
a24122,a24124,a24126,a24128,a24130,a24132,a24134,a24136,a24138,a24140,a24142,a24144,a24146,a24148,a24150,
a24152,a24154,a24156,a24158,a24160,a24162,a24164,a24166,a24168,a24170,a24172,a24174,a24176,a24178,a24180,
a24182,a24184,a24186,a24188,a24190,a24192,a24194,a24196,a24198,a24200,a24202,a24204,a24206,a24208,a24210,
a24212,a24214,a24216,a24218,a24220,a24222,a24224,a24226,a24228,a24230,a24232,a24234,a24236,a24238,a24240,
a24242,a24244,a24246,a24248,a24250,a24252,a24254,a24256,a24258,a24260,a24262,a24264,a24266,a24268,a24270,
a24272,a24274,a24276,a24278,a24280,a24282,a24284,a24286,a24288,a24290,a24292,a24294,a24296,a24298,a24300,
a24302,a24304,a24306,a24308,a24310,a24312,a24314,a24316,a24318,a24320,a24322,a24324,a24326,a24328,a24330,
a24332,a24334,a24336,a24338,a24340,a24342,a24344,a24346,a24348,a24350,a24352,a24354,a24356,a24358,a24360,
a24362,a24364,a24366,a24368,a24370,a24372,a24374,a24376,a24378,a24380,a24382,a24384,a24386,a24388,a24390,
a24392,a24394,a24396,a24398,a24400,a24402,a24404,a24406,a24408,a24410,a24412,a24414,a24416,a24418,a24420,
a24422,a24424,a24426,a24428,a24430,a24432,a24434,a24436,a24438,a24440,a24444,a24446,a24448,a24450,a24452,
a24454,a24456,a24458,a24460,a24462,a24464,a24466,a24468,a24470,a24472,a24474,a24476,a24478,a24480,a24482,
a24484,a24486,a24488,a24490,a24492,a24494,a24496,a24498,a24500,a24502,a24504,a24506,a24508,a24510,a24512,
a24514,a24516,a24518,a24520,a24522,a24524,a24526,a24528,a24530,a24532,a24534,a24536,a24538,a24540,a24542,
a24544,a24546,a24548,a24550,a24552,a24554,a24556,a24558,a24560,a24562,a24564,a24566,a24568,a24570,a24572,
a24574,a24576,a24578,a24580,a24582,a24584,a24586,a24588,a24590,a24592,a24594,a24596,a24598,a24600,a24602,
a24604,a24606,a24608,a24610,a24612,a24614,a24616,a24618,a24620,a24622,a24624,a24626,a24628,a24630,a24632,
a24634,a24636,a24638,a24640,a24642,a24644,a24646,a24648,a24650,a24652,a24654,a24656,a24658,a24662,a24664,
a24666,a24668,a24670,a24672,a24674,a24676,a24678,a24680,a24682,a24684,a24686,a24688,a24690,a24692,a24694,
a24696,a24698,a24700,a24702,a24704,a24706,a24708,a24710,a24712,a24714,a24716,a24718,a24722,a24724,a24726,
a24730,a24732,a24734,a24736,a24738,a24742,a24744,a24746,a24750,a24752,a24754,a24756,a24758,a24760,a24762,
a24766,a24768,a24770,a24774,a24776,a24778,a24780,a24782,a24786,a24788,a24790,a24794,a24796,a24798,a24800,
a24802,a24804,a24806,a24808,a24810,a24814,a24816,a24818,a24822,a24824,a24826,a24828,a24830,a24832,a24834,
a24836,a24838,a24840,a24842,a24844,a24848,a24850,a24852,a24856,a24858,a24860,a24862,a24864,a24868,a24870,
a24872,a24876,a24878,a24880,a24882,a24884,a24886,a24888,a24892,a24894,a24896,a24900,a24902,a24904,a24906,
a24908,a24912,a24914,a24916,a24920,a24922,a24924,a24926,a24928,a24930,a24932,a24934,a24936,a24940,a24942,
a24944,a24948,a24950,a24952,a24954,a24956,a24958,a24960,a24962,a24964,a24966,a24968,a24972,a24974,a24976,
a24980,a24982,a24984,a24986,a24988,a24992,a24994,a24996,a25000,a25002,a25004,a25006,a25008,a25010,a25012,
a25016,a25018,a25020,a25024,a25026,a25028,a25030,a25032,a25036,a25038,a25040,a25044,a25046,a25048,a25050,
a25052,a25054,a25056,a25058,a25060,a25064,a25066,a25068,a25072,a25074,a25076,a25078,a25080,a25082,a25084,
a25086,a25088,a25090,a25092,a25096,a25098,a25100,a25104,a25106,a25108,a25110,a25112,a25116,a25118,a25120,
a25124,a25126,a25128,a25130,a25132,a25134,a25136,a25140,a25142,a25144,a25148,a25150,a25152,a25154,a25156,
a25160,a25162,a25164,a25168,a25170,a25172,a25174,a25176,a25178,a25180,a25182,a25184,a25188,a25190,a25192,
a25196,a25198,a25200,a25202,a25204,a25206,a25208,a25210,a25212,a25214,a25216,a25220,a25222,a25224,a25228,
a25230,a25232,a25234,a25236,a25240,a25242,a25244,a25248,a25250,a25252,a25254,a25256,a25258,a25260,a25264,
a25266,a25268,a25272,a25274,a25276,a25278,a25280,a25284,a25286,a25288,a25292,a25294,a25296,a25298,a25300,
a25302,a25304,a25306,a25308,a25312,a25314,a25316,a25320,a25322,a25324,a25326,a25328,a25330,a25332,a25334,
a25336,a25338,a25340,a25344,a25346,a25348,a25352,a25354,a25356,a25358,a25360,a25364,a25366,a25368,a25372,
a25374,a25376,a25378,a25380,a25382,a25384,a25388,a25390,a25392,a25396,a25398,a25400,a25402,a25404,a25408,
a25410,a25412,a25416,a25418,a25420,a25422,a25424,a25426,a25428,a25430,a25432,a25436,a25438,a25440,a25444,
a25446,a25448,a25450,a25452,a25454,a25456,a25458,a25460,a25462,a25464,a25468,a25470,a25472,a25476,a25478,
a25480,a25482,a25484,a25488,a25490,a25492,a25496,a25498,a25500,a25502,a25504,a25506,a25508,a25512,a25514,
a25516,a25520,a25522,a25524,a25526,a25528,a25532,a25534,a25536,a25540,a25542,a25544,a25546,a25548,a25550,
a25552,a25554,a25556,a25560,a25562,a25564,a25568,a25570,a25572,a25574,a25576,a25578,a25580,a25582,a25584,
a25586,a25588,a25592,a25594,a25596,a25600,a25602,a25604,a25606,a25608,a25612,a25614,a25616,a25620,a25622,
a25624,a25626,a25628,a25630,a25632,a25636,a25638,a25640,a25644,a25646,a25648,a25650,a25652,a25656,a25658,
a25660,a25664,a25666,a25668,a25670,a25672,a25674,a25676,a25678,a25680,a25684,a25686,a25688,a25692,a25694,
a25696,a25698,a25700,a25702,a25704,a25706,a25708,a25710,a25712,a25714,a25716,a25718,a25720,a25722,a25724,
a25726,a25728,a25730,a25732,a25734,a25736,a25738,a25740,a25742,a25744,a25746,a25748,a25750,a25752,a25754,
a25756,a25758,a25760,a25762,a25764,a25766,a25768,a25770,a25772,a25774,a25776,a25778,a25780,a25782,a25784,
a25786,a25788,a25790,a25792,a25794,a25796,a25798,a25800,a25802,a25804,a25806,a25808,a25810,a25812,a25814,
a25816,a25818,a25820,a25822,a25824,a25826,a25828,a25830,a25832,a25834,a25836,a25838,a25840,a25842,a25844,
a25846,a25848,a25850,a25852,a25854,a25856,a25858,a25860,a25862,a25864,a25866,a25868,a25870,a25872,a25874,
a25876,a25878,a25880,a25882,a25884,a25886,a25888,a25890,a25892,a25894,a25896,a25898,a25900,a25902,a25904,
a25906,a25908,a25910,a25912,a25914,a25916,a25918,a25920,a25922,a25924,a25926,a25928,a25930,a25932,a25934,
a25936,a25938,a25940,a25942,a25944,a25946,a25948,a25950,a25952,a25954,a25956,a25958,a25960,a25962,a25964,
a25966,a25968,a25970,a25972,a25974,a25976,a25978,a25980,a25982,a25984,a25986,a25988,a25990,a25992,a25994,
a25996,a25998,a26000,a26002,a26004,a26006,a26008,a26010,a26012,a26014,a26016,a26018,a26020,a26022,a26024,
a26026,a26028,a26030,a26032,a26034,a26036,a26038,a26040,a26042,a26044,a26046,a26048,a26050,a26052,a26054,
a26056,a26058,a26060,a26062,a26064,a26066,a26068,a26070,a26072,a26074,a26076,a26078,a26080,a26082,a26084,
a26086,a26088,a26090,a26092,a26094,a26096,a26098,a26100,a26102,a26104,a26106,a26108,a26110,a26112,a26114,
a26116,a26118,a26120,a26122,a26124,a26126,a26128,a26130,a26132,a26134,a26136,a26138,a26140,a26142,a26144,
a26146,a26148,a26150,a26152,a26154,a26156,a26158,a26160,a26162,a26164,a26166,a26168,a26170,a26172,a26174,
a26176,a26178,a26180,a26182,a26184,a26186,a26188,a26190,a26192,a26194,a26196,a26198,a26200,a26202,a26204,
a26206,a26208,a26210,a26212,a26214,a26216,a26218,a26220,a26222,a26224,a26226,a26228,a26230,a26232,a26234,
a26236,a26238,a26240,a26242,a26244,a26246,a26248,a26250,a26252,a26254,a26256,a26258,a26260,a26262,a26264,
a26266,a26268,a26270,a26272,a26274,a26276,a26278,a26280,a26282,a26284,a26286,a26288,a26290,a26292,a26294,
a26296,a26298,a26300,a26302,a26304,a26306,a26308,a26310,a26312,a26314,a26316,a26318,a26320,a26322,a26324,
a26326,a26328,a26330,a26332,a26334,a26336,a26338,a26340,a26342,a26344,a26346,a26348,a26350,a26352,a26354,
a26356,a26358,a26360,a26362,a26364,a26366,a26368,a26370,a26372,a26374,a26376,a26378,a26380,a26382,a26384,
a26386,a26388,a26390,a26392,a26394,a26396,a26398,a26400,a26402,a26404,a26406,a26408,a26410,a26412,a26414,
a26416,a26418,a26420,a26422,a26424,a26426,a26428,a26430,a26432,a26434,a26436,a26438,a26440,a26442,a26444,
a26446,a26448,a26450,a26452,a26454,a26456,a26458,a26460,a26462,a26464,a26466,a26468,a26470,a26472,a26474,
a26476,a26478,a26480,a26482,a26484,a26486,a26488,a26490,a26492,a26494,a26496,a26498,a26500,a26502,a26504,
a26506,a26508,a26510,a26512,a26514,a26516,a26518,a26520,a26522,a26524,a26526,a26528,a26530,a26532,a26534,
a26536,a26538,a26540,a26542,a26544,a26546,a26548,a26550,a26552,a26554,a26556,a26558,a26560,a26562,a26564,
a26566,a26568,a26570,a26572,a26574,a26576,a26578,a26580,a26582,a26584,a26586,a26588,a26590,a26592,a26594,
a26596,a26598,a26600,a26602,a26606,a26608,a26610,a26612,a26618,a26620,a26624,a26626,a26628,a26630,a26632,
a26634,a26638,a26640,a26642,a26644,a26646,a26648,a26650,a26652,a26654,a26656,a26658,a26660,a26662,a26664,
a26666,a26668,a26670,a26672,a26674,a26676,a26678,a26680,a26682,a26684,a26686,a26688,a26690,a26692,a26694,
a26696,a26698,a26700,a26702,a26704,a26706,a26708,a26710,a26712,a26714,a26716,a26718,a26720,a26722,a26724,
a26726,a26728,a26730,a26732,a26734,a26736,a26738,a26740,a26742,a26744,a26746,a26748,a26750,a26752,a26754,
a26756,a26758,a26760,a26762,a26764,a26766,a26768,a26770,a26772,a26774,a26776,a26778,a26780,a26782,a26784,
a26786,a26788,a26790,a26792,a26794,a26796,a26798,a26800,a26802,a26804,a26806,a26808,a26810,a26812,a26814,
a26816,a26818,a26820,a26822,a26824,a26826,a26828,a26830,a26832,a26834,a26836,a26838,a26840,a26842,a26844,
a26846,a26848,a26850,a26852,a26854,a26856,a26858,a26860,a26862,a26864,a26866,a26868,a26870,a26872,a26874,
a26876,a26878,a26880,a26882,a26884,a26886,a26888,a26890,a26892,a26894,a26896,a26898,a26900,a26902,a26904,
a26906,a26908,a26910,a26912,a26914,a26916,a26918,a26920,a26922,a26924,a26926,a26928,a26930,a26932,a26934,
a26936,a26938,a26940,a26942,a26944,a26946,a26948,a26950,a26952,a26954,a26956,a26958,a26960,a26962,a26964,
a26966,a26968,a26970,a26972,a26974,a26976,a26978,a26980,a26982,a26984,a26986,a26988,a26990,a26992,a26994,
a26996,a26998,a27000,a27002,a27004,a27006,a27008,a27010,a27012,a27014,a27016,a27018,a27020,a27022,a27024,
a27026,a27028,a27030,a27032,a27034,a27036,a27038,a27040,a27042,a27044,a27046,a27048,a27050,a27052,a27054,
a27056,a27058,a27062,a27064,a27066,a27068,a27070,a27072,a27074,a27076,a27078,a27080,a27082,a27084,a27086,
a27088,a27090,a27092,a27094,a27096,a27098,a27100,a27102,a27104,a27106,a27110,a27112,a27114,a27116,a27118,
a27120,a27122,a27124,a27126,a27128,a27130,a27132,a27134,a27136,a27138,a27140,a27142,a27144,a27146,a27148,
a27150,a27152,a27154,a27158,a27160,a27162,a27164,a27166,a27168,a27170,a27172,a27174,a27176,a27178,a27180,
a27182,a27184,a27186,a27188,a27190,a27192,a27194,a27196,a27198,a27200,a27202,a27206,a27208,a27210,a27212,
a27214,a27216,a27218,a27220,a27222,a27224,a27226,a27228,a27230,a27232,a27234,a27236,a27238,a27240,a27242,
a27244,a27246,a27248,a27250,a27254,a27256,a27258,a27260,a27262,a27264,a27266,a27268,a27270,a27272,a27274,
a27276,a27278,a27280,a27282,a27284,a27286,a27288,a27290,a27292,a27294,a27296,a27298,a27302,a27304,a27306,
a27308,a27310,a27312,a27314,a27316,a27318,a27320,a27322,a27324,a27326,a27328,a27330,a27332,a27334,a27336,
a27338,a27340,a27342,a27344,a27346,a27350,a27352,a27354,a27356,a27358,a27360,a27362,a27364,a27366,a27368,
a27370,a27372,a27374,a27376,a27378,a27380,a27384,a27386,a27388,a27390,a27392,a27394,a27396,a27400,a27402,
a27404,a27406,a27408,a27410,a27412,a27416,a27418,a27420,a27422,a27424,a27426,a27428,a27432,a27434,a27436,
a27438,a27440,a27442,a27444,a27446,a27448,a27450,a27456,a27458,a27462,a27464,a27468,a27470,a27474,a27476,
a27480,a27482,a27486,a27488,a27492,a27494,a27496,a27500,a27502,a27504,a27506,a27508,a27510,a27512,a27514,
a27516,a27518,a27520,a27522,a27524,a27526,a27528,a27530,a27532,a27534,a27536,a27538,a27540,a27542,a27544,
a27546,a27548,a27550,a27552,a27554,a27556,a27558,a27560,a27562,a27564,a27566,a27568,a27570,a27574,a27576,
a27578,a27580,a27582,a27584,a27586,a27590,a27592,a27594,a27596,a27598,a27600,a27602,a27604,a27606,a27608,
a27610,a27612,a27614,a27616,a27618,a27620,a27622,a27624,a27626,a27628,a27632,a27634,a27636,a27638,a27640,
a27642,a27644,a27646,a27648,a27650,a27652,a27654,a27656,a27658,a27660,a27662,a27666,a27668,a27670,a27672,
a27674,a27676,a27678,a27680,a27682,a27686,a27688,a27690,a27692,a27694,a27696,a27700,a27702,a27704,a27706,
a27708,a27710,a27712,a27714,a27716,a27718,a27720,a27722,a27724,a27726,a27728,a27730,a27732,a27736,a27738,
a27740,a27742,a27744,a27746,a27748,a27750,a27752,a27754,a27756,a27758,a27760,a27762,a27764,a27766,a27770,
a27772,a27774,a27776,a27778,a27780,a27782,a27784,a27786,a27788,a27792,a27794,a27796,a27798,a27800,a27804,
a27806,a27808,a27810,a27812,a27814,a27816,a27818,a27820,a27822,a27824,a27826,a27828,a27830,a27832,a27834,
a27836,a27840,a27842,a27844,a27846,a27848,a27850,a27852,a27854,a27856,a27858,a27860,a27862,a27864,a27866,
a27868,a27870,a27874,a27876,a27878,a27880,a27882,a27884,a27886,a27888,a27892,a27894,a27896,a27898,a27900,
a27904,a27906,a27908,a27910,a27912,a27914,a27916,a27918,a27920,a27922,a27924,a27926,a27928,a27930,a27932,
a27934,a27936,a27940,a27942,a27944,a27946,a27948,a27950,a27952,a27954,a27956,a27958,a27960,a27962,a27964,
a27966,a27968,a27970,a27974,a27976,a27978,a27980,a27982,a27984,a27986,a27988,a27990,a27992,a27994,a27996,
a27998,a28000,a28002,a28006,a28008,a28010,a28012,a28014,a28016,a28018,a28020,a28022,a28024,a28026,a28028,
a28030,a28032,a28034,a28036,a28038,a28040,a28042,a28044,a28046,a28048,a28050,a28052,a28054,a28056,a28058,
a28060,a28062,a28064,a28066,a28068,a28070,a28074,a28076,a28078,a28080,a28084,a28086,a28088,a28090,a28092,
a28094,a28096,a28098,a28100,a28102,a28104,a28106,a28108,a28110,a28112,a28114,a28116,a28118,a28120,a28122,
a28124,a28126,a28128,a28130,a28132,a28134,a28136,a28138,a28140,a28142,a28144,a28146,a28148,a28150,a28152,
a28154,a28156,a28158,a28160,a28162,a28164,a28166,a28168,a28170,a28172,a28174,a28176,a28178,a28180,a28182,
a28184,a28186,a28188,a28190,a28192,a28194,a28196,a28198,a28200,a28202,a28204,a28206,a28208,a28210,a28212,
a28214,a28216,a28218,a28220,a28222,a28224,a28226,a28228,a28232,a28234,a28236,a28238,a28240,a28242,a28244,
a28246,a28248,a28250,a28252,a28256,a28258,a28260,a28262,a28264,a28266,a28268,a28270,a28272,a28274,a28276,
a28280,a28282,a28284,a28286,a28288,a28290,a28292,a28294,a28296,a28298,a28300,a28304,a28306,a28308,a28310,
a28312,a28316,a28318,a28322,a28324,a28328,a28330,a28334,a28336,a28340,a28342,a28346,a28348,a28352,a28354,
a28358,a28360,a28364,a28366,a28370,a28372,a28374,a28376,a28378,a28382,a28384,a28388,a28390,a28394,a28396,
a28400,a28402,a28406,a28408,a28412,a28414,a28418,a28420,a28424,a28426,a28430,a28432,a28436,a28438,a28440,
a28442,a28444,a28448,a28450,a28454,a28456,a28460,a28462,a28466,a28468,a28472,a28474,a28478,a28480,a28484,
a28486,a28490,a28492,a28496,a28498,a28502,a28504,a28506,a28508,a28510,a28514,a28516,a28520,a28522,a28526,
a28528,a28532,a28534,a28538,a28540,a28544,a28546,a28550,a28552,a28556,a28558,a28562,a28564,a28568,a28570,
a28572,a28574,a28576,a28580,a28582,a28586,a28588,a28592,a28594,a28598,a28600,a28604,a28606,a28610,a28612,
a28616,a28618,a28622,a28624,a28628,a28630,a28634,a28636,a28638,a28640,a28642,a28646,a28648,a28652,a28654,
a28658,a28660,a28664,a28666,a28670,a28672,a28676,a28678,a28682,a28684,a28688,a28690,a28694,a28696,a28700,
a28702,a28704,a28706,a28708,a28712,a28714,a28718,a28720,a28724,a28726,a28730,a28732,a28736,a28738,a28742,
a28744,a28748,a28750,a28754,a28756,a28760,a28762,a28766,a28768,a28770,a28772,a28774,a28778,a28780,a28784,
a28786,a28790,a28792,a28796,a28798,a28802,a28804,a28808,a28810,a28814,a28816,a28820,a28822,a28826,a28828,
a28832,a28836,a28838,a28840,a28842,a28844,a28846,a28848,a28850,a28852,a28854,a28856,a28858,a28860,a28862,
a28864,a28868,a28870,a28872,a28874,a28876,a28880,a28884,a28886,a28890,a28892,a28896,a28898,a28902,a28904,
a28908,a28910,a28914,a28916,a28920,a28922,a28926,a28928,a28930,a28932,a28934,a28936,a28940,a28944,a28946,
a28948,a28950,a28952,a28954,a28956,a28958,a28960,a28962,a28964,a28966,a28968,a28970,a28974,a28976,a28978,
a28980,a28982,a28984,a28986,a28988,a28990,a28992,a28994,a28996,a28998,a29000,a29002,a29004,a29006,a29008,
a29010,a29012,a29014,a29016,a29018,a29020,a29022,a29024,a29026,a29028,a29030,a29032,a29034,a29036,a29038,
a29040,a29042,a29044,a29046,a29048,a29050,a29052,a29054,a29056,a29060,a29062,a29064,a29066,a29068,a29070,
a29074,a29076,a29078,a29080,a29082,a29086,a29088,a29090,a29092,a29094,a29098,a29100,a29104,a29106,a29110,
a29112,a29116,a29118,a29124,a29126,a29128,a29130,a29134,a29136,a29138,a29140,a29142,a29146,a29148,a29150,
a29152,a29156,a29158,a29162,a29164,a29166,a29168,a29172,a29174,a29176,a29178,a29182,a29184,a29186,a29188,
a29192,a29194,a29196,a29198,a29202,a29204,a29206,a29208,a29212,a29214,a29216,a29218,a29222,a29224,a29226,
a29228,a29232,a29234,a29236,a29238,a29242,a29244,a29246,a29250,a29252,a29256,a29258,a29260,a29264,a29266,
a29268,a29272,a29274,a29276,a29278,a29280,a29282,a29284,a29286,a29288,a29290,a29292,a29294,a29296,a29298,
a29300,a29302,a29304,a29306,a29308,a29310,a29312,a29314,a29316,a29318,a29320,a29322,a29324,a29326,a29328,
a29330,a29332,a29334,a29336,a29338,a29342,a29344,a29346,a29348,a29350,a29352,a29354,a29356,a29358,a29360,
a29362,a29364,a29366,a29368,a29370,a29372,a29374,a29376,a29378,a29380,a29382,a29384,a29386,a29388,a29392,
a29394,a29396,a29398,a29400,a29402,a29404,a29406,a29410,a29412,a29414,a29416,a29418,a29420,a29422,a29424,
a29428,a29430,a29432,a29434,a29436,a29438,a29442,a29444,a29446,a29448,a29450,a29452,a29454,a29456,a29458,
a29460,a29462,a29464,a29466,a29468,a29470,a29472,a29474,a29476,a29478,a29480,a29482,a29484,a29486,a29488,
a29490,a29492,a29494,a29496,a29498,a29500,a29502,a29504,a29506,a29508,a29510,a29512,a29514,a29516,a29518,
a29520,a29522,a29524,a29526,a29528,a29530,a29532,a29534,a29536,a29538,a29540,a29542,a29544,a29546,a29548,
a29550,a29552,a29554,a29556,a29558,a29560,a29562,a29564,a29566,a29568,a29570,a29572,a29574,a29576,a29578,
a29580,a29582,a29584,a29586,a29588,a29590,a29592,a29594,a29596,a29598,a29600,a29602,a29604,a29606,a29608,
a29610,a29612,a29614,a29616,a29618,a29620,a29622,a29624,a29626,a29628,a29630,a29632,a29634,a29636,a29638,
a29640,a29642,a29644,a29646,a29648,a29650,a29652,a29654,a29656,a29658,a29660,a29662,a29664,a29666,a29668,
a29670,a29672,a29674,a29676,a29678,a29680,a29682,a29684,a29686,a29688,a29690,a29692,a29694,a29696,a29698,
a29700,a29702,a29704,a29706,a29708,a29710,a29712,a29714,a29716,a29718,a29720,a29722,a29724,a29726,a29728,
a29730,a29732,a29734,a29736,a29738,a29740,a29742,a29744,a29746,a29748,a29750,a29752,a29754,a29756,a29758,
a29760,a29762,a29764,a29766,a29768,a29770,a29772,a29774,a29776,a29778,a29780,a29782,a29784,a29786,a29788,
a29790,a29792,a29794,a29796,a29798,a29800,a29802,a29804,a29806,a29808,a29810,a29812,a29814,a29816,a29818,
a29820,a29822,a29824,a29826,a29828,a29830,a29832,a29834,a29836,a29838,a29840,a29842,a29844,a29846,a29848,
a29850,a29852,a29854,a29856,a29858,a29860,a29862,a29864,a29866,a29868,a29870,a29872,a29874,a29876,a29878,
a29880,a29882,a29884,a29886,a29888,a29890,a29892,a29894,a29896,a29898,a29900,a29902,a29904,a29906,a29908,
a29910,a29912,a29914,a29916,a29918,a29920,a29922,a29924,a29926,a29928,a29930,a29932,a29934,a29936,a29938,
a29940,a29942,a29944,a29946,a29948,a29950,a29952,a29954,a29956,a29958,a29960,a29962,a29964,a29966,a29968,
a29970,a29972,a29974,a29976,a29978,a29980,a29982,a29984,a29986,a29988,a29990,a29992,a29994,a29996,a29998,
a30000,a30002,a30004,a30006,a30008,a30010,a30012,a30014,a30016,a30018,a30020,a30022,a30024,a30026,a30028,
a30030,a30032,a30034,a30036,a30038,a30040,a30042,a30044,a30046,a30048,a30050,a30052,a30054,a30056,a30058,
a30060,a30062,a30064,a30066,a30068,a30070,a30072,a30074,a30076,a30078,a30080,a30082,a30084,a30086,a30088,
a30090,a30092,a30094,a30096,a30098,a30100,a30102,a30104,a30106,a30108,a30110,a30112,a30114,a30116,a30118,
a30120,a30122,a30124,a30126,a30128,a30130,a30132,a30134,a30136,a30138,a30140,a30142,a30144,a30146,a30148,
a30150,a30152,a30154,a30156,a30158,a30160,a30162,a30164,a30166,a30168,a30170,a30172,a30174,a30176,a30178,
a30180,a30182,a30184,a30186,a30188,a30190,a30192,a30194,a30196,a30198,a30200,a30202,a30204,a30206,a30208,
a30210,a30212,a30214,a30216,a30218,a30220,a30222,a30224,a30226,a30228,a30230,a30232,a30234,a30236,a30238,
a30240,a30242,a30244,a30246,a30248,a30250,a30252,a30254,a30256,a30258,a30260,a30262,a30264,a30266,a30268,
a30270,a30272,a30274,a30276,a30278,a30280,a30282,a30284,a30286,a30288,a30290,a30292,a30294,a30296,a30298,
a30300,a30302,a30304,a30306,a30308,a30310,a30312,a30314,a30316,a30320,a30322,a30324,a30326,a30328,a30330,
a30332,a30334,a30336,a30338,a30340,a30342,a30344,a30346,a30348,a30350,a30354,a30356,a30358,a30360,a30362,
a30364,a30368,a30370,a30372,a30374,a30376,a30378,a30380,a30382,a30386,a30388,a30390,a30394,a30396,a30398,
a30400,a30402,a30404,a30406,a30408,a30412,a30414,a30418,a30420,a30422,a30424,a30426,a30430,a30432,a30436,
a30438,a30440,a30442,a30444,a30446,a30448,a30450,a30452,a30454,a30456,a30458,a30460,a30462,a30464,a30466,
a30470,a30472,a30474,a30476,a30478,a30480,a30484,a30486,a30488,a30492,a30494,a30498,a30500,a30502,a30504,
a30508,a30510,a30512,a30514,a30516,a30518,a30520,a30522,a30524,a30526,a30528,a30530,a30532,a30534,a30536,
a30538,a30540,a30542,a30544,a30546,a30548,a30550,a30552,a30554,a30556,a30558,a30560,a30562,a30564,a30566,
a30568,a30570,a30572,a30574,a30576,a30578,a30580,a30582,a30584,a30586,a30588,a30590,a30592,a30594,a30596,
a30598,a30600,a30602,a30604,a30606,a30608,a30610,a30612,a30614,a30616,a30618,a30620,a30622,a30624,a30626,
a30628,a30630,a30632,a30634,a30636,a30638,a30640,a30642,a30644,a30646,a30648,a30650,a30652,a30654,a30656,
a30658,a30660,a30662,a30664,a30666,a30668,a30670,a30672,a30674,a30676,a30678,a30680,a30682,a30684,a30686,
a30688,a30690,a30692,a30694,a30696,a30698,a30700,a30702,a30704,a30706,a30708,a30710,a30712,a30714,a30716,
a30718,a30720,a30722,a30724,a30726,a30728,a30730,a30732,a30734,a30736,a30738,a30740,a30742,a30744,a30746,
a30748,a30750,a30752,a30754,a30756,a30758,a30760,a30762,a30764,a30766,a30768,a30770,a30772,a30774,a30776,
a30778,a30780,a30782,a30784,a30786,a30788,a30790,a30792,a30794,a30796,a30798,a30800,a30802,a30804,a30806,
a30808,a30810,a30812,a30814,a30816,a30818,a30820,a30822,a30824,a30826,a30828,a30830,a30832,a30834,a30836,
a30838,a30840,a30842,a30844,a30846,a30848,a30850,a30852,a30854,a30856,a30858,a30860,a30862,a30864,a30866,
a30868,a30870,a30872,a30874,a30876,a30878,a30880,a30882,a30884,a30886,a30888,a30890,a30892,a30894,a30896,
a30898,a30900,a30902,a30904,a30906,a30908,a30910,a30912,a30914,a30916,a30918,a30920,a30922,a30924,a30926,
a30928,a30930,a30932,a30934,a30936,a30938,a30940,a30942,a30944,a30946,a30948,a30950,a30952,a30954,a30956,
a30958,a30960,a30962,a30964,a30966,a30968,a30970,a30972,a30974,a30976,a30978,a30980,a30982,a30984,a30986,
a30988,a30990,a30992,a30994,a30996,a30998,a31000,a31002,a31004,a31006,a31008,a31010,a31012,a31014,a31016,
a31018,a31020,a31022,a31024,a31026,a31028,a31030,a31032,a31034,a31036,a31038,a31040,a31042,a31044,a31046,
a31048,a31050,a31052,a31054,a31056,a31058,a31060,a31062,a31064,a31066,a31068,a31070,a31072,a31074,a31076,
a31078,a31080,a31082,a31084,a31086,a31088,a31090,a31092,a31094,a31096,a31098,a31100,a31102,a31104,a31106,
a31108,a31110,a31112,a31114,a31116,a31118,a31120,a31122,a31124,a31126,a31128,a31130,a31132,a31134,a31136,
a31138,a31140,a31142,a31144,a31146,a31148,a31150,a31152,a31154,a31156,a31158,a31160,a31162,a31164,a31166,
a31168,a31170,a31172,a31174,a31176,a31178,a31180,a31182,a31184,a31186,a31188,a31190,a31192,a31194,a31196,
a31198,a31200,a31202,a31204,a31206,a31208,a31210,a31212,a31214,a31216,a31218,a31220,a31222,a31224,a31226,
a31228,a31230,a31232,a31234,a31236,a31238,a31240,a31242,a31244,a31246,a31248,a31250,a31252,a31254,a31256,
a31258,a31260,a31262,a31264,a31266,a31268,a31270,a31272,a31274,a31276,a31278,a31280,a31282,a31284,a31286,
a31288,a31290,a31292,a31294,a31296,a31298,a31300,a31302,a31304,a31306,a31308,a31310,a31312,a31314,a31316,
a31318,a31320,a31322,a31324,a31326,a31328,a31330,a31332,a31334,a31336,a31338,a31340,a31342,a31344,a31346,
a31348,a31350,a31352,a31354,a31356,a31358,a31360,a31362,a31364,a31366,a31368,a31370,a31372,a31374,a31376,
a31378,a31380,a31382,a31384,a31386,a31388,a31390,a31392,a31394,a31396,a31398,a31400,a31402,a31404,a31406,
a31408,a31410,a31412,a31414,a31416,a31418,a31420,a31422,a31424,a31426,a31428,a31430,a31432,a31434,a31436,
a31438,a31440,a31442,a31444,a31446,a31448,a31450,a31452,a31454,a31456,a31458,a31460,a31462,a31464,a31466,
a31468,a31470,a31472,a31474,a31476,a31478,a31480,a31482,a31484,a31486,a31488,a31490,a31492,a31494,a31496,
a31498,a31500,a31502,a31504,a31506,a31508,a31510,a31512,a31514,a31516,a31518,a31520,a31522,a31524,a31526,
a31528,a31530,a31532,a31534,a31536,a31538,a31540,a31542,a31544,a31546,a31548,a31550,a31552,a31554,a31556,
a31558,a31560,a31562,a31564,a31566,a31568,a31570,a31572,a31574,a31576,a31578,a31580,a31582,a31584,a31586,
a31588,a31590,a31592,a31594,a31596,a31598,a31600,a31602,a31604,a31606,a31608,a31610,a31612,a31614,a31616,
a31618,a31620,a31622,a31624,a31626,a31628,a31630,a31632,a31634,a31636,a31638,a31640,a31642,a31644,a31646,
a31648,a31650,a31652,a31654,a31656,a31658,a31660,a31662,a31664,a31666,a31668,a31670,a31672,a31674,a31676,
a31678,a31680,a31682,a31684,a31686,a31688,a31690,a31692,a31694,a31696,a31698,a31700,a31702,a31704,a31706,
a31708,a31710,a31712,a31714,a31716,a31718,a31720,a31722,a31724,a31726,a31728,a31730,a31732,a31734,a31736,
a31738,a31740,a31742,a31744,a31746,a31748,a31750,a31752,a31754,a31756,a31758,a31760,a31762,a31764,a31766,
a31768,a31770,a31772,a31774,a31776,a31778,a31780,a31782,a31784,a31786,a31788,a31790,a31792,a31794,a31796,
a31798,a31800,a31802,a31804,a31806,a31808,a31810,a31812,a31814,a31816,a31818,a31820,a31822,a31824,a31826,
a31828,a31830,a31832,a31834,a31836,a31838,a31840,a31842,a31844,a31846,a31848,a31850,a31852,a31854,a31856,
a31858,a31860,a31862,a31864,a31866,a31868,a31870,a31872,a31874,a31876,a31878,a31880,a31882,a31884,a31886,
a31888,a31890,a31892,a31894,a31896,a31898,a31900,a31902,a31904,a31906,a31908,a31910,a31912,a31914,a31916,
a31918,a31920,a31922,a31924,a31926,a31928,a31930,a31932,a31934,a31936,a31938,a31940,a31942,a31944,a31946,
a31948,a31950,a31952,a31954,a31956,a31958,a31960,a31962,a31964,a31966,a31968,a31970,a31972,a31974,a31976,
a31978,a31980,a31982,a31984,a31986,a31988,a31990,a31992,a31994,a31996,a31998,a32000,a32002,a32004,a32006,
a32008,a32010,a32012,a32014,a32016,a32018,a32020,a32022,a32024,a32026,a32030,a32032,a32034,a32036,a32038,
a32040,a32042,a32044,a32046,a32048,a32050,a32052,a32054,a32056,a32058,a32060,a32062,a32064,a32066,a32068,
a32070,a32072,a32074,a32076,a32078,a32080,a32082,a32084,a32086,a32088,a32090,a32092,a32094,a32096,a32098,
a32100,a32102,a32104,a32106,a32108,a32110,a32112,a32114,a32116,a32118,a32120,a32122,a32124,a32126,a32128,
a32130,a32132,a32134,a32136,a32138,a32140,a32142,a32144,a32146,a32148,a32150,a32152,a32154,a32156,a32158,
a32160,a32162,a32164,a32166,a32168,a32170,a32172,a32174,a32176,a32178,a32180,a32182,a32184,a32186,a32188,
a32190,a32192,a32194,a32196,a32198,a32200,a32202,a32204,a32206,a32208,a32210,a32212,a32214,a32216,a32218,
a32220,a32222,a32224,a32226,a32228,a32230,a32232,a32234,a32236,a32238,a32240,a32242,a32244,a32246,a32248,
a32250,a32252,a32254,a32256,a32258,a32260,a32262,a32264,a32266,a32268,a32270,a32272,a32274,a32276,a32278,
a32280,a32282,a32284,a32286,a32288,a32290,a32292,a32294,a32296,a32298,a32300,a32302,a32304,a32306,a32308,
a32310,a32312,a32314,a32316,a32318,a32320,a32322,a32324,a32326,a32328,a32330,a32332,a32334,a32336,a32338,
a32340,a32342,a32344,a32346,a32348,a32350,a32352,a32354,a32356,a32358,a32360,a32362,a32364,a32366,a32368,
a32370,a32372,a32374,a32376,a32378,a32380,a32382,a32384,a32386,a32388,a32390,a32392,a32394,a32396,a32398,
a32400,a32402,a32404,a32406,a32408,a32410,a32412,a32414,a32416,a32418,a32420,a32422,a32424,a32426,a32428,
a32430,a32432,a32434,a32436,a32438,a32440,a32442,a32444,a32446,a32448,a32450,a32452,a32454,a32456,a32458,
a32460,a32462,a32464,a32466,a32468,a32470,a32472,a32474,a32476,a32478,a32480,a32482,a32484,a32486,a32488,
a32490,a32492,a32494,a32496,a32498,a32500,a32502,a32504,a32506,a32508,a32510,a32512,a32514,a32516,a32518,
a32520,a32522,a32524,a32526,a32528,a32530,a32532,a32534,a32536,a32538,a32540,a32542,a32544,a32546,a32550,
a32552,a32554,a32556,a32558,a32560,a32562,p0;

reg l492,l494,l496,l498,l500,l502,l504,l506,l508,l510,l512,l514,l516,l518,l520,
l522,l524,l526,l528,l530,l532,l534,l536,l538,l540,l542,l544,l546,l548,l550,
l552,l554,l556,l558,l560,l562,l564,l566,l568,l570,l572,l574,l576,l578,l580,
l582,l584,l586,l588,l590,l592,l594,l596,l598,l600,l602,l604,l606,l608,l610,
l612,l614,l616,l618,l620,l622,l624,l626,l628,l630,l632,l634,l636,l638,l640,
l642,l644,l646,l648,l650,l652,l654,l656,l658,l660,l662,l664,l666,l668,l670,
l672,l674,l676,l678,l680,l682,l684,l686,l688,l690,l692,l694,l696,l698,l700,
l702,l704,l706,l708,l710,l712,l714,l716,l718,l720,l722,l724,l726,l728,l730,
l732,l734,l736,l738,l740,l742,l744,l746,l748,l750,l752,l754,l756,l758,l760,
l762,l764,l766,l768,l770,l772,l774,l776,l778,l780,l782,l784,l786,l788,l790,
l792,l794,l796,l798,l800,l802,l804,l806,l808,l810,l812,l814,l816,l818,l820,
l822,l824,l826,l828,l830,l832,l834,l836,l838,l840,l842,l844,l846,l848,l850,
l852,l854,l856,l858,l860,l862,l864,l866,l868,l870,l872,l874,l876,l878,l880,
l882,l884,l886,l888,l890,l892,l894,l896,l898,l900,l902,l904,l906,l908,l910,
l912,l914,l916,l918,l920,l922,l924,l926,l928,l930,l932,l934,l936,l938,l940,
l942,l944,l946,l948,l950,l952,l954,l956,l958,l960,l962,l964,l966,l968,l970,
l972,l974,l976,l978,l980,l982,l984,l986,l988,l990,l992,l994,l996,l998,l1000,
l1002,l1004,l1006,l1008,l1010,l1012,l1014,l1016,l1018,l1020,l1022,l1024,l1026,l1028,l1030,
l1032,l1034,l1036,l1038,l1040,l1042,l1044,l1046,l1048,l1050,l1052,l1054,l1056,l1058,l1060,
l1062,l1064,l1066,l1068,l1070,l1072,l1074,l1076,l1078,l1080,l1082,l1084,l1086,l1088,l1090,
l1092,l1094,l1096,l1098,l1100,l1102,l1104,l1106,l1108,l1110,l1112,l1114,l1116,l1118,l1120,
l1122,l1124,l1126,l1128,l1130,l1132,l1134,l1136,l1138,l1140,l1142,l1144,l1146,l1148,l1150,
l1152,l1154,l1156,l1158,l1160,l1162,l1164,l1166,l1168,l1170,l1172,l1174,l1176,l1178,l1180,
l1182,l1184,l1186,l1188,l1190,l1192,l1194,l1196,l1198,l1200,l1202,l1204,l1206,l1208,l1210,
l1212,l1214,l1216,l1218,l1220,l1222,l1224,l1226,l1228,l1230,l1232,l1234,l1236,l1238,l1240,
l1242,l1244,l1246,l1248,l1250,l1252,l1254,l1256,l1258,l1260,l1262,l1264,l1266,l1268,l1270,
l1272,l1274,l1276,l1278,l1280,l1282,l1284,l1286,l1288,l1290,l1292,l1294,l1296,l1298,l1300,
l1302,l1304,l1306,l1308,l1310,l1312,l1314,l1316,l1318,l1320,l1322,l1324,l1326,l1328,l1330,
l1332,l1334,l1336,l1338,l1340,l1342,l1344,l1346,l1348,l1350,l1352,l1354,l1356,l1358,l1360,
l1362,l1364,l1366,l1368,l1370,l1372,l1374,l1376,l1378,l1380,l1382,l1384,l1386,l1388,l1390,
l1392,l1394,l1396,l1398,l1400,l1402,l1404,l1406,l1408,l1410,l1412,l1414,l1416,l1418,l1420,
l1422,l1424,l1426,l1428,l1430,l1432,l1434,l1436,l1438,l1440,l1442,l1444,l1446,l1448,l1450,
l1452,l1454,l1456,l1458,l1460,l1462,l1464,l1466,l1468,l1470,l1472,l1474,l1476,l1478,l1480,
l1482,l1484,l1486,l1488,l1490,l1492,l1494,l1496,l1498,l1500,l1502,l1504,l1506,l1508,l1510,
l1512,l1514,l1516,l1518,l1520,l1522,l1524,l1526,l1528,l1530,l1532,l1534,l1536,l1538,l1540,
l1542,l1544,l1546,l1548,l1550,l1552,l1554,l1556,l1558,l1560,l1562,l1564,l1566,l1568,l1570,
l1572,l1574,l1576,l1578,l1580,l1582,l1584,l1586,l1588,l1590,l1592,l1594,l1596,l1598,l1600,
l1602,l1604,l1606,l1608,l1610,l1612,l1614,l1616,l1618,l1620,l1622,l1624,l1626,l1628,l1630,
l1632,l1634,l1636,l1638,l1640,l1642,l1644,l1646,l1648,l1650,l1652,l1654,l1656,l1658,l1660,
l1662,l1664,l1666,l1668,l1670,l1672,l1674,l1676,l1678,l1680,l1682,l1684,l1686;

initial
begin
   l492 = 0;
   l494 = 0;
   l496 = 0;
   l498 = 0;
   l500 = 0;
   l502 = 0;
   l504 = 0;
   l506 = 0;
   l508 = 0;
   l510 = 0;
   l512 = 0;
   l514 = 0;
   l516 = 0;
   l518 = 0;
   l520 = 0;
   l522 = 0;
   l524 = 0;
   l526 = 0;
   l528 = 0;
   l530 = 0;
   l532 = 0;
   l534 = 0;
   l536 = 0;
   l538 = 0;
   l540 = 0;
   l542 = 0;
   l544 = 0;
   l546 = 0;
   l548 = 0;
   l550 = 0;
   l552 = 0;
   l554 = 0;
   l556 = 0;
   l558 = 0;
   l560 = 0;
   l562 = 0;
   l564 = 0;
   l566 = 0;
   l568 = 0;
   l570 = 0;
   l572 = 0;
   l574 = 0;
   l576 = 0;
   l578 = 0;
   l580 = 0;
   l582 = 0;
   l584 = 0;
   l586 = 0;
   l588 = 0;
   l590 = 0;
   l592 = 0;
   l594 = 0;
   l596 = 0;
   l598 = 0;
   l600 = 0;
   l602 = 0;
   l604 = 0;
   l606 = 0;
   l608 = 0;
   l610 = 0;
   l612 = 0;
   l614 = 0;
   l616 = 0;
   l618 = 0;
   l620 = 0;
   l622 = 0;
   l624 = 0;
   l626 = 0;
   l628 = 0;
   l630 = 0;
   l632 = 0;
   l634 = 0;
   l636 = 0;
   l638 = 0;
   l640 = 0;
   l642 = 0;
   l644 = 0;
   l646 = 0;
   l648 = 0;
   l650 = 0;
   l652 = 0;
   l654 = 0;
   l656 = 0;
   l658 = 0;
   l660 = 0;
   l662 = 0;
   l664 = 0;
   l666 = 0;
   l668 = 0;
   l670 = 0;
   l672 = 0;
   l674 = 0;
   l676 = 0;
   l678 = 0;
   l680 = 0;
   l682 = 0;
   l684 = 0;
   l686 = 0;
   l688 = 0;
   l690 = 0;
   l692 = 0;
   l694 = 0;
   l696 = 0;
   l698 = 0;
   l700 = 0;
   l702 = 0;
   l704 = 0;
   l706 = 0;
   l708 = 0;
   l710 = 0;
   l712 = 0;
   l714 = 0;
   l716 = 0;
   l718 = 0;
   l720 = 0;
   l722 = 0;
   l724 = 0;
   l726 = 0;
   l728 = 0;
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
   l802 = 0;
   l804 = 0;
   l806 = 0;
   l808 = 0;
   l810 = 0;
   l812 = 0;
   l814 = 0;
   l816 = 0;
   l818 = 0;
   l820 = 0;
   l822 = 0;
   l824 = 0;
   l826 = 0;
   l828 = 0;
   l830 = 0;
   l832 = 0;
   l834 = 0;
   l836 = 0;
   l838 = 0;
   l840 = 0;
   l842 = 0;
   l844 = 0;
   l846 = 0;
   l848 = 0;
   l850 = 0;
   l852 = 0;
   l854 = 0;
   l856 = 0;
   l858 = 0;
   l860 = 0;
   l862 = 0;
   l864 = 0;
   l866 = 0;
   l868 = 0;
   l870 = 0;
   l872 = 0;
   l874 = 0;
   l876 = 0;
   l878 = 0;
   l880 = 0;
   l882 = 0;
   l884 = 0;
   l886 = 0;
   l888 = 0;
   l890 = 0;
   l892 = 0;
   l894 = 0;
   l896 = 0;
   l898 = 0;
   l900 = 0;
   l902 = 0;
   l904 = 0;
   l906 = 0;
   l908 = 0;
   l910 = 0;
   l912 = 0;
   l914 = 0;
   l916 = 0;
   l918 = 0;
   l920 = 0;
   l922 = 0;
   l924 = 0;
   l926 = 0;
   l928 = 0;
   l930 = 0;
   l932 = 0;
   l934 = 0;
   l936 = 0;
   l938 = 0;
   l940 = 0;
   l942 = 0;
   l944 = 0;
   l946 = 0;
   l948 = 0;
   l950 = 0;
   l952 = 0;
   l954 = 0;
   l956 = 0;
   l958 = 0;
   l960 = 0;
   l962 = 0;
   l964 = 0;
   l966 = 0;
   l968 = 0;
   l970 = 0;
   l972 = 0;
   l974 = 0;
   l976 = 0;
   l978 = 0;
   l980 = 0;
   l982 = 0;
   l984 = 0;
   l986 = 0;
   l988 = 0;
   l990 = 0;
   l992 = 0;
   l994 = 0;
   l996 = 0;
   l998 = 0;
   l1000 = 0;
   l1002 = 0;
   l1004 = 0;
   l1006 = 0;
   l1008 = 0;
   l1010 = 0;
   l1012 = 0;
   l1014 = 0;
   l1016 = 0;
   l1018 = 0;
   l1020 = 0;
   l1022 = 0;
   l1024 = 0;
   l1026 = 0;
   l1028 = 0;
   l1030 = 0;
   l1032 = 0;
   l1034 = 0;
   l1036 = 0;
   l1038 = 0;
   l1040 = 0;
   l1042 = 0;
   l1044 = 0;
   l1046 = 0;
   l1048 = 0;
   l1050 = 0;
   l1052 = 0;
   l1054 = 0;
   l1056 = 0;
   l1058 = 0;
   l1060 = 0;
   l1062 = 0;
   l1064 = 0;
   l1066 = 0;
   l1068 = 0;
   l1070 = 0;
   l1072 = 0;
   l1074 = 0;
   l1076 = 0;
   l1078 = 0;
   l1080 = 0;
   l1082 = 0;
   l1084 = 0;
   l1086 = 0;
   l1088 = 0;
   l1090 = 0;
   l1092 = 0;
   l1094 = 0;
   l1096 = 0;
   l1098 = 0;
   l1100 = 0;
   l1102 = 0;
   l1104 = 0;
   l1106 = 0;
   l1108 = 0;
   l1110 = 0;
   l1112 = 0;
   l1114 = 0;
   l1116 = 0;
   l1118 = 0;
   l1120 = 0;
   l1122 = 0;
   l1124 = 0;
   l1126 = 0;
   l1128 = 0;
   l1130 = 0;
   l1132 = 0;
   l1134 = 0;
   l1136 = 0;
   l1138 = 0;
   l1140 = 0;
   l1142 = 0;
   l1144 = 0;
   l1146 = 0;
   l1148 = 0;
   l1150 = 0;
   l1152 = 0;
   l1154 = 0;
   l1156 = 0;
   l1158 = 0;
   l1160 = 0;
   l1162 = 0;
   l1164 = 0;
   l1166 = 0;
   l1168 = 0;
   l1170 = 0;
   l1172 = 0;
   l1174 = 0;
   l1176 = 0;
   l1178 = 0;
   l1180 = 0;
   l1182 = 0;
   l1184 = 0;
   l1186 = 0;
   l1188 = 0;
   l1190 = 0;
   l1192 = 0;
   l1194 = 0;
   l1196 = 0;
   l1198 = 0;
   l1200 = 0;
   l1202 = 0;
   l1204 = 0;
   l1206 = 0;
   l1208 = 0;
   l1210 = 0;
   l1212 = 0;
   l1214 = 0;
   l1216 = 0;
   l1218 = 0;
   l1220 = 0;
   l1222 = 0;
   l1224 = 0;
   l1226 = 0;
   l1228 = 0;
   l1230 = 0;
   l1232 = 0;
   l1234 = 0;
   l1236 = 0;
   l1238 = 0;
   l1240 = 0;
   l1242 = 0;
   l1244 = 0;
   l1246 = 0;
   l1248 = 0;
   l1250 = 0;
   l1252 = 0;
   l1254 = 0;
   l1256 = 0;
   l1258 = 0;
   l1260 = 0;
   l1262 = 0;
   l1264 = 0;
   l1266 = 0;
   l1268 = 0;
   l1270 = 0;
   l1272 = 0;
   l1274 = 0;
   l1276 = 0;
   l1278 = 0;
   l1280 = 0;
   l1282 = 0;
   l1284 = 0;
   l1286 = 0;
   l1288 = 0;
   l1290 = 0;
   l1292 = 0;
   l1294 = 0;
   l1296 = 0;
   l1298 = 0;
   l1300 = 0;
   l1302 = 0;
   l1304 = 0;
   l1306 = 0;
   l1308 = 0;
   l1310 = 0;
   l1312 = 0;
   l1314 = 0;
   l1316 = 0;
   l1318 = 0;
   l1320 = 0;
   l1322 = 0;
   l1324 = 0;
   l1326 = 0;
   l1328 = 0;
   l1330 = 0;
   l1332 = 0;
   l1334 = 0;
   l1336 = 0;
   l1338 = 0;
   l1340 = 0;
   l1342 = 0;
   l1344 = 0;
   l1346 = 0;
   l1348 = 0;
   l1350 = 0;
   l1352 = 0;
   l1354 = 0;
   l1356 = 0;
   l1358 = 0;
   l1360 = 0;
   l1362 = 0;
   l1364 = 0;
   l1366 = 0;
   l1368 = 0;
   l1370 = 0;
   l1372 = 0;
   l1374 = 0;
   l1376 = 0;
   l1378 = 0;
   l1380 = 0;
   l1382 = 0;
   l1384 = 0;
   l1386 = 0;
   l1388 = 0;
   l1390 = 0;
   l1392 = 0;
   l1394 = 0;
   l1396 = 0;
   l1398 = 0;
   l1400 = 0;
   l1402 = 0;
   l1404 = 0;
   l1406 = 0;
   l1408 = 0;
   l1410 = 0;
   l1412 = 0;
   l1414 = 0;
   l1416 = 0;
   l1418 = 0;
   l1420 = 0;
   l1422 = 0;
   l1424 = 0;
   l1426 = 0;
   l1428 = 0;
   l1430 = 0;
   l1432 = 0;
   l1434 = 0;
   l1436 = 0;
   l1438 = 0;
   l1440 = 0;
   l1442 = 0;
   l1444 = 0;
   l1446 = 0;
   l1448 = 0;
   l1450 = 0;
   l1452 = 0;
   l1454 = 0;
   l1456 = 0;
   l1458 = 0;
   l1460 = 0;
   l1462 = 0;
   l1464 = 0;
   l1466 = 0;
   l1468 = 0;
   l1470 = 0;
   l1472 = 0;
   l1474 = 0;
   l1476 = 0;
   l1478 = 0;
   l1480 = 0;
   l1482 = 0;
   l1484 = 0;
   l1486 = 0;
   l1488 = 0;
   l1490 = 0;
   l1492 = 0;
   l1494 = 0;
   l1496 = 0;
   l1498 = 0;
   l1500 = 0;
   l1502 = 0;
   l1504 = 0;
   l1506 = 0;
   l1508 = 0;
   l1510 = 0;
   l1512 = 0;
   l1514 = 0;
   l1516 = 0;
   l1518 = 0;
   l1520 = 0;
   l1522 = 0;
   l1524 = 0;
   l1526 = 0;
   l1528 = 0;
   l1530 = 0;
   l1532 = 0;
   l1534 = 0;
   l1536 = 0;
   l1538 = 0;
   l1540 = 0;
   l1542 = 0;
   l1544 = 0;
   l1546 = 0;
   l1548 = 0;
   l1550 = 0;
   l1552 = 0;
   l1554 = 0;
   l1556 = 0;
   l1558 = 0;
   l1560 = 0;
   l1562 = 0;
   l1564 = 0;
   l1566 = 0;
   l1568 = 0;
   l1570 = 0;
   l1572 = 0;
   l1574 = 0;
   l1576 = 0;
   l1578 = 0;
   l1580 = 0;
   l1582 = 0;
   l1584 = 0;
   l1586 = 0;
   l1588 = 0;
   l1590 = 0;
   l1592 = 0;
   l1594 = 0;
   l1596 = 0;
   l1598 = 0;
   l1600 = 0;
   l1602 = 0;
   l1604 = 0;
   l1606 = 0;
   l1608 = 0;
   l1610 = 0;
   l1612 = 0;
   l1614 = 0;
   l1616 = 0;
   l1618 = 0;
   l1620 = 0;
   l1622 = 0;
   l1624 = 0;
   l1626 = 0;
   l1628 = 0;
   l1630 = 0;
   l1632 = 0;
   l1634 = 0;
   l1636 = 0;
   l1638 = 0;
   l1640 = 0;
   l1642 = 0;
   l1644 = 0;
   l1646 = 0;
   l1648 = 0;
   l1650 = 0;
   l1652 = 0;
   l1654 = 0;
   l1656 = 0;
   l1658 = 0;
   l1660 = 0;
   l1662 = 0;
   l1664 = 0;
   l1666 = 0;
   l1668 = 0;
   l1670 = 0;
   l1672 = 0;
   l1674 = 0;
   l1676 = 0;
   l1678 = 0;
   l1680 = 0;
   l1682 = 0;
   l1684 = 0;
   l1686 = 0;
end

always @(posedge a6662)
   l492 <= a6662;

always @(posedge a6682)
   l494 <= a6682;

always @(posedge a6690)
   l496 <= a6690;

always @(posedge a6696)
   l498 <= a6696;

always @(posedge a6702)
   l500 <= a6702;

always @(posedge a6708)
   l502 <= a6708;

always @(posedge na6710)
   l504 <= na6710;

always @(posedge l1684)
   l506 <= l1684;

always @(posedge l510)
   l508 <= l510;

always @(posedge l514)
   l510 <= l514;

always @(posedge a6712)
   l512 <= a6712;

always @(posedge l966)
   l514 <= l966;

always @(posedge l1678)
   l516 <= l1678;

always @(posedge a6074)
   l518 <= a6074;

always @(posedge a6920)
   l520 <= a6920;

always @(posedge a7152)
   l522 <= a7152;

always @(posedge a7352)
   l524 <= a7352;

always @(posedge a7590)
   l526 <= a7590;

always @(posedge a7812)
   l528 <= a7812;

always @(posedge a7852)
   l530 <= a7852;

always @(posedge a7864)
   l532 <= a7864;

always @(posedge a7900)
   l534 <= a7900;

always @(posedge a7930)
   l536 <= a7930;

always @(posedge a7942)
   l538 <= a7942;

always @(posedge a7954)
   l540 <= a7954;

always @(posedge a7966)
   l542 <= a7966;

always @(posedge a7978)
   l544 <= a7978;

always @(posedge a7990)
   l546 <= a7990;

always @(posedge a8002)
   l548 <= a8002;

always @(posedge a8020)
   l550 <= a8020;

always @(posedge a16268)
   l552 <= a16268;

always @(posedge a16274)
   l554 <= a16274;

always @(posedge a16280)
   l556 <= a16280;

always @(posedge a16286)
   l558 <= a16286;

always @(posedge a16292)
   l560 <= a16292;

always @(posedge a16298)
   l562 <= a16298;

always @(posedge a16304)
   l564 <= a16304;

always @(posedge a16310)
   l566 <= a16310;

always @(posedge a16660)
   l568 <= a16660;

always @(posedge a16800)
   l570 <= a16800;

always @(posedge a16936)
   l572 <= a16936;

always @(posedge a17072)
   l574 <= a17072;

always @(posedge a17208)
   l576 <= a17208;

always @(posedge a17342)
   l578 <= a17342;

always @(posedge a17476)
   l580 <= a17476;

always @(posedge a17610)
   l582 <= a17610;

always @(posedge a17742)
   l584 <= a17742;

always @(posedge a17872)
   l586 <= a17872;

always @(posedge a15370)
   l588 <= a15370;

always @(posedge a15474)
   l590 <= a15474;

always @(posedge a15578)
   l592 <= a15578;

always @(posedge a15682)
   l594 <= a15682;

always @(posedge a15786)
   l596 <= a15786;

always @(posedge a15884)
   l598 <= a15884;

always @(posedge a15982)
   l600 <= a15982;

always @(posedge na2430)
   l602 <= na2430;

always @(posedge a17882)
   l604 <= a17882;

always @(posedge na2432)
   l606 <= na2432;

always @(posedge na2436)
   l608 <= na2436;

always @(posedge a17900)
   l610 <= a17900;

always @(posedge a17916)
   l612 <= a17916;

always @(posedge na2434)
   l614 <= na2434;

always @(posedge na5594)
   l616 <= na5594;

always @(posedge na5596)
   l618 <= na5596;

always @(posedge na5600)
   l620 <= na5600;

always @(posedge na5598)
   l622 <= na5598;

always @(posedge a6592)
   l624 <= a6592;

always @(posedge a6476)
   l626 <= a6476;

always @(posedge a6548)
   l628 <= a6548;

always @(posedge a6512)
   l630 <= a6512;

always @(posedge na17918)
   l632 <= na17918;

always @(posedge na17920)
   l634 <= na17920;

always @(posedge na17922)
   l636 <= na17922;

always @(posedge na17924)
   l638 <= na17924;

always @(posedge a15314)
   l640 <= a15314;

always @(posedge a6522)
   l642 <= a6522;

always @(posedge a6566)
   l644 <= a6566;

always @(posedge a6608)
   l646 <= a6608;

always @(posedge a6494)
   l648 <= a6494;

always @(posedge a18026)
   l650 <= a18026;

always @(posedge na18028)
   l652 <= na18028;

always @(posedge na6410)
   l654 <= na6410;

always @(posedge na6404)
   l656 <= na6404;

always @(posedge a6424)
   l658 <= a6424;

always @(posedge a6448)
   l660 <= a6448;

always @(posedge a18098)
   l662 <= a18098;

always @(posedge z0)
   l664 <= z0;

always @(posedge a19208)
   l666 <= a19208;

always @(posedge a19248)
   l668 <= a19248;

always @(posedge a19262)
   l670 <= a19262;

always @(posedge a19274)
   l672 <= a19274;

always @(posedge a19282)
   l674 <= a19282;

always @(posedge a19292)
   l676 <= a19292;

always @(posedge a19300)
   l678 <= a19300;

always @(posedge a19308)
   l680 <= a19308;

always @(posedge a19318)
   l682 <= a19318;

always @(posedge a19326)
   l684 <= a19326;

always @(posedge a19334)
   l686 <= a19334;

always @(posedge a19342)
   l688 <= a19342;

always @(posedge a19348)
   l690 <= a19348;

always @(posedge a19354)
   l692 <= a19354;

always @(posedge a19360)
   l694 <= a19360;

always @(posedge a19336)
   l696 <= a19336;

always @(posedge na16352)
   l698 <= na16352;

always @(posedge na19362)
   l700 <= na19362;

always @(posedge a6346)
   l702 <= a6346;

always @(posedge a19364)
   l704 <= a19364;

always @(posedge a19924)
   l706 <= a19924;

always @(posedge a19912)
   l708 <= a19912;

always @(posedge a19834)
   l710 <= a19834;

always @(posedge a19808)
   l712 <= a19808;

always @(posedge a19770)
   l714 <= a19770;

always @(posedge a19732)
   l716 <= a19732;

always @(posedge a19698)
   l718 <= a19698;

always @(posedge a19664)
   l720 <= a19664;

always @(posedge a19630)
   l722 <= a19630;

always @(posedge a19926)
   l724 <= a19926;

always @(posedge a19938)
   l726 <= a19938;

always @(posedge a19944)
   l728 <= a19944;

always @(posedge a19950)
   l730 <= a19950;

always @(posedge a19956)
   l732 <= a19956;

always @(posedge a19962)
   l734 <= a19962;

always @(posedge a19968)
   l736 <= a19968;

always @(posedge a19974)
   l738 <= a19974;

always @(posedge a19980)
   l740 <= a19980;

always @(posedge a19986)
   l742 <= a19986;

always @(posedge a19992)
   l744 <= a19992;

always @(posedge a16070)
   l746 <= a16070;

always @(posedge a20004)
   l748 <= a20004;

always @(posedge a20010)
   l750 <= a20010;

always @(posedge a20016)
   l752 <= a20016;

always @(posedge a20022)
   l754 <= a20022;

always @(posedge a20028)
   l756 <= a20028;

always @(posedge a20034)
   l758 <= a20034;

always @(posedge a20040)
   l760 <= a20040;

always @(posedge a20046)
   l762 <= a20046;

always @(posedge a20052)
   l764 <= a20052;

always @(posedge a20058)
   l766 <= a20058;

always @(posedge a20060)
   l768 <= a20060;

always @(posedge a20072)
   l770 <= a20072;

always @(posedge a20078)
   l772 <= a20078;

always @(posedge a20084)
   l774 <= a20084;

always @(posedge a20090)
   l776 <= a20090;

always @(posedge a20096)
   l778 <= a20096;

always @(posedge a20102)
   l780 <= a20102;

always @(posedge a20108)
   l782 <= a20108;

always @(posedge a20114)
   l784 <= a20114;

always @(posedge a20120)
   l786 <= a20120;

always @(posedge a20126)
   l788 <= a20126;

always @(posedge a20128)
   l790 <= a20128;

always @(posedge a20140)
   l792 <= a20140;

always @(posedge a20146)
   l794 <= a20146;

always @(posedge a20152)
   l796 <= a20152;

always @(posedge a20158)
   l798 <= a20158;

always @(posedge a20164)
   l800 <= a20164;

always @(posedge a20170)
   l802 <= a20170;

always @(posedge a20176)
   l804 <= a20176;

always @(posedge a20182)
   l806 <= a20182;

always @(posedge a20188)
   l808 <= a20188;

always @(posedge a20194)
   l810 <= a20194;

always @(posedge a20196)
   l812 <= a20196;

always @(posedge a20208)
   l814 <= a20208;

always @(posedge a20214)
   l816 <= a20214;

always @(posedge a20220)
   l818 <= a20220;

always @(posedge a20226)
   l820 <= a20226;

always @(posedge a20232)
   l822 <= a20232;

always @(posedge a20238)
   l824 <= a20238;

always @(posedge a20244)
   l826 <= a20244;

always @(posedge a20250)
   l828 <= a20250;

always @(posedge a20256)
   l830 <= a20256;

always @(posedge a20262)
   l832 <= a20262;

always @(posedge a20264)
   l834 <= a20264;

always @(posedge a20276)
   l836 <= a20276;

always @(posedge a20282)
   l838 <= a20282;

always @(posedge a20288)
   l840 <= a20288;

always @(posedge a20294)
   l842 <= a20294;

always @(posedge a20300)
   l844 <= a20300;

always @(posedge a20306)
   l846 <= a20306;

always @(posedge a20312)
   l848 <= a20312;

always @(posedge a20318)
   l850 <= a20318;

always @(posedge a20324)
   l852 <= a20324;

always @(posedge a20330)
   l854 <= a20330;

always @(posedge a20332)
   l856 <= a20332;

always @(posedge a20344)
   l858 <= a20344;

always @(posedge a20350)
   l860 <= a20350;

always @(posedge a20356)
   l862 <= a20356;

always @(posedge a20362)
   l864 <= a20362;

always @(posedge a20368)
   l866 <= a20368;

always @(posedge a20374)
   l868 <= a20374;

always @(posedge a20380)
   l870 <= a20380;

always @(posedge a20386)
   l872 <= a20386;

always @(posedge a20392)
   l874 <= a20392;

always @(posedge a20398)
   l876 <= a20398;

always @(posedge a8042)
   l878 <= a8042;

always @(posedge a20412)
   l880 <= a20412;

always @(posedge a20418)
   l882 <= a20418;

always @(posedge a20424)
   l884 <= a20424;

always @(posedge a20430)
   l886 <= a20430;

always @(posedge a20436)
   l888 <= a20436;

always @(posedge a20442)
   l890 <= a20442;

always @(posedge a20448)
   l892 <= a20448;

always @(posedge a20454)
   l894 <= a20454;

always @(posedge a20460)
   l896 <= a20460;

always @(posedge a20466)
   l898 <= a20466;

always @(posedge a20564)
   l900 <= a20564;

always @(posedge a20636)
   l902 <= a20636;

always @(posedge a20666)
   l904 <= a20666;

always @(posedge a20716)
   l906 <= a20716;

always @(posedge a20762)
   l908 <= a20762;

always @(posedge a20800)
   l910 <= a20800;

always @(posedge a20816)
   l912 <= a20816;

always @(posedge a20836)
   l914 <= a20836;

always @(posedge a20854)
   l916 <= a20854;

always @(posedge a20870)
   l918 <= a20870;

always @(posedge na20872)
   l920 <= na20872;

always @(posedge na20874)
   l922 <= na20874;

always @(posedge na20876)
   l924 <= na20876;

always @(posedge na20878)
   l926 <= na20878;

always @(posedge a6384)
   l928 <= a6384;

always @(posedge a6372)
   l930 <= a6372;

always @(posedge a6362)
   l932 <= a6362;

always @(posedge a6394)
   l934 <= a6394;

always @(posedge a19886)
   l936 <= a19886;

always @(posedge a19494)
   l938 <= a19494;

always @(posedge a20898)
   l940 <= a20898;

always @(posedge na21812)
   l942 <= na21812;

always @(posedge a22630)
   l944 <= a22630;

always @(posedge na6674)
   l946 <= na6674;

always @(posedge z1)
   l948 <= z1;

always @(posedge a22638)
   l950 <= a22638;

always @(posedge a22656)
   l952 <= a22656;

always @(posedge a22664)
   l954 <= a22664;

always @(posedge a22668)
   l956 <= a22668;

always @(posedge a22670)
   l958 <= a22670;

always @(posedge a22676)
   l960 <= a22676;

always @(posedge l964)
   l962 <= l964;

always @(posedge z2)
   l964 <= z2;

always @(posedge l968)
   l966 <= l968;

always @(posedge na11396)
   l968 <= na11396;

always @(posedge z3)
   l970 <= z3;

always @(posedge z4)
   l972 <= z4;

always @(posedge z5)
   l974 <= z5;

always @(posedge z6)
   l976 <= z6;

always @(posedge a15296)
   l978 <= a15296;

always @(posedge a22688)
   l980 <= a22688;

always @(posedge a22696)
   l982 <= a22696;

always @(posedge a22706)
   l984 <= a22706;

always @(posedge a22712)
   l986 <= a22712;

always @(posedge a22686)
   l988 <= a22686;

always @(posedge a24442)
   l990 <= a24442;

always @(posedge a24660)
   l992 <= a24660;

always @(posedge a26604)
   l994 <= a26604;

always @(posedge a26614)
   l996 <= a26614;

always @(posedge a26616)
   l998 <= a26616;

always @(posedge a26622)
   l1000 <= a26622;

always @(posedge a10920)
   l1002 <= a10920;

always @(posedge a10962)
   l1004 <= a10962;

always @(posedge a10816)
   l1006 <= a10816;

always @(posedge a10876)
   l1008 <= a10876;

always @(posedge a27060)
   l1010 <= a27060;

always @(posedge a11278)
   l1012 <= a11278;

always @(posedge a22600)
   l1014 <= a22600;

always @(posedge a15956)
   l1016 <= a15956;

always @(posedge a22172)
   l1018 <= a22172;

always @(posedge a27108)
   l1020 <= a27108;

always @(posedge a15858)
   l1022 <= a15858;

always @(posedge a22230)
   l1024 <= a22230;

always @(posedge a27156)
   l1026 <= a27156;

always @(posedge a15760)
   l1028 <= a15760;

always @(posedge a22288)
   l1030 <= a22288;

always @(posedge a27204)
   l1032 <= a27204;

always @(posedge a15656)
   l1034 <= a15656;

always @(posedge a22346)
   l1036 <= a22346;

always @(posedge a27252)
   l1038 <= a27252;

always @(posedge a15552)
   l1040 <= a15552;

always @(posedge a22404)
   l1042 <= a22404;

always @(posedge a27300)
   l1044 <= a27300;

always @(posedge a15448)
   l1046 <= a15448;

always @(posedge a22462)
   l1048 <= a22462;

always @(posedge a27348)
   l1050 <= a27348;

always @(posedge a27382)
   l1052 <= a27382;

always @(posedge a11380)
   l1054 <= a11380;

always @(posedge a22520)
   l1056 <= a22520;

always @(posedge a27398)
   l1058 <= a27398;

always @(posedge a27414)
   l1060 <= a27414;

always @(posedge a27430)
   l1062 <= a27430;

always @(posedge a11040)
   l1064 <= a11040;

always @(posedge a27454)
   l1066 <= a27454;

always @(posedge a27460)
   l1068 <= a27460;

always @(posedge a27466)
   l1070 <= a27466;

always @(posedge a27472)
   l1072 <= a27472;

always @(posedge a27478)
   l1074 <= a27478;

always @(posedge a27484)
   l1076 <= a27484;

always @(posedge a27490)
   l1078 <= a27490;

always @(posedge a27498)
   l1080 <= a27498;

always @(posedge a28230)
   l1082 <= a28230;

always @(posedge a28254)
   l1084 <= a28254;

always @(posedge a28004)
   l1086 <= a28004;

always @(posedge a28082)
   l1088 <= a28082;

always @(posedge a28278)
   l1090 <= a28278;

always @(posedge a28302)
   l1092 <= a28302;

always @(posedge a27902)
   l1094 <= a27902;

always @(posedge a27890)
   l1096 <= a27890;

always @(posedge a27802)
   l1098 <= a27802;

always @(posedge a27790)
   l1100 <= a27790;

always @(posedge a27698)
   l1102 <= a27698;

always @(posedge a27684)
   l1104 <= a27684;

always @(posedge a27588)
   l1106 <= a27588;

always @(posedge a27572)
   l1108 <= a27572;

always @(posedge a28314)
   l1110 <= a28314;

always @(posedge a28320)
   l1112 <= a28320;

always @(posedge a28326)
   l1114 <= a28326;

always @(posedge a28332)
   l1116 <= a28332;

always @(posedge a28338)
   l1118 <= a28338;

always @(posedge a28344)
   l1120 <= a28344;

always @(posedge a28350)
   l1122 <= a28350;

always @(posedge a28356)
   l1124 <= a28356;

always @(posedge a28362)
   l1126 <= a28362;

always @(posedge a28368)
   l1128 <= a28368;

always @(posedge a24820)
   l1130 <= a24820;

always @(posedge a24812)
   l1132 <= a24812;

always @(posedge a24792)
   l1134 <= a24792;

always @(posedge a24784)
   l1136 <= a24784;

always @(posedge a24772)
   l1138 <= a24772;

always @(posedge a24764)
   l1140 <= a24764;

always @(posedge a24748)
   l1142 <= a24748;

always @(posedge a24740)
   l1144 <= a24740;

always @(posedge a24728)
   l1146 <= a24728;

always @(posedge a24720)
   l1148 <= a24720;

always @(posedge na26802)
   l1150 <= na26802;

always @(posedge a28380)
   l1152 <= a28380;

always @(posedge a28386)
   l1154 <= a28386;

always @(posedge a28392)
   l1156 <= a28392;

always @(posedge a28398)
   l1158 <= a28398;

always @(posedge a28404)
   l1160 <= a28404;

always @(posedge a28410)
   l1162 <= a28410;

always @(posedge a28416)
   l1164 <= a28416;

always @(posedge a28422)
   l1166 <= a28422;

always @(posedge a28428)
   l1168 <= a28428;

always @(posedge a28434)
   l1170 <= a28434;

always @(posedge a25690)
   l1172 <= a25690;

always @(posedge a25682)
   l1174 <= a25682;

always @(posedge a25662)
   l1176 <= a25662;

always @(posedge a25654)
   l1178 <= a25654;

always @(posedge a25642)
   l1180 <= a25642;

always @(posedge a25634)
   l1182 <= a25634;

always @(posedge a25618)
   l1184 <= a25618;

always @(posedge a25610)
   l1186 <= a25610;

always @(posedge a25598)
   l1188 <= a25598;

always @(posedge a25590)
   l1190 <= a25590;

always @(posedge na26780)
   l1192 <= na26780;

always @(posedge a28446)
   l1194 <= a28446;

always @(posedge a28452)
   l1196 <= a28452;

always @(posedge a28458)
   l1198 <= a28458;

always @(posedge a28464)
   l1200 <= a28464;

always @(posedge a28470)
   l1202 <= a28470;

always @(posedge a28476)
   l1204 <= a28476;

always @(posedge a28482)
   l1206 <= a28482;

always @(posedge a28488)
   l1208 <= a28488;

always @(posedge a28494)
   l1210 <= a28494;

always @(posedge a28500)
   l1212 <= a28500;

always @(posedge a25566)
   l1214 <= a25566;

always @(posedge a25558)
   l1216 <= a25558;

always @(posedge a25538)
   l1218 <= a25538;

always @(posedge a25530)
   l1220 <= a25530;

always @(posedge a25518)
   l1222 <= a25518;

always @(posedge a25510)
   l1224 <= a25510;

always @(posedge a25494)
   l1226 <= a25494;

always @(posedge a25486)
   l1228 <= a25486;

always @(posedge a25474)
   l1230 <= a25474;

always @(posedge a25466)
   l1232 <= a25466;

always @(posedge na26752)
   l1234 <= na26752;

always @(posedge a28512)
   l1236 <= a28512;

always @(posedge a28518)
   l1238 <= a28518;

always @(posedge a28524)
   l1240 <= a28524;

always @(posedge a28530)
   l1242 <= a28530;

always @(posedge a28536)
   l1244 <= a28536;

always @(posedge a28542)
   l1246 <= a28542;

always @(posedge a28548)
   l1248 <= a28548;

always @(posedge a28554)
   l1250 <= a28554;

always @(posedge a28560)
   l1252 <= a28560;

always @(posedge a28566)
   l1254 <= a28566;

always @(posedge a25442)
   l1256 <= a25442;

always @(posedge a25434)
   l1258 <= a25434;

always @(posedge a25414)
   l1260 <= a25414;

always @(posedge a25406)
   l1262 <= a25406;

always @(posedge a25394)
   l1264 <= a25394;

always @(posedge a25386)
   l1266 <= a25386;

always @(posedge a25370)
   l1268 <= a25370;

always @(posedge a25362)
   l1270 <= a25362;

always @(posedge a25350)
   l1272 <= a25350;

always @(posedge a25342)
   l1274 <= a25342;

always @(posedge na26724)
   l1276 <= na26724;

always @(posedge a28578)
   l1278 <= a28578;

always @(posedge a28584)
   l1280 <= a28584;

always @(posedge a28590)
   l1282 <= a28590;

always @(posedge a28596)
   l1284 <= a28596;

always @(posedge a28602)
   l1286 <= a28602;

always @(posedge a28608)
   l1288 <= a28608;

always @(posedge a28614)
   l1290 <= a28614;

always @(posedge a28620)
   l1292 <= a28620;

always @(posedge a28626)
   l1294 <= a28626;

always @(posedge a28632)
   l1296 <= a28632;

always @(posedge a25318)
   l1298 <= a25318;

always @(posedge a25310)
   l1300 <= a25310;

always @(posedge a25290)
   l1302 <= a25290;

always @(posedge a25282)
   l1304 <= a25282;

always @(posedge a25270)
   l1306 <= a25270;

always @(posedge a25262)
   l1308 <= a25262;

always @(posedge a25246)
   l1310 <= a25246;

always @(posedge a25238)
   l1312 <= a25238;

always @(posedge a25226)
   l1314 <= a25226;

always @(posedge a25218)
   l1316 <= a25218;

always @(posedge na26696)
   l1318 <= na26696;

always @(posedge a28644)
   l1320 <= a28644;

always @(posedge a28650)
   l1322 <= a28650;

always @(posedge a28656)
   l1324 <= a28656;

always @(posedge a28662)
   l1326 <= a28662;

always @(posedge a28668)
   l1328 <= a28668;

always @(posedge a28674)
   l1330 <= a28674;

always @(posedge a28680)
   l1332 <= a28680;

always @(posedge a28686)
   l1334 <= a28686;

always @(posedge a28692)
   l1336 <= a28692;

always @(posedge a28698)
   l1338 <= a28698;

always @(posedge a25194)
   l1340 <= a25194;

always @(posedge a25186)
   l1342 <= a25186;

always @(posedge a25166)
   l1344 <= a25166;

always @(posedge a25158)
   l1346 <= a25158;

always @(posedge a25146)
   l1348 <= a25146;

always @(posedge a25138)
   l1350 <= a25138;

always @(posedge a25122)
   l1352 <= a25122;

always @(posedge a25114)
   l1354 <= a25114;

always @(posedge a25102)
   l1356 <= a25102;

always @(posedge a25094)
   l1358 <= a25094;

always @(posedge na26668)
   l1360 <= na26668;

always @(posedge a28710)
   l1362 <= a28710;

always @(posedge a28716)
   l1364 <= a28716;

always @(posedge a28722)
   l1366 <= a28722;

always @(posedge a28728)
   l1368 <= a28728;

always @(posedge a28734)
   l1370 <= a28734;

always @(posedge a28740)
   l1372 <= a28740;

always @(posedge a28746)
   l1374 <= a28746;

always @(posedge a28752)
   l1376 <= a28752;

always @(posedge a28758)
   l1378 <= a28758;

always @(posedge a28764)
   l1380 <= a28764;

always @(posedge a25070)
   l1382 <= a25070;

always @(posedge a25062)
   l1384 <= a25062;

always @(posedge a25042)
   l1386 <= a25042;

always @(posedge a25034)
   l1388 <= a25034;

always @(posedge a25022)
   l1390 <= a25022;

always @(posedge a25014)
   l1392 <= a25014;

always @(posedge a24998)
   l1394 <= a24998;

always @(posedge a24990)
   l1396 <= a24990;

always @(posedge a24978)
   l1398 <= a24978;

always @(posedge a24970)
   l1400 <= a24970;

always @(posedge a26636)
   l1402 <= a26636;

always @(posedge a28776)
   l1404 <= a28776;

always @(posedge a28782)
   l1406 <= a28782;

always @(posedge a28788)
   l1408 <= a28788;

always @(posedge a28794)
   l1410 <= a28794;

always @(posedge a28800)
   l1412 <= a28800;

always @(posedge a28806)
   l1414 <= a28806;

always @(posedge a28812)
   l1416 <= a28812;

always @(posedge a28818)
   l1418 <= a28818;

always @(posedge a28824)
   l1420 <= a28824;

always @(posedge a28830)
   l1422 <= a28830;

always @(posedge a24946)
   l1424 <= a24946;

always @(posedge a24938)
   l1426 <= a24938;

always @(posedge a24918)
   l1428 <= a24918;

always @(posedge a24910)
   l1430 <= a24910;

always @(posedge a24898)
   l1432 <= a24898;

always @(posedge a24890)
   l1434 <= a24890;

always @(posedge a24874)
   l1436 <= a24874;

always @(posedge a24866)
   l1438 <= a24866;

always @(posedge a24854)
   l1440 <= a24854;

always @(posedge a24846)
   l1442 <= a24846;

always @(posedge a22946)
   l1444 <= a22946;

always @(posedge a22778)
   l1446 <= a22778;

always @(posedge a22806)
   l1448 <= a22806;

always @(posedge a22834)
   l1450 <= a22834;

always @(posedge a22862)
   l1452 <= a22862;

always @(posedge a22890)
   l1454 <= a22890;

always @(posedge a22918)
   l1456 <= a22918;

always @(posedge a22750)
   l1458 <= a22750;

always @(posedge a28834)
   l1460 <= a28834;

always @(posedge na28842)
   l1462 <= na28842;

always @(posedge na28854)
   l1464 <= na28854;

always @(posedge a28866)
   l1466 <= a28866;

always @(posedge a28878)
   l1468 <= a28878;

always @(posedge z7)
   l1470 <= z7;

always @(posedge a28882)
   l1472 <= a28882;

always @(posedge a28888)
   l1474 <= a28888;

always @(posedge a28894)
   l1476 <= a28894;

always @(posedge a28900)
   l1478 <= a28900;

always @(posedge a28906)
   l1480 <= a28906;

always @(posedge a28912)
   l1482 <= a28912;

always @(posedge a28918)
   l1484 <= a28918;

always @(posedge a28924)
   l1486 <= a28924;

always @(posedge a21698)
   l1488 <= a21698;

always @(posedge na24508)
   l1490 <= na24508;

always @(posedge na1690)
   l1492 <= na1690;

always @(posedge l1496)
   l1494 <= l1496;

always @(posedge z8)
   l1496 <= z8;

always @(posedge a28938)
   l1498 <= a28938;

always @(posedge a28942)
   l1500 <= a28942;

always @(posedge a28972)
   l1502 <= a28972;

always @(posedge a17616)
   l1504 <= a17616;

always @(posedge a29058)
   l1506 <= a29058;

always @(posedge a29072)
   l1508 <= a29072;

always @(posedge a29084)
   l1510 <= a29084;

always @(posedge a29096)
   l1512 <= a29096;

always @(posedge a17748)
   l1514 <= a17748;

always @(posedge a17488)
   l1516 <= a17488;

always @(posedge a17350)
   l1518 <= a17350;

always @(posedge a17216)
   l1520 <= a17216;

always @(posedge a17082)
   l1522 <= a17082;

always @(posedge a16950)
   l1524 <= a16950;

always @(posedge a16808)
   l1526 <= a16808;

always @(posedge a16674)
   l1528 <= a16674;

always @(posedge a16356)
   l1530 <= a16356;

always @(posedge a29102)
   l1532 <= a29102;

always @(posedge a29108)
   l1534 <= a29108;

always @(posedge a29114)
   l1536 <= a29114;

always @(posedge a29120)
   l1538 <= a29120;

always @(posedge a28072)
   l1540 <= a28072;

always @(posedge a29122)
   l1542 <= a29122;

always @(posedge a27972)
   l1544 <= a27972;

always @(posedge a27938)
   l1546 <= a27938;

always @(posedge a27872)
   l1548 <= a27872;

always @(posedge a27838)
   l1550 <= a27838;

always @(posedge a27768)
   l1552 <= a27768;

always @(posedge a27734)
   l1554 <= a27734;

always @(posedge a27664)
   l1556 <= a27664;

always @(posedge a27630)
   l1558 <= a27630;

always @(posedge a29132)
   l1560 <= a29132;

always @(posedge a27452)
   l1562 <= a27452;

always @(posedge na27436)
   l1564 <= na27436;

always @(posedge a29144)
   l1566 <= a29144;

always @(posedge a29154)
   l1568 <= a29154;

always @(posedge a29160)
   l1570 <= a29160;

always @(posedge a19484)
   l1572 <= a19484;

always @(posedge a19474)
   l1574 <= a19474;

always @(posedge a19510)
   l1576 <= a19510;

always @(posedge a19518)
   l1578 <= a19518;

always @(posedge a19526)
   l1580 <= a19526;

always @(posedge a19534)
   l1582 <= a19534;

always @(posedge a29170)
   l1584 <= a29170;

always @(posedge a29180)
   l1586 <= a29180;

always @(posedge a29190)
   l1588 <= a29190;

always @(posedge a29200)
   l1590 <= a29200;

always @(posedge a29210)
   l1592 <= a29210;

always @(posedge a29220)
   l1594 <= a29220;

always @(posedge a29230)
   l1596 <= a29230;

always @(posedge a29240)
   l1598 <= a29240;

always @(posedge na29242)
   l1600 <= na29242;

always @(posedge a29340)
   l1602 <= a29340;

always @(posedge z9)
   l1604 <= z9;

always @(posedge a29390)
   l1606 <= a29390;

always @(posedge a29408)
   l1608 <= a29408;

always @(posedge a29426)
   l1610 <= a29426;

always @(posedge a29440)
   l1612 <= a29440;

always @(posedge a30318)
   l1614 <= a30318;

always @(posedge a30352)
   l1616 <= a30352;

always @(posedge na30354)
   l1618 <= na30354;

always @(posedge na30356)
   l1620 <= na30356;

always @(posedge na30358)
   l1622 <= na30358;

always @(posedge a30366)
   l1624 <= a30366;

always @(posedge na2330)
   l1626 <= na2330;

always @(posedge na2332)
   l1628 <= na2332;

always @(posedge na2336)
   l1630 <= na2336;

always @(posedge a30384)
   l1632 <= a30384;

always @(posedge na30386)
   l1634 <= na30386;

always @(posedge a30392)
   l1636 <= a30392;

always @(posedge na2334)
   l1638 <= na2334;

always @(posedge a30410)
   l1640 <= a30410;

always @(posedge a30416)
   l1642 <= a30416;

always @(posedge a30428)
   l1644 <= a30428;

always @(posedge a30434)
   l1646 <= a30434;

always @(posedge a30468)
   l1648 <= a30468;

always @(posedge a30482)
   l1650 <= a30482;

always @(posedge a30490)
   l1652 <= a30490;

always @(posedge a30496)
   l1654 <= a30496;

always @(posedge a30506)
   l1656 <= a30506;

always @(posedge a32028)
   l1658 <= a32028;

always @(posedge a32548)
   l1660 <= a32548;

always @(posedge na32550)
   l1662 <= na32550;

always @(posedge a29254)
   l1664 <= a29254;

always @(posedge na32552)
   l1666 <= na32552;

always @(posedge a29248)
   l1668 <= a29248;

always @(posedge na32554)
   l1670 <= na32554;

always @(posedge a29262)
   l1672 <= a29262;

always @(posedge na32556)
   l1674 <= na32556;

always @(posedge a29270)
   l1676 <= a29270;

always @(posedge l1680)
   l1678 <= l1680;

always @(posedge na32562)
   l1680 <= na32562;

always @(posedge na15294)
   l1682 <= na15294;

always @(posedge a32564)
   l1684 <= a32564;

always @(posedge c1)
   l1686 <= c1;


assign a6662 = ~a6660 & a6658;
assign a6682 = a6680 & ~a6674;
assign a6690 = ~a6688 & ~a6684;
assign a6696 = ~a6694 & ~a6692;
assign a6702 = ~a6700 & ~a6698;
assign a6708 = ~a6706 & ~a6704;
assign na6710 = ~a6710;
assign a6712 = a6338 & ~a6336;
assign a6074 = ~a6072 & i4;
assign a6920 = ~a6918 & ~a6910;
assign a7152 = ~a7150 & ~a7148;
assign a7352 = ~a7350 & ~a7348;
assign a7590 = ~a7588 & ~a7586;
assign a7812 = ~a7810 & ~a7808;
assign a7852 = ~a7850 & ~a7848;
assign a7864 = ~a7862 & ~a7854;
assign a7900 = ~a7898 & ~a7896;
assign a7930 = ~a7928 & ~a7926;
assign a7942 = ~a7940 & ~a7932;
assign a7954 = ~a7952 & ~a7944;
assign a7966 = ~a7964 & ~a7956;
assign a7978 = ~a7976 & ~a7968;
assign a7990 = ~a7988 & ~a7980;
assign a8002 = ~a8000 & ~a7992;
assign a8020 = ~a8018 & ~a8016;
assign a16268 = ~a16266 & ~a16264;
assign a16274 = ~a16272 & ~a16270;
assign a16280 = ~a16278 & ~a16276;
assign a16286 = ~a16284 & ~a16282;
assign a16292 = ~a16290 & ~a16288;
assign a16298 = ~a16296 & ~a16294;
assign a16304 = ~a16302 & ~a16300;
assign a16310 = ~a16308 & ~a16306;
assign a16660 = ~a16658 & a16466;
assign a16800 = ~a16798 & a16780;
assign a16936 = ~a16934 & a16914;
assign a17072 = ~a17070 & a17056;
assign a17208 = ~a17206 & a17188;
assign a17342 = ~a17340 & a17322;
assign a17476 = ~a17474 & a17456;
assign a17610 = ~a17608 & a17594;
assign a17742 = ~a17740 & a17724;
assign a17872 = ~a17870 & a17854;
assign a15370 = ~a15368 & ~a15366;
assign a15474 = ~a15472 & ~a15470;
assign a15578 = ~a15576 & ~a15574;
assign a15682 = ~a15680 & ~a15678;
assign a15786 = ~a15784 & ~a15782;
assign a15884 = ~a15882 & ~a15880;
assign a15982 = ~a15980 & ~a15978;
assign na2430 = ~a2430;
assign a17882 = ~a17880 & a17878;
assign na2432 = ~a2432;
assign na2436 = ~a2436;
assign a17900 = ~a17898 & a17896;
assign a17916 = ~a17914 & a17912;
assign na2434 = ~a2434;
assign na5594 = ~a5594;
assign na5596 = ~a5596;
assign na5600 = ~a5600;
assign na5598 = ~a5598;
assign a6592 = ~a6590 & ~a6584;
assign a6476 = ~a6474 & ~a6464;
assign a6548 = ~a6546 & ~a6538;
assign a6512 = ~a6510 & ~a6508;
assign na17918 = ~a17918;
assign na17920 = ~a17920;
assign na17922 = ~a17922;
assign na17924 = ~a17924;
assign a15314 = ~a15312 & ~a15310;
assign a6522 = ~a6520 & ~a6518;
assign a6566 = ~a6564 & ~a6554;
assign a6608 = ~a6606 & ~a6598;
assign a6494 = ~a6492 & ~a6482;
assign a18026 = a18024 & a17974;
assign na18028 = ~a18028;
assign na6410 = ~a6410;
assign na6404 = ~a6404;
assign a6424 = ~a6422 & ~a6348;
assign a6448 = ~a6446 & ~a6430;
assign a18098 = ~a18096 & a18034;
assign z0 = l494;
assign a19208 = ~a19206 & a19178;
assign a19248 = ~a19246 & ~a19244;
assign a19262 = ~a19260 & ~a19258;
assign a19274 = ~a19272 & ~a19270;
assign a19282 = ~a19280 & ~a19278;
assign a19292 = ~a19290 & ~a19288;
assign a19300 = ~a19298 & ~a19296;
assign a19308 = ~a19306 & ~a19304;
assign a19318 = ~a19316 & ~a19314;
assign a19326 = ~a19324 & ~a19322;
assign a19334 = ~a19332 & ~a19330;
assign a19342 = ~a19340 & ~a19338;
assign a19348 = ~a19346 & ~a19344;
assign a19354 = ~a19352 & ~a19350;
assign a19360 = ~a19358 & ~a19356;
assign a19336 = a11112 & a6934;
assign na16352 = ~a16352;
assign na19362 = ~a19362;
assign a6346 = a6344 & ~a2262;
assign a19364 = a11186 & i480;
assign a19924 = ~a19922 & ~a19920;
assign a19912 = ~a19910 & ~a19898;
assign a19834 = ~a19832 & ~a19830;
assign a19808 = ~a19806 & ~a19800;
assign a19770 = ~a19768 & ~a19762;
assign a19732 = ~a19730 & ~a19724;
assign a19698 = ~a19696 & ~a19690;
assign a19664 = ~a19662 & ~a19656;
assign a19630 = ~a19628 & ~a19546;
assign a19926 = ~a16052 & ~a6682;
assign a19938 = ~a19936 & ~a19934;
assign a19944 = ~a19942 & ~a19940;
assign a19950 = ~a19948 & ~a19946;
assign a19956 = ~a19954 & ~a19952;
assign a19962 = ~a19960 & ~a19958;
assign a19968 = ~a19966 & ~a19964;
assign a19974 = ~a19972 & ~a19970;
assign a19980 = ~a19978 & ~a19976;
assign a19986 = ~a19984 & ~a19982;
assign a19992 = ~a19990 & ~a19988;
assign a16070 = ~a16068 & ~a7952;
assign a20004 = ~a20002 & ~a20000;
assign a20010 = ~a20008 & ~a20006;
assign a20016 = ~a20014 & ~a20012;
assign a20022 = ~a20020 & ~a20018;
assign a20028 = ~a20026 & ~a20024;
assign a20034 = ~a20032 & ~a20030;
assign a20040 = ~a20038 & ~a20036;
assign a20046 = ~a20044 & ~a20042;
assign a20052 = ~a20050 & ~a20048;
assign a20058 = ~a20056 & ~a20054;
assign a20060 = ~a16080 & ~a6682;
assign a20072 = ~a20070 & ~a20068;
assign a20078 = ~a20076 & ~a20074;
assign a20084 = ~a20082 & ~a20080;
assign a20090 = ~a20088 & ~a20086;
assign a20096 = ~a20094 & ~a20092;
assign a20102 = ~a20100 & ~a20098;
assign a20108 = ~a20106 & ~a20104;
assign a20114 = ~a20112 & ~a20110;
assign a20120 = ~a20118 & ~a20116;
assign a20126 = ~a20124 & ~a20122;
assign a20128 = ~a16090 & ~a6682;
assign a20140 = ~a20138 & ~a20136;
assign a20146 = ~a20144 & ~a20142;
assign a20152 = ~a20150 & ~a20148;
assign a20158 = ~a20156 & ~a20154;
assign a20164 = ~a20162 & ~a20160;
assign a20170 = ~a20168 & ~a20166;
assign a20176 = ~a20174 & ~a20172;
assign a20182 = ~a20180 & ~a20178;
assign a20188 = ~a20186 & ~a20184;
assign a20194 = ~a20192 & ~a20190;
assign a20196 = ~a16100 & ~a6682;
assign a20208 = ~a20206 & ~a20204;
assign a20214 = ~a20212 & ~a20210;
assign a20220 = ~a20218 & ~a20216;
assign a20226 = ~a20224 & ~a20222;
assign a20232 = ~a20230 & ~a20228;
assign a20238 = ~a20236 & ~a20234;
assign a20244 = ~a20242 & ~a20240;
assign a20250 = ~a20248 & ~a20246;
assign a20256 = ~a20254 & ~a20252;
assign a20262 = ~a20260 & ~a20258;
assign a20264 = ~a16110 & ~a6682;
assign a20276 = ~a20274 & ~a20272;
assign a20282 = ~a20280 & ~a20278;
assign a20288 = ~a20286 & ~a20284;
assign a20294 = ~a20292 & ~a20290;
assign a20300 = ~a20298 & ~a20296;
assign a20306 = ~a20304 & ~a20302;
assign a20312 = ~a20310 & ~a20308;
assign a20318 = ~a20316 & ~a20314;
assign a20324 = ~a20322 & ~a20320;
assign a20330 = ~a20328 & ~a20326;
assign a20332 = ~a16120 & ~a6682;
assign a20344 = ~a20342 & ~a20340;
assign a20350 = ~a20348 & ~a20346;
assign a20356 = ~a20354 & ~a20352;
assign a20362 = ~a20360 & ~a20358;
assign a20368 = ~a20366 & ~a20364;
assign a20374 = ~a20372 & ~a20370;
assign a20380 = ~a20378 & ~a20376;
assign a20386 = ~a20384 & ~a20382;
assign a20392 = ~a20390 & ~a20388;
assign a20398 = ~a20396 & ~a20394;
assign a8042 = ~a8040 & ~a7862;
assign a20412 = ~a20410 & ~a20408;
assign a20418 = ~a20416 & ~a20414;
assign a20424 = ~a20422 & ~a20420;
assign a20430 = ~a20428 & ~a20426;
assign a20436 = ~a20434 & ~a20432;
assign a20442 = ~a20440 & ~a20438;
assign a20448 = ~a20446 & ~a20444;
assign a20454 = ~a20452 & ~a20450;
assign a20460 = ~a20458 & ~a20456;
assign a20466 = ~a20464 & ~a20462;
assign a20564 = ~a20562 & a20474;
assign a20636 = ~a20634 & a20574;
assign a20666 = ~a20664 & a20644;
assign a20716 = ~a20714 & a20678;
assign a20762 = ~a20760 & a20724;
assign a20800 = ~a20798 & a20770;
assign a20816 = ~a20814 & a20808;
assign a20836 = ~a20834 & a20822;
assign a20854 = ~a20852 & a20846;
assign a20870 = ~a20868 & a20862;
assign na20872 = ~a20872;
assign na20874 = ~a20874;
assign na20876 = ~a20876;
assign na20878 = ~a20878;
assign a6384 = ~a6382 & a6380;
assign a6372 = ~a6370 & a6368;
assign a6362 = ~a6360 & a6356;
assign a6394 = ~a6392 & a6390;
assign a19886 = ~a19884 & ~a19882;
assign a19494 = ~a19492 & ~a19490;
assign a20898 = a20896 & a15298;
assign na21812 = ~a21812;
assign a22630 = a22628 & a13494;
assign na6674 = ~a6674;
assign z1 = l946;
assign a22638 = ~a22636 & ~a22632;
assign a22656 = ~a22654 & ~a22646;
assign a22664 = ~a22662 & ~a15338;
assign a22668 = ~a22666 & ~a22654;
assign a22670 = ~a15336 & ~l958;
assign a22676 = ~a22674 & ~a22672;
assign z2 = l508;
assign na11396 = ~a11396;
assign z3 = l962;
assign z4 = l970;
assign z5 = l972;
assign z6 = l974;
assign a15296 = ~a15294 & a11420;
assign a22688 = ~a22686 & ~a22684;
assign a22696 = ~a22694 & ~a22686;
assign a22706 = a22704 & ~a22686;
assign a22712 = ~a22710 & ~a22686;
assign a22686 = a22636 & i416;
assign a24442 = ~a24440 & a22714;
assign a24660 = ~a24658 & ~a24656;
assign a26604 = ~a26602 & ~a26550;
assign a26614 = ~a26612 & ~a26610;
assign a26616 = ~a22624 & ~a8048;
assign a26622 = ~a26620 & ~a26618;
assign a10920 = ~a10918 & ~a6520;
assign a10962 = ~a10960 & ~a6564;
assign a10816 = ~a10814 & ~a6606;
assign a10876 = ~a10874 & ~a6492;
assign a27060 = ~a27058 & ~a6492;
assign a11278 = ~a11276 & a11218;
assign a22600 = ~a22598 & ~a22590;
assign a15956 = ~a15954 & a15910;
assign a22172 = ~a22170 & ~a22160;
assign a27108 = ~a27106 & ~a27104;
assign a15858 = ~a15856 & a15812;
assign a22230 = ~a22228 & ~a22220;
assign a27156 = ~a27154 & ~a27152;
assign a15760 = ~a15758 & a15714;
assign a22288 = ~a22286 & ~a22278;
assign a27204 = ~a27202 & ~a27200;
assign a15656 = ~a15654 & a15610;
assign a22346 = ~a22344 & ~a22336;
assign a27252 = ~a27250 & ~a27248;
assign a15552 = ~a15550 & a15506;
assign a22404 = ~a22402 & ~a22394;
assign a27300 = ~a27298 & ~a27296;
assign a15448 = ~a15446 & a15402;
assign a22462 = ~a22460 & ~a22452;
assign a27348 = ~a27346 & ~a27344;
assign a27382 = ~a27380 & ~a27378;
assign a11380 = ~a11378 & a11308;
assign a22520 = ~a22518 & ~a22510;
assign a27398 = ~a27396 & ~a6606;
assign a27414 = ~a27412 & ~a6564;
assign a27430 = ~a27428 & ~a6520;
assign a11040 = ~a11038 & ~a10968;
assign a27454 = a27452 & a27446;
assign a27460 = ~a27458 & ~a27456;
assign a27466 = ~a27464 & ~a27462;
assign a27472 = ~a27470 & ~a27468;
assign a27478 = ~a27476 & ~a27474;
assign a27484 = ~a27482 & ~a27480;
assign a27490 = ~a27488 & ~a27486;
assign a27498 = a27496 & ~a27492;
assign a28230 = ~a28228 & ~a28224;
assign a28254 = ~a28252 & ~a28248;
assign a28004 = a28002 & l584;
assign a28082 = a28080 & a17872;
assign a28278 = ~a28276 & ~a28272;
assign a28302 = ~a28300 & ~a28296;
assign a27902 = a27900 & a17610;
assign a27890 = a27888 & a17476;
assign a27802 = a27800 & a17342;
assign a27790 = a27788 & a17208;
assign a27698 = a27696 & a17072;
assign a27684 = a27682 & a16936;
assign a27588 = a27586 & a16800;
assign a27572 = a27570 & a16660;
assign a28314 = ~a28312 & ~a28304;
assign a28320 = ~a28318 & ~a28316;
assign a28326 = ~a28324 & ~a28322;
assign a28332 = ~a28330 & ~a28328;
assign a28338 = ~a28336 & ~a28334;
assign a28344 = ~a28342 & ~a28340;
assign a28350 = ~a28348 & ~a28346;
assign a28356 = ~a28354 & ~a28352;
assign a28362 = ~a28360 & ~a28358;
assign a28368 = ~a28366 & ~a28364;
assign a24820 = ~a24818 & ~a24816;
assign a24812 = ~a24810 & ~a24808;
assign a24792 = ~a24790 & ~a24788;
assign a24784 = ~a24782 & ~a24780;
assign a24772 = ~a24770 & ~a24768;
assign a24764 = ~a24762 & ~a24760;
assign a24748 = ~a24746 & ~a24744;
assign a24740 = ~a24738 & ~a24736;
assign a24728 = ~a24726 & ~a24724;
assign a24720 = ~a24718 & ~a24716;
assign na26802 = ~a26802;
assign a28380 = ~a28378 & ~a28370;
assign a28386 = ~a28384 & ~a28382;
assign a28392 = ~a28390 & ~a28388;
assign a28398 = ~a28396 & ~a28394;
assign a28404 = ~a28402 & ~a28400;
assign a28410 = ~a28408 & ~a28406;
assign a28416 = ~a28414 & ~a28412;
assign a28422 = ~a28420 & ~a28418;
assign a28428 = ~a28426 & ~a28424;
assign a28434 = ~a28432 & ~a28430;
assign a25690 = ~a25688 & ~a25686;
assign a25682 = ~a25680 & ~a25678;
assign a25662 = ~a25660 & ~a25658;
assign a25654 = ~a25652 & ~a25650;
assign a25642 = ~a25640 & ~a25638;
assign a25634 = ~a25632 & ~a25630;
assign a25618 = ~a25616 & ~a25614;
assign a25610 = ~a25608 & ~a25606;
assign a25598 = ~a25596 & ~a25594;
assign a25590 = ~a25588 & ~a25586;
assign na26780 = ~a26780;
assign a28446 = ~a28444 & ~a28436;
assign a28452 = ~a28450 & ~a28448;
assign a28458 = ~a28456 & ~a28454;
assign a28464 = ~a28462 & ~a28460;
assign a28470 = ~a28468 & ~a28466;
assign a28476 = ~a28474 & ~a28472;
assign a28482 = ~a28480 & ~a28478;
assign a28488 = ~a28486 & ~a28484;
assign a28494 = ~a28492 & ~a28490;
assign a28500 = ~a28498 & ~a28496;
assign a25566 = ~a25564 & ~a25562;
assign a25558 = ~a25556 & ~a25554;
assign a25538 = ~a25536 & ~a25534;
assign a25530 = ~a25528 & ~a25526;
assign a25518 = ~a25516 & ~a25514;
assign a25510 = ~a25508 & ~a25506;
assign a25494 = ~a25492 & ~a25490;
assign a25486 = ~a25484 & ~a25482;
assign a25474 = ~a25472 & ~a25470;
assign a25466 = ~a25464 & ~a25462;
assign na26752 = ~a26752;
assign a28512 = ~a28510 & ~a28502;
assign a28518 = ~a28516 & ~a28514;
assign a28524 = ~a28522 & ~a28520;
assign a28530 = ~a28528 & ~a28526;
assign a28536 = ~a28534 & ~a28532;
assign a28542 = ~a28540 & ~a28538;
assign a28548 = ~a28546 & ~a28544;
assign a28554 = ~a28552 & ~a28550;
assign a28560 = ~a28558 & ~a28556;
assign a28566 = ~a28564 & ~a28562;
assign a25442 = ~a25440 & ~a25438;
assign a25434 = ~a25432 & ~a25430;
assign a25414 = ~a25412 & ~a25410;
assign a25406 = ~a25404 & ~a25402;
assign a25394 = ~a25392 & ~a25390;
assign a25386 = ~a25384 & ~a25382;
assign a25370 = ~a25368 & ~a25366;
assign a25362 = ~a25360 & ~a25358;
assign a25350 = ~a25348 & ~a25346;
assign a25342 = ~a25340 & ~a25338;
assign na26724 = ~a26724;
assign a28578 = ~a28576 & ~a28568;
assign a28584 = ~a28582 & ~a28580;
assign a28590 = ~a28588 & ~a28586;
assign a28596 = ~a28594 & ~a28592;
assign a28602 = ~a28600 & ~a28598;
assign a28608 = ~a28606 & ~a28604;
assign a28614 = ~a28612 & ~a28610;
assign a28620 = ~a28618 & ~a28616;
assign a28626 = ~a28624 & ~a28622;
assign a28632 = ~a28630 & ~a28628;
assign a25318 = ~a25316 & ~a25314;
assign a25310 = ~a25308 & ~a25306;
assign a25290 = ~a25288 & ~a25286;
assign a25282 = ~a25280 & ~a25278;
assign a25270 = ~a25268 & ~a25266;
assign a25262 = ~a25260 & ~a25258;
assign a25246 = ~a25244 & ~a25242;
assign a25238 = ~a25236 & ~a25234;
assign a25226 = ~a25224 & ~a25222;
assign a25218 = ~a25216 & ~a25214;
assign na26696 = ~a26696;
assign a28644 = ~a28642 & ~a28634;
assign a28650 = ~a28648 & ~a28646;
assign a28656 = ~a28654 & ~a28652;
assign a28662 = ~a28660 & ~a28658;
assign a28668 = ~a28666 & ~a28664;
assign a28674 = ~a28672 & ~a28670;
assign a28680 = ~a28678 & ~a28676;
assign a28686 = ~a28684 & ~a28682;
assign a28692 = ~a28690 & ~a28688;
assign a28698 = ~a28696 & ~a28694;
assign a25194 = ~a25192 & ~a25190;
assign a25186 = ~a25184 & ~a25182;
assign a25166 = ~a25164 & ~a25162;
assign a25158 = ~a25156 & ~a25154;
assign a25146 = ~a25144 & ~a25142;
assign a25138 = ~a25136 & ~a25134;
assign a25122 = ~a25120 & ~a25118;
assign a25114 = ~a25112 & ~a25110;
assign a25102 = ~a25100 & ~a25098;
assign a25094 = ~a25092 & ~a25090;
assign na26668 = ~a26668;
assign a28710 = ~a28708 & ~a28700;
assign a28716 = ~a28714 & ~a28712;
assign a28722 = ~a28720 & ~a28718;
assign a28728 = ~a28726 & ~a28724;
assign a28734 = ~a28732 & ~a28730;
assign a28740 = ~a28738 & ~a28736;
assign a28746 = ~a28744 & ~a28742;
assign a28752 = ~a28750 & ~a28748;
assign a28758 = ~a28756 & ~a28754;
assign a28764 = ~a28762 & ~a28760;
assign a25070 = ~a25068 & ~a25066;
assign a25062 = ~a25060 & ~a25058;
assign a25042 = ~a25040 & ~a25038;
assign a25034 = ~a25032 & ~a25030;
assign a25022 = ~a25020 & ~a25018;
assign a25014 = ~a25012 & ~a25010;
assign a24998 = ~a24996 & ~a24994;
assign a24990 = ~a24988 & ~a24986;
assign a24978 = ~a24976 & ~a24974;
assign a24970 = ~a24968 & ~a24966;
assign a26636 = ~a26634 & ~a26628;
assign a28776 = ~a28774 & ~a28766;
assign a28782 = ~a28780 & ~a28778;
assign a28788 = ~a28786 & ~a28784;
assign a28794 = ~a28792 & ~a28790;
assign a28800 = ~a28798 & ~a28796;
assign a28806 = ~a28804 & ~a28802;
assign a28812 = ~a28810 & ~a28808;
assign a28818 = ~a28816 & ~a28814;
assign a28824 = ~a28822 & ~a28820;
assign a28830 = ~a28828 & ~a28826;
assign a24946 = ~a24944 & ~a24942;
assign a24938 = ~a24936 & ~a24934;
assign a24918 = ~a24916 & ~a24914;
assign a24910 = ~a24908 & ~a24906;
assign a24898 = ~a24896 & ~a24894;
assign a24890 = ~a24888 & ~a24886;
assign a24874 = ~a24872 & ~a24870;
assign a24866 = ~a24864 & ~a24862;
assign a24854 = ~a24852 & ~a24850;
assign a24846 = ~a24844 & ~a24842;
assign a22946 = ~a22944 & ~a22942;
assign a22778 = ~a22776 & ~a22774;
assign a22806 = ~a22804 & ~a22802;
assign a22834 = ~a22832 & ~a22830;
assign a22862 = ~a22860 & ~a22858;
assign a22890 = ~a22888 & ~a22886;
assign a22918 = ~a22916 & ~a22914;
assign a22750 = ~a22748 & ~a22746;
assign a28834 = ~a28832 & ~a13508;
assign na28842 = ~a28842;
assign na28854 = ~a28854;
assign a28866 = ~a28864 & ~a28860;
assign a28878 = ~a28876 & ~a28872;
assign z7 = l976;
assign a28882 = a28880 & ~a1690;
assign a28888 = ~a28886 & ~a28884;
assign a28894 = ~a28892 & ~a28890;
assign a28900 = ~a28898 & ~a28896;
assign a28906 = ~a28904 & ~a28902;
assign a28912 = ~a28910 & ~a28908;
assign a28918 = ~a28916 & ~a28914;
assign a28924 = ~a28922 & ~a28920;
assign a21698 = ~a21696 & ~a6682;
assign na24508 = ~a24508;
assign na1690 = ~a1690;
assign z8 = l988;
assign a28938 = ~a28936 & ~a28934;
assign a28942 = a28940 & a26966;
assign a28972 = a28970 & a28964;
assign a17616 = ~a17614 & ~a17612;
assign a29058 = ~a29056 & ~a29054;
assign a29072 = ~a29070 & ~a29068;
assign a29084 = ~a29082 & ~a29080;
assign a29096 = ~a29094 & ~a29092;
assign a17748 = ~a17746 & ~a17744;
assign a17488 = ~a17486 & ~a17484;
assign a17350 = ~a17348 & ~a17346;
assign a17216 = ~a17214 & ~a17212;
assign a17082 = ~a17080 & ~a17078;
assign a16950 = ~a16948 & ~a16946;
assign a16808 = ~a16806 & ~a16804;
assign a16674 = ~a16672 & ~a16670;
assign a16356 = ~a16354 & ~a16346;
assign a29102 = ~a29100 & ~a29098;
assign a29108 = ~a29106 & ~a29104;
assign a29114 = ~a29112 & ~a29110;
assign a29120 = ~a29118 & ~a29116;
assign a28072 = a28070 & l586;
assign a29122 = ~a28036 & l584;
assign a27972 = a27970 & l582;
assign a27938 = a27936 & l580;
assign a27872 = a27870 & l578;
assign a27838 = a27836 & l576;
assign a27768 = a27766 & ~a5572;
assign a27734 = a27732 & ~a5556;
assign a27664 = a27662 & ~a5548;
assign a27630 = a27628 & ~a5542;
assign a29132 = a29130 & ~a19362;
assign a27452 = a27450 & ~l962;
assign na27436 = ~a27436;
assign a29144 = a29142 & ~a29140;
assign a29154 = ~a29152 & a20890;
assign a29160 = a29158 & ~l946;
assign a19484 = ~a19482 & ~a19480;
assign a19474 = ~a19472 & ~a19470;
assign a19510 = ~a19508 & ~a19506;
assign a19518 = ~a19516 & ~a19514;
assign a19526 = ~a19524 & ~a19522;
assign a19534 = ~a19532 & ~a19530;
assign a29170 = ~a29168 & ~a7996;
assign a29180 = ~a29178 & ~a6914;
assign a29190 = ~a29188 & ~a7984;
assign a29200 = ~a29198 & ~a7972;
assign a29210 = ~a29208 & ~a7960;
assign a29220 = ~a29218 & ~a7948;
assign a29230 = ~a29228 & ~a7936;
assign a29240 = ~a29238 & ~a7858;
assign na29242 = ~a29242;
assign a29340 = a29338 & a29316;
assign z9 = l664;
assign a29390 = ~a29388 & a29382;
assign a29408 = ~a29406 & a29404;
assign a29426 = ~a29424 & a29422;
assign a29440 = ~a29438 & a29436;
assign a30318 = a30316 & a22624;
assign a30352 = ~a30350 & a30342;
assign na30354 = ~a30354;
assign na30356 = ~a30356;
assign na30358 = ~a30358;
assign a30366 = ~a30364 & ~a30362;
assign na2330 = ~a2330;
assign na2332 = ~a2332;
assign na2336 = ~a2336;
assign a30384 = ~a30382 & a30380;
assign na30386 = ~a30386;
assign a30392 = ~a30390 & ~a30388;
assign na2334 = ~a2334;
assign a30410 = ~a30408 & a30406;
assign a30416 = ~a30414 & ~a30412;
assign a30428 = ~a30426 & a30424;
assign a30434 = ~a30432 & ~a30430;
assign a30468 = ~a30466 & ~l664;
assign a30482 = ~a30480 & ~a30472;
assign a30490 = ~a30488 & ~a30484;
assign a30496 = ~a30494 & ~a30492;
assign a30506 = ~a30504 & ~a30498;
assign a32028 = ~a32026 & a30674;
assign a32548 = ~a32546 & a32518;
assign na32550 = ~a32550;
assign a29254 = ~a29252 & ~a29250;
assign na32552 = ~a32552;
assign a29248 = ~a29246 & ~a29244;
assign na32554 = ~a32554;
assign a29262 = ~a29260 & ~a29258;
assign na32556 = ~a32556;
assign a29270 = ~a29268 & ~a29266;
assign na32562 = ~a32562;
assign na15294 = ~a15294;
assign a32564 = a6330 & l516;
assign c1 = 1;
assign a1688 = l1686 & ~l662;
assign a1690 = l1686 & ~l504;
assign a1692 = l1686 & ~l660;
assign a1694 = l1686 & ~l648;
assign a1696 = ~i16 & ~i14;
assign a1698 = a1696 & ~i10;
assign a1700 = ~a1696 & i10;
assign a1702 = ~a1700 & ~i8;
assign a1704 = ~a1702 & ~a1698;
assign a1706 = a1696 & i10;
assign a1708 = ~a1696 & ~i10;
assign a1710 = ~a1708 & ~a1706;
assign a1712 = ~a1710 & ~i8;
assign a1714 = a1710 & i8;
assign a1716 = ~a1714 & ~a1712;
assign a1718 = ~a1716 & i62;
assign a1720 = a1718 & a1704;
assign a1722 = ~a1720 & ~l1686;
assign a1724 = l1686 & l646;
assign a1726 = ~a1724 & ~a1722;
assign a1728 = a1716 & ~i62;
assign a1730 = ~a1728 & ~a1718;
assign a1732 = ~a1730 & ~l1686;
assign a1734 = l1686 & l642;
assign a1736 = ~a1734 & ~a1732;
assign a1738 = ~a1718 & ~a1704;
assign a1740 = ~a1738 & ~a1720;
assign a1742 = ~a1740 & ~l1686;
assign a1744 = l1686 & l644;
assign a1746 = ~a1744 & ~a1742;
assign a1748 = a1746 & a1736;
assign a1750 = a1748 & a1726;
assign a1752 = a1750 & a1694;
assign a1754 = ~a1746 & a1736;
assign a1756 = a1754 & a1694;
assign a1758 = a1756 & ~a1726;
assign a1760 = ~a1758 & ~a1752;
assign a1762 = ~a1706 & ~i20;
assign a1764 = i22 & i10;
assign a1766 = ~i24 & i14;
assign a1768 = ~a1766 & ~a1696;
assign a1770 = a1768 & a1764;
assign a1772 = a1770 & ~a1762;
assign a1774 = ~a1762 & i10;
assign a1776 = a1766 & i22;
assign a1778 = a1776 & a1774;
assign a1780 = a1700 & ~i22;
assign a1782 = a1780 & a1762;
assign a1784 = ~a1782 & ~a1778;
assign a1786 = a1784 & ~a1772;
assign a1788 = a1786 & ~i18;
assign a1790 = a1788 & ~a1696;
assign a1792 = a1790 & i12;
assign a1794 = ~a1790 & ~i12;
assign a1796 = ~a1794 & ~a1792;
assign a1798 = ~a1796 & i10;
assign a1800 = a1788 & a1708;
assign a1802 = ~a1800 & ~a1798;
assign a1804 = ~a1802 & i26;
assign a1806 = a1802 & ~i26;
assign a1808 = ~a1806 & ~a1804;
assign a1810 = ~a1808 & i8;
assign a1812 = ~a1802 & ~i8;
assign a1814 = ~a1812 & ~a1810;
assign a1816 = ~a1814 & i28;
assign a1818 = a1764 & a1762;
assign a1820 = a1774 & ~i22;
assign a1822 = ~a1820 & ~a1818;
assign a1824 = ~a1822 & a1766;
assign a1826 = i16 & ~i14;
assign a1828 = a1826 & a1818;
assign a1830 = ~a1828 & ~a1824;
assign a1832 = i24 & i14;
assign a1834 = a1832 & a1818;
assign a1836 = a1820 & a1768;
assign a1838 = ~a1836 & ~a1834;
assign a1840 = a1838 & a1830;
assign a1842 = ~a1840 & a1788;
assign a1844 = ~a1706 & ~i30;
assign a1846 = a1844 & a1842;
assign a1848 = ~a1700 & i32;
assign a1850 = ~a1848 & a1786;
assign a1852 = a1850 & ~a1846;
assign a1854 = ~a1852 & ~a1788;
assign a1856 = a1852 & ~i18;
assign a1858 = ~a1856 & ~a1854;
assign a1860 = a1858 & ~a1696;
assign a1862 = ~a1860 & ~i34;
assign a1864 = a1860 & i34;
assign a1866 = ~a1864 & ~a1792;
assign a1868 = a1866 & ~a1862;
assign a1870 = ~a1864 & ~a1862;
assign a1872 = ~a1870 & a1792;
assign a1874 = ~a1872 & ~a1868;
assign a1876 = a1874 & ~a1796;
assign a1878 = ~a1874 & a1796;
assign a1880 = ~a1878 & i10;
assign a1882 = a1880 & ~a1876;
assign a1884 = a1858 & a1708;
assign a1886 = ~a1884 & ~a1882;
assign a1888 = a1886 & ~i36;
assign a1890 = ~a1886 & i36;
assign a1892 = ~a1890 & ~a1804;
assign a1894 = a1892 & ~a1888;
assign a1896 = ~a1890 & ~a1888;
assign a1898 = ~a1896 & a1804;
assign a1900 = ~a1898 & ~a1894;
assign a1902 = a1900 & ~a1808;
assign a1904 = ~a1900 & a1808;
assign a1906 = ~a1904 & i8;
assign a1908 = a1906 & ~a1902;
assign a1910 = ~a1886 & ~i8;
assign a1912 = ~a1910 & ~a1908;
assign a1914 = a1912 & ~i38;
assign a1916 = ~a1912 & i38;
assign a1918 = ~a1916 & ~a1914;
assign a1920 = a1918 & ~a1816;
assign a1922 = ~a1918 & a1816;
assign a1924 = ~a1922 & ~a1920;
assign a1926 = a1814 & ~i28;
assign a1928 = ~a1926 & ~a1816;
assign a1930 = a1928 & ~a1924;
assign a1932 = ~a1916 & ~a1816;
assign a1934 = ~a1932 & ~a1914;
assign a1936 = ~a1892 & ~a1888;
assign a1938 = ~a1866 & ~a1862;
assign a1940 = a1854 & i22;
assign a1942 = ~a1854 & ~i22;
assign a1944 = ~a1942 & ~a1940;
assign a1946 = a1944 & ~a1696;
assign a1948 = ~a1946 & ~i40;
assign a1950 = a1946 & i40;
assign a1952 = ~a1950 & ~a1948;
assign a1954 = a1952 & ~a1938;
assign a1956 = ~a1952 & a1938;
assign a1958 = ~a1956 & ~a1954;
assign a1960 = ~a1958 & a1878;
assign a1962 = a1958 & ~a1878;
assign a1964 = ~a1962 & i10;
assign a1966 = a1964 & ~a1960;
assign a1968 = a1944 & a1708;
assign a1970 = ~a1968 & ~a1966;
assign a1972 = a1970 & ~i42;
assign a1974 = ~a1970 & i42;
assign a1976 = ~a1974 & ~a1972;
assign a1978 = a1976 & ~a1936;
assign a1980 = ~a1976 & a1936;
assign a1982 = ~a1980 & ~a1978;
assign a1984 = ~a1982 & a1904;
assign a1986 = a1982 & ~a1904;
assign a1988 = ~a1986 & i8;
assign a1990 = a1988 & ~a1984;
assign a1992 = ~a1970 & ~i8;
assign a1994 = ~a1992 & ~a1990;
assign a1996 = a1994 & ~i44;
assign a1998 = ~a1994 & i44;
assign a2000 = ~a1998 & ~a1996;
assign a2002 = a2000 & ~a1934;
assign a2004 = ~a2000 & a1934;
assign a2006 = ~a2004 & ~a2002;
assign a2008 = ~a2006 & a1930;
assign a2010 = ~a1998 & ~a1934;
assign a2012 = ~a2010 & ~a1996;
assign a2014 = ~a1974 & ~a1936;
assign a2016 = ~a2014 & ~a1972;
assign a2018 = ~a1950 & ~a1938;
assign a2020 = ~a2018 & ~a1948;
assign a2022 = a1940 & i46;
assign a2024 = ~a1940 & ~i46;
assign a2026 = ~a2024 & ~a2022;
assign a2028 = a2026 & ~a1696;
assign a2030 = ~a2028 & ~i48;
assign a2032 = a2028 & i48;
assign a2034 = ~a2032 & ~a2030;
assign a2036 = a2034 & ~a2020;
assign a2038 = ~a2034 & a2020;
assign a2040 = ~a2038 & ~a2036;
assign a2042 = ~a2040 & a1960;
assign a2044 = a2040 & ~a1960;
assign a2046 = ~a2044 & i10;
assign a2048 = a2046 & ~a2042;
assign a2050 = a2026 & a1708;
assign a2052 = ~a2050 & ~a2048;
assign a2054 = a2052 & ~i50;
assign a2056 = ~a2052 & i50;
assign a2058 = ~a2056 & ~a2054;
assign a2060 = a2058 & ~a2016;
assign a2062 = ~a2058 & a2016;
assign a2064 = ~a2062 & ~a2060;
assign a2066 = ~a2064 & a1984;
assign a2068 = a2064 & ~a1984;
assign a2070 = ~a2068 & i8;
assign a2072 = a2070 & ~a2066;
assign a2074 = ~a2052 & ~i8;
assign a2076 = ~a2074 & ~a2072;
assign a2078 = a2076 & ~i52;
assign a2080 = ~a2076 & i52;
assign a2082 = ~a2080 & ~a2078;
assign a2084 = a2082 & ~a2012;
assign a2086 = ~a2082 & a2012;
assign a2088 = ~a2086 & ~a2084;
assign a2090 = ~a2088 & a2008;
assign a2092 = ~a2080 & ~a2012;
assign a2094 = ~a2092 & ~a2078;
assign a2096 = ~a2056 & ~a2016;
assign a2098 = ~a2096 & ~a2054;
assign a2100 = ~a2032 & ~a2020;
assign a2102 = ~a2100 & ~a2030;
assign a2104 = a2022 & i54;
assign a2106 = ~a2022 & ~i54;
assign a2108 = ~a2106 & ~a2104;
assign a2110 = a2108 & ~a1696;
assign a2112 = ~a2110 & ~i56;
assign a2114 = a2110 & i56;
assign a2116 = ~a2114 & ~a2112;
assign a2118 = a2116 & ~a2102;
assign a2120 = ~a2116 & a2102;
assign a2122 = ~a2120 & ~a2118;
assign a2124 = ~a2122 & a2042;
assign a2126 = a2122 & ~a2042;
assign a2128 = ~a2126 & i10;
assign a2130 = a2128 & ~a2124;
assign a2132 = a2108 & a1708;
assign a2134 = ~a2132 & ~a2130;
assign a2136 = a2134 & ~i58;
assign a2138 = ~a2134 & i58;
assign a2140 = ~a2138 & ~a2136;
assign a2142 = a2140 & ~a2098;
assign a2144 = ~a2140 & a2098;
assign a2146 = ~a2144 & ~a2142;
assign a2148 = ~a2146 & a2066;
assign a2150 = a2146 & ~a2066;
assign a2152 = ~a2150 & i8;
assign a2154 = a2152 & ~a2148;
assign a2156 = ~a2134 & ~i8;
assign a2158 = ~a2156 & ~a2154;
assign a2160 = a2158 & ~i60;
assign a2162 = ~a2158 & i60;
assign a2164 = ~a2162 & ~a2160;
assign a2166 = a2164 & ~a2094;
assign a2168 = ~a2164 & a2094;
assign a2170 = ~a2168 & ~a2166;
assign a2172 = ~a2170 & a2090;
assign a2174 = a2104 & ~a1696;
assign a2176 = ~a2114 & ~a2102;
assign a2178 = ~a2176 & ~a2112;
assign a2180 = ~a2178 & ~a2174;
assign a2182 = ~a2180 & a2124;
assign a2184 = a2182 & i10;
assign a2186 = ~a2174 & ~i10;
assign a2188 = a2180 & ~a2124;
assign a2190 = ~a2188 & ~a2186;
assign a2192 = a2190 & ~a2184;
assign a2194 = ~a2138 & ~a2098;
assign a2196 = ~a2194 & ~a2136;
assign a2198 = a2196 & a2192;
assign a2200 = ~a2196 & ~a2192;
assign a2202 = ~a2200 & ~a2198;
assign a2204 = a2202 & a2148;
assign a2206 = ~a2202 & ~a2148;
assign a2208 = ~a2206 & i8;
assign a2210 = a2208 & ~a2204;
assign a2212 = a2192 & ~i8;
assign a2214 = ~a2212 & ~a2210;
assign a2216 = ~a2162 & ~a2094;
assign a2218 = ~a2216 & ~a2160;
assign a2220 = a2218 & ~a2214;
assign a2222 = ~a2218 & a2214;
assign a2224 = ~a2222 & ~a2220;
assign a2226 = a2224 & a2172;
assign a2228 = ~a2204 & ~a2198;
assign a2230 = ~a2228 & i8;
assign a2232 = ~a2230 & ~a2184;
assign a2234 = a2232 & ~a2220;
assign a2236 = ~a2234 & i62;
assign a2238 = a2236 & a2226;
assign a2240 = ~a2238 & i6;
assign a2242 = a2240 & ~l1686;
assign a2244 = l1686 & l518;
assign a2246 = ~a2244 & ~a2242;
assign a2248 = a2246 & ~a1690;
assign a2250 = ~a2248 & ~a1760;
assign a2252 = ~a2250 & a1692;
assign a2254 = a2250 & ~a1692;
assign a2256 = ~a2254 & ~a2252;
assign a2258 = ~a2256 & ~a1690;
assign a2260 = l1686 & ~l658;
assign a2262 = l508 & l506;
assign a2264 = l512 & l510;
assign a2266 = l1686 & ~l600;
assign a2268 = l1686 & ~l532;
assign a2270 = l1686 & ~l604;
assign a2272 = a2270 & l630;
assign a2274 = l1686 & ~l630;
assign a2276 = a2274 & l604;
assign a2278 = ~a2276 & ~a2272;
assign a2280 = l1686 & ~l610;
assign a2282 = a2280 & l628;
assign a2284 = l1686 & ~l628;
assign a2286 = a2284 & l610;
assign a2288 = ~a2286 & ~a2282;
assign a2290 = a2288 & a2278;
assign a2292 = l1686 & ~l624;
assign a2294 = l1686 & ~l626;
assign a2296 = l1686 & ~l492;
assign a2298 = a2296 & l612;
assign a2300 = a2298 & a2294;
assign a2302 = l1686 & ~l612;
assign a2304 = ~a2302 & ~a2296;
assign a2306 = a2304 & ~a2294;
assign a2308 = ~a2306 & ~a2300;
assign a2310 = ~a2308 & ~a2292;
assign a2312 = a2302 & a2296;
assign a2314 = a2312 & a2294;
assign a2316 = a2302 & l492;
assign a2318 = a2316 & ~a2294;
assign a2320 = ~a2318 & ~a2314;
assign a2322 = ~a2320 & a2292;
assign a2324 = ~a2322 & ~a2310;
assign a2326 = ~a2324 & a2290;
assign a2328 = ~a2326 & ~a2262;
assign a2330 = l1686 & ~l602;
assign a2332 = l1686 & ~l606;
assign a2334 = l1686 & ~l614;
assign a2336 = l1686 & ~l608;
assign a2338 = a2304 & ~a2280;
assign a2340 = a2338 & ~a2336;
assign a2342 = a2316 & ~a2280;
assign a2344 = a2342 & a2336;
assign a2346 = ~a2344 & ~a2340;
assign a2348 = ~a2346 & ~a2334;
assign a2350 = a2298 & ~a2280;
assign a2352 = ~a2350 & ~a2336;
assign a2354 = a2312 & ~a2280;
assign a2356 = ~a2354 & a2336;
assign a2358 = ~a2356 & ~a2352;
assign a2360 = a2358 & a2334;
assign a2362 = ~a2360 & ~a2348;
assign a2364 = ~a2362 & ~a2332;
assign a2366 = a2304 & a2280;
assign a2368 = ~a2366 & ~a2336;
assign a2370 = a2316 & a2280;
assign a2372 = ~a2370 & a2336;
assign a2374 = ~a2372 & ~a2368;
assign a2376 = ~a2374 & ~a2334;
assign a2378 = ~a2376 & a2332;
assign a2380 = a2298 & a2280;
assign a2382 = ~a2380 & ~a2336;
assign a2384 = a2312 & a2280;
assign a2386 = ~a2384 & a2336;
assign a2388 = ~a2386 & ~a2382;
assign a2390 = ~a2388 & a2334;
assign a2392 = ~a2390 & a2378;
assign a2394 = ~a2392 & ~a2364;
assign a2396 = ~a2394 & a2270;
assign a2398 = ~a2396 & ~a2330;
assign a2400 = a2346 & a2334;
assign a2402 = ~a2400 & ~a2376;
assign a2404 = ~a2402 & ~a2332;
assign a2406 = ~a2342 & ~a2336;
assign a2408 = ~a2350 & a2336;
assign a2410 = ~a2408 & ~a2406;
assign a2412 = ~a2410 & a2332;
assign a2414 = ~a2412 & ~a2404;
assign a2416 = a2414 & ~a2270;
assign a2418 = ~a2416 & a2330;
assign a2420 = ~a2418 & ~a2398;
assign a2422 = ~a2420 & l506;
assign a2424 = a2422 & l508;
assign a2426 = ~a2424 & ~a2328;
assign a2428 = ~a2426 & ~a2264;
assign a2430 = l1686 & ~l616;
assign a2432 = l1686 & ~l618;
assign a2434 = l1686 & ~l622;
assign a2436 = l1686 & ~l620;
assign a2438 = ~a2436 & a2338;
assign a2440 = a2436 & a2342;
assign a2442 = ~a2440 & ~a2438;
assign a2444 = ~a2442 & ~a2434;
assign a2446 = ~a2436 & ~a2350;
assign a2448 = a2436 & ~a2354;
assign a2450 = ~a2448 & ~a2446;
assign a2452 = a2450 & a2434;
assign a2454 = ~a2452 & ~a2444;
assign a2456 = ~a2454 & ~a2432;
assign a2458 = ~a2436 & ~a2380;
assign a2460 = a2436 & ~a2384;
assign a2462 = ~a2460 & ~a2458;
assign a2464 = ~a2462 & a2434;
assign a2466 = ~a2436 & ~a2366;
assign a2468 = a2436 & ~a2370;
assign a2470 = ~a2468 & ~a2466;
assign a2472 = ~a2470 & ~a2434;
assign a2474 = ~a2472 & ~a2464;
assign a2476 = a2474 & a2432;
assign a2478 = ~a2476 & ~a2456;
assign a2480 = ~a2478 & a2270;
assign a2482 = ~a2480 & ~a2430;
assign a2484 = a2442 & a2434;
assign a2486 = ~a2484 & ~a2472;
assign a2488 = ~a2486 & ~a2432;
assign a2490 = ~a2436 & ~a2342;
assign a2492 = a2436 & ~a2350;
assign a2494 = ~a2492 & ~a2490;
assign a2496 = ~a2494 & a2432;
assign a2498 = ~a2496 & ~a2488;
assign a2500 = a2498 & ~a2270;
assign a2502 = ~a2500 & a2430;
assign a2504 = ~a2502 & ~a2482;
assign a2506 = ~a2504 & ~l506;
assign a2508 = ~a2506 & ~a2422;
assign a2510 = ~a2508 & l512;
assign a2512 = a2510 & l510;
assign a2514 = ~a2512 & ~a2428;
assign a2516 = ~a2514 & a2268;
assign a2518 = ~a2516 & ~a2266;
assign a2520 = ~a2514 & ~a2268;
assign a2522 = ~a2520 & a2266;
assign a2524 = ~a2522 & ~a2518;
assign a2526 = l1686 & ~l598;
assign a2528 = a2526 & l538;
assign a2530 = a2528 & ~a2524;
assign a2532 = a2520 & ~a2266;
assign a2534 = a2516 & a2266;
assign a2536 = ~a2534 & ~a2532;
assign a2538 = a2536 & ~a2528;
assign a2540 = ~a2538 & ~a2530;
assign a2542 = l1686 & ~l596;
assign a2544 = a2542 & l540;
assign a2546 = a2544 & ~a2540;
assign a2548 = l1686 & ~l538;
assign a2550 = ~a2548 & ~a2536;
assign a2552 = a2548 & a2524;
assign a2554 = ~a2552 & ~a2550;
assign a2556 = ~a2554 & ~a2526;
assign a2558 = ~a2536 & a2526;
assign a2560 = ~a2558 & ~a2556;
assign a2562 = a2560 & ~a2544;
assign a2564 = ~a2562 & ~a2546;
assign a2566 = l1686 & ~l542;
assign a2568 = ~i70 & ~i68;
assign a2570 = ~a2568 & i72;
assign a2572 = i76 & i74;
assign a2574 = i80 & i78;
assign a2576 = a2574 & a2572;
assign a2578 = a2576 & a2570;
assign a2580 = ~a2578 & ~i82;
assign a2582 = i86 & i84;
assign a2584 = i90 & i88;
assign a2586 = a2584 & i92;
assign a2588 = a2586 & a2582;
assign a2590 = a1696 & ~i94;
assign a2592 = ~a1696 & ~i96;
assign a2594 = ~a2592 & ~a2590;
assign a2596 = a2594 & ~a2588;
assign a2598 = ~a2596 & a1712;
assign a2600 = a2598 & ~a2580;
assign a2602 = a1712 & ~i84;
assign a2604 = i98 & i82;
assign a2606 = ~i98 & ~i82;
assign a2608 = ~a2606 & ~a2604;
assign a2610 = a2608 & ~a2578;
assign a2612 = ~a2610 & a2598;
assign a2614 = a2604 & i100;
assign a2616 = ~a2604 & ~i100;
assign a2618 = ~a2616 & ~a2614;
assign a2620 = a2618 & ~a2578;
assign a2622 = ~a2620 & a2598;
assign a2624 = ~a2614 & ~i102;
assign a2626 = a2614 & i102;
assign a2628 = ~a2626 & ~a2578;
assign a2630 = a2628 & ~a2624;
assign a2632 = ~a2630 & a2598;
assign a2634 = a2626 & i70;
assign a2636 = ~a2626 & ~i70;
assign a2638 = ~a2636 & ~a2634;
assign a2640 = ~a2638 & ~a2578;
assign a2642 = a2640 & a2598;
assign a2644 = a2634 & i68;
assign a2646 = ~a2634 & ~i68;
assign a2648 = ~a2646 & ~a2578;
assign a2650 = a2648 & ~a2644;
assign a2652 = ~a2650 & a2598;
assign a2654 = a2644 & i80;
assign a2656 = ~a2644 & ~i80;
assign a2658 = ~a2656 & ~a2654;
assign a2660 = ~a2658 & ~a2578;
assign a2662 = a2660 & a2598;
assign a2664 = a2654 & i72;
assign a2666 = ~a2654 & ~i72;
assign a2668 = ~a2666 & ~a2664;
assign a2670 = ~a2668 & ~a2578;
assign a2672 = a1712 & ~i88;
assign a2674 = ~a2672 & i90;
assign a2676 = a2674 & a2598;
assign a2678 = a2670 & a2598;
assign a2680 = a2664 & i78;
assign a2682 = ~a2664 & ~i78;
assign a2684 = ~a2682 & ~a2680;
assign a2686 = ~a2684 & ~a2578;
assign a2688 = a1712 & ~i92;
assign a2690 = ~a2688 & a2676;
assign a2692 = a2686 & a2598;
assign a2694 = a2680 & i76;
assign a2696 = ~a2680 & ~i76;
assign a2698 = ~a2696 & ~a2694;
assign a2700 = ~a2698 & ~a2578;
assign a2702 = a1712 & ~i86;
assign a2704 = ~a2702 & a2690;
assign a2706 = a2700 & a2598;
assign a2708 = ~a2694 & ~i74;
assign a2710 = a2704 & ~a2602;
assign a2712 = ~a2710 & ~a2708;
assign a2714 = ~a2712 & a2602;
assign a2716 = ~a2714 & ~a2706;
assign a2718 = a2712 & ~a2602;
assign a2720 = ~a2718 & ~a2716;
assign a2722 = ~a2720 & a2704;
assign a2724 = ~a2722 & ~a2700;
assign a2726 = ~a2724 & a2602;
assign a2728 = ~a2726 & ~a2692;
assign a2730 = a2724 & ~a2602;
assign a2732 = ~a2730 & ~a2728;
assign a2734 = a2602 & i86;
assign a2736 = ~a2688 & a2674;
assign a2738 = a2736 & a2734;
assign a2740 = a2738 & ~a2720;
assign a2742 = ~a2740 & a2712;
assign a2744 = ~a2742 & a2702;
assign a2746 = ~a2744 & ~a2732;
assign a2748 = a2742 & ~a2702;
assign a2750 = ~a2748 & ~a2746;
assign a2752 = ~a2750 & a2690;
assign a2754 = a2752 & a2686;
assign a2756 = ~a2752 & ~a2686;
assign a2758 = ~a2756 & ~a2754;
assign a2760 = a2758 & a2602;
assign a2762 = ~a2760 & ~a2678;
assign a2764 = ~a2758 & ~a2602;
assign a2766 = ~a2764 & ~a2762;
assign a2768 = ~a2750 & a2736;
assign a2770 = a2768 & a2602;
assign a2772 = a2770 & ~a2724;
assign a2774 = ~a2770 & a2724;
assign a2776 = ~a2774 & ~a2772;
assign a2778 = ~a2776 & ~a2754;
assign a2780 = ~a2778 & a2702;
assign a2782 = ~a2780 & ~a2766;
assign a2784 = a2778 & ~a2702;
assign a2786 = ~a2784 & ~a2782;
assign a2788 = a2768 & a2702;
assign a2790 = ~a2788 & a2742;
assign a2792 = a2790 & ~a2772;
assign a2794 = ~a2792 & a2688;
assign a2796 = ~a2794 & ~a2786;
assign a2798 = a2792 & ~a2688;
assign a2800 = ~a2798 & ~a2796;
assign a2802 = ~a2800 & a2676;
assign a2804 = ~a2802 & ~a2670;
assign a2806 = a2802 & a2670;
assign a2808 = ~a2806 & ~a2804;
assign a2810 = a2808 & a2602;
assign a2812 = ~a2810 & ~a2662;
assign a2814 = ~a2808 & ~a2602;
assign a2816 = ~a2814 & ~a2812;
assign a2818 = ~a2800 & a2674;
assign a2820 = a2818 & a2602;
assign a2822 = a2820 & a2758;
assign a2824 = ~a2820 & ~a2758;
assign a2826 = ~a2824 & ~a2822;
assign a2828 = ~a2826 & ~a2806;
assign a2830 = a2826 & a2806;
assign a2832 = ~a2830 & ~a2828;
assign a2834 = a2832 & a2702;
assign a2836 = ~a2834 & ~a2816;
assign a2838 = ~a2832 & ~a2702;
assign a2840 = ~a2838 & ~a2836;
assign a2842 = a2818 & a2702;
assign a2844 = a2842 & ~a2778;
assign a2846 = ~a2842 & a2778;
assign a2848 = ~a2846 & ~a2844;
assign a2850 = ~a2822 & ~a2806;
assign a2852 = ~a2850 & ~a2824;
assign a2854 = ~a2852 & ~a2848;
assign a2856 = a2852 & a2848;
assign a2858 = ~a2856 & ~a2854;
assign a2860 = a2858 & a2688;
assign a2862 = ~a2860 & ~a2840;
assign a2864 = ~a2858 & ~a2688;
assign a2866 = ~a2864 & ~a2862;
assign a2868 = a2818 & a2688;
assign a2870 = ~a2868 & a2792;
assign a2872 = ~a2852 & ~a2844;
assign a2874 = ~a2872 & ~a2846;
assign a2876 = ~a2874 & a2870;
assign a2878 = ~a2876 & a2672;
assign a2880 = ~a2878 & ~a2866;
assign a2882 = a2876 & ~a2672;
assign a2884 = ~a2882 & ~a2880;
assign a2886 = ~a2884 & i90;
assign a2888 = a2886 & a2598;
assign a2890 = a2888 & a2660;
assign a2892 = ~a2888 & ~a2660;
assign a2894 = ~a2892 & ~a2890;
assign a2896 = a2894 & a2602;
assign a2898 = ~a2896 & ~a2652;
assign a2900 = ~a2894 & ~a2602;
assign a2902 = ~a2900 & ~a2898;
assign a2904 = a2886 & a2602;
assign a2906 = a2904 & a2808;
assign a2908 = ~a2904 & ~a2808;
assign a2910 = ~a2908 & ~a2906;
assign a2912 = ~a2910 & ~a2890;
assign a2914 = a2910 & a2890;
assign a2916 = ~a2914 & ~a2912;
assign a2918 = a2916 & a2702;
assign a2920 = ~a2918 & ~a2902;
assign a2922 = ~a2916 & ~a2702;
assign a2924 = ~a2922 & ~a2920;
assign a2926 = a2886 & a2702;
assign a2928 = a2926 & a2832;
assign a2930 = ~a2926 & ~a2832;
assign a2932 = ~a2930 & ~a2928;
assign a2934 = ~a2906 & ~a2890;
assign a2936 = ~a2934 & ~a2908;
assign a2938 = ~a2936 & ~a2932;
assign a2940 = a2936 & a2932;
assign a2942 = ~a2940 & ~a2938;
assign a2944 = a2942 & a2688;
assign a2946 = ~a2944 & ~a2924;
assign a2948 = ~a2942 & ~a2688;
assign a2950 = ~a2948 & ~a2946;
assign a2952 = a2886 & a2688;
assign a2954 = a2952 & a2858;
assign a2956 = ~a2952 & ~a2858;
assign a2958 = ~a2956 & ~a2954;
assign a2960 = ~a2936 & ~a2928;
assign a2962 = ~a2960 & ~a2930;
assign a2964 = ~a2962 & ~a2958;
assign a2966 = a2962 & a2958;
assign a2968 = ~a2966 & ~a2964;
assign a2970 = a2968 & a2672;
assign a2972 = ~a2970 & ~a2950;
assign a2974 = ~a2968 & ~a2672;
assign a2976 = ~a2974 & ~a2972;
assign a2978 = a1712 & ~i90;
assign a2980 = a2886 & a2672;
assign a2982 = ~a2980 & a2876;
assign a2984 = ~a2962 & ~a2954;
assign a2986 = ~a2984 & ~a2956;
assign a2988 = ~a2986 & a2982;
assign a2990 = ~a2988 & a2978;
assign a2992 = ~a2990 & ~a2976;
assign a2994 = a2988 & ~a2978;
assign a2996 = ~a2994 & ~a2992;
assign a2998 = ~a2996 & a2598;
assign a3000 = a2998 & ~a2650;
assign a3002 = ~a2998 & a2650;
assign a3004 = ~a3002 & ~a3000;
assign a3006 = a3004 & a2602;
assign a3008 = ~a3006 & ~a2642;
assign a3010 = ~a3004 & ~a2602;
assign a3012 = ~a3010 & ~a3008;
assign a3014 = ~a2996 & a2602;
assign a3016 = ~a3014 & ~a2894;
assign a3018 = a3014 & a2894;
assign a3020 = ~a3018 & ~a3016;
assign a3022 = ~a3020 & ~a3000;
assign a3024 = a3020 & a3000;
assign a3026 = ~a3024 & ~a3022;
assign a3028 = a3026 & a2702;
assign a3030 = ~a3028 & ~a3012;
assign a3032 = ~a3026 & ~a2702;
assign a3034 = ~a3032 & ~a3030;
assign a3036 = ~a2996 & a2702;
assign a3038 = a3036 & a2916;
assign a3040 = ~a3036 & ~a2916;
assign a3042 = ~a3040 & ~a3038;
assign a3044 = ~a3018 & ~a3000;
assign a3046 = ~a3044 & ~a3016;
assign a3048 = ~a3046 & ~a3042;
assign a3050 = a3046 & a3042;
assign a3052 = ~a3050 & ~a3048;
assign a3054 = a3052 & a2688;
assign a3056 = ~a3054 & ~a3034;
assign a3058 = ~a3052 & ~a2688;
assign a3060 = ~a3058 & ~a3056;
assign a3062 = ~a2996 & a2688;
assign a3064 = a3062 & a2942;
assign a3066 = ~a3062 & ~a2942;
assign a3068 = ~a3066 & ~a3064;
assign a3070 = ~a3046 & ~a3038;
assign a3072 = ~a3070 & ~a3040;
assign a3074 = ~a3072 & ~a3068;
assign a3076 = a3072 & a3068;
assign a3078 = ~a3076 & ~a3074;
assign a3080 = a3078 & a2672;
assign a3082 = ~a3080 & ~a3060;
assign a3084 = ~a3078 & ~a2672;
assign a3086 = ~a3084 & ~a3082;
assign a3088 = ~a2996 & a2672;
assign a3090 = a3088 & a2968;
assign a3092 = ~a3088 & ~a2968;
assign a3094 = ~a3092 & ~a3090;
assign a3096 = ~a3072 & ~a3064;
assign a3098 = ~a3096 & ~a3066;
assign a3100 = ~a3098 & ~a3094;
assign a3102 = a3098 & a3094;
assign a3104 = ~a3102 & ~a3100;
assign a3106 = a3104 & a2978;
assign a3108 = ~a3106 & ~a3086;
assign a3110 = ~a3104 & ~a2978;
assign a3112 = ~a2996 & a2978;
assign a3114 = ~a3112 & a2988;
assign a3116 = ~a3098 & ~a3090;
assign a3118 = ~a3116 & ~a3092;
assign a3120 = ~a3118 & a3114;
assign a3122 = ~a3120 & ~a3110;
assign a3124 = a3122 & ~a3108;
assign a3126 = ~a3124 & a2598;
assign a3128 = a3126 & a2640;
assign a3130 = ~a3126 & ~a2640;
assign a3132 = ~a3130 & ~a3128;
assign a3134 = a3132 & a2602;
assign a3136 = ~a3134 & ~a2632;
assign a3138 = ~a3132 & ~a2602;
assign a3140 = ~a3138 & ~a3136;
assign a3142 = ~a3124 & a2602;
assign a3144 = ~a3142 & ~a3004;
assign a3146 = a3142 & a3004;
assign a3148 = ~a3146 & ~a3144;
assign a3150 = ~a3148 & ~a3128;
assign a3152 = a3148 & a3128;
assign a3154 = ~a3152 & ~a3150;
assign a3156 = a3154 & a2702;
assign a3158 = ~a3156 & ~a3140;
assign a3160 = ~a3154 & ~a2702;
assign a3162 = ~a3160 & ~a3158;
assign a3164 = ~a3146 & ~a3128;
assign a3166 = ~a3164 & ~a3144;
assign a3168 = ~a3124 & a2702;
assign a3170 = ~a3168 & ~a3026;
assign a3172 = a3168 & a3026;
assign a3174 = ~a3172 & ~a3170;
assign a3176 = ~a3174 & ~a3166;
assign a3178 = a3174 & a3166;
assign a3180 = ~a3178 & ~a3176;
assign a3182 = a3180 & a2688;
assign a3184 = ~a3182 & ~a3162;
assign a3186 = ~a3180 & ~a2688;
assign a3188 = ~a3186 & ~a3184;
assign a3190 = ~a3124 & a2688;
assign a3192 = a3190 & a3052;
assign a3194 = ~a3190 & ~a3052;
assign a3196 = ~a3194 & ~a3192;
assign a3198 = ~a3172 & ~a3166;
assign a3200 = ~a3198 & ~a3170;
assign a3202 = ~a3200 & ~a3196;
assign a3204 = a3200 & a3196;
assign a3206 = ~a3204 & ~a3202;
assign a3208 = a3206 & a2672;
assign a3210 = ~a3208 & ~a3188;
assign a3212 = ~a3206 & ~a2672;
assign a3214 = ~a3212 & ~a3210;
assign a3216 = ~a3124 & a2672;
assign a3218 = a3216 & a3078;
assign a3220 = ~a3216 & ~a3078;
assign a3222 = ~a3220 & ~a3218;
assign a3224 = ~a3200 & ~a3192;
assign a3226 = ~a3224 & ~a3194;
assign a3228 = ~a3226 & ~a3222;
assign a3230 = a3226 & a3222;
assign a3232 = ~a3230 & ~a3228;
assign a3234 = a3232 & a2978;
assign a3236 = ~a3234 & ~a3214;
assign a3238 = ~a3124 & a2978;
assign a3240 = a3238 & a3104;
assign a3242 = ~a3238 & ~a3104;
assign a3244 = ~a3242 & ~a3240;
assign a3246 = ~a3226 & ~a3218;
assign a3248 = ~a3246 & ~a3220;
assign a3250 = ~a3248 & ~a3244;
assign a3252 = a3248 & a3244;
assign a3254 = ~a3232 & ~a2978;
assign a3256 = ~a3254 & ~a3252;
assign a3258 = a3256 & ~a3250;
assign a3260 = a3258 & ~a3236;
assign a3262 = ~a3260 & a2598;
assign a3264 = a3262 & ~a2630;
assign a3266 = ~a3262 & a2630;
assign a3268 = ~a3266 & ~a3264;
assign a3270 = a3268 & a2602;
assign a3272 = ~a3270 & ~a2622;
assign a3274 = ~a3268 & ~a2602;
assign a3276 = ~a3274 & ~a3272;
assign a3278 = ~a3260 & a2602;
assign a3280 = ~a3278 & ~a3132;
assign a3282 = a3278 & a3132;
assign a3284 = ~a3282 & ~a3280;
assign a3286 = ~a3284 & ~a3264;
assign a3288 = a3284 & a3264;
assign a3290 = ~a3288 & ~a3286;
assign a3292 = a3290 & a2702;
assign a3294 = ~a3292 & ~a3276;
assign a3296 = ~a3290 & ~a2702;
assign a3298 = ~a3296 & ~a3294;
assign a3300 = ~a3282 & ~a3264;
assign a3302 = ~a3300 & ~a3280;
assign a3304 = ~a3260 & a2702;
assign a3306 = ~a3304 & ~a3154;
assign a3308 = a3304 & a3154;
assign a3310 = ~a3308 & ~a3306;
assign a3312 = ~a3310 & ~a3302;
assign a3314 = a3310 & a3302;
assign a3316 = ~a3314 & ~a3312;
assign a3318 = a3316 & a2688;
assign a3320 = ~a3318 & ~a3298;
assign a3322 = ~a3316 & ~a2688;
assign a3324 = ~a3322 & ~a3320;
assign a3326 = ~a3308 & ~a3302;
assign a3328 = ~a3326 & ~a3306;
assign a3330 = ~a3260 & a2688;
assign a3332 = ~a3330 & ~a3180;
assign a3334 = a3330 & a3180;
assign a3336 = ~a3334 & ~a3332;
assign a3338 = ~a3336 & ~a3328;
assign a3340 = a3336 & a3328;
assign a3342 = ~a3340 & ~a3338;
assign a3344 = a3342 & a2672;
assign a3346 = ~a3344 & ~a3324;
assign a3348 = ~a3342 & ~a2672;
assign a3350 = ~a3348 & ~a3346;
assign a3352 = ~a3260 & a2672;
assign a3354 = a3352 & a3206;
assign a3356 = ~a3352 & ~a3206;
assign a3358 = ~a3356 & ~a3354;
assign a3360 = ~a3334 & ~a3328;
assign a3362 = ~a3360 & ~a3332;
assign a3364 = ~a3362 & ~a3358;
assign a3366 = a3362 & a3358;
assign a3368 = ~a3366 & ~a3364;
assign a3370 = a3368 & a2978;
assign a3372 = ~a3370 & ~a3350;
assign a3374 = ~a3260 & a2978;
assign a3376 = a3374 & a3232;
assign a3378 = ~a3374 & ~a3232;
assign a3380 = ~a3378 & ~a3376;
assign a3382 = ~a3362 & ~a3354;
assign a3384 = ~a3382 & ~a3356;
assign a3386 = ~a3384 & ~a3380;
assign a3388 = a3384 & a3380;
assign a3390 = ~a3368 & ~a2978;
assign a3392 = ~a3390 & ~a3388;
assign a3394 = a3392 & ~a3386;
assign a3396 = a3394 & ~a3372;
assign a3398 = ~a3396 & a2598;
assign a3400 = a3398 & ~a2620;
assign a3402 = ~a3398 & a2620;
assign a3404 = ~a3402 & ~a3400;
assign a3406 = a3404 & a2602;
assign a3408 = ~a3406 & ~a2612;
assign a3410 = ~a3404 & ~a2602;
assign a3412 = ~a3410 & ~a3408;
assign a3414 = ~a3396 & a2602;
assign a3416 = ~a3414 & ~a3268;
assign a3418 = a3414 & a3268;
assign a3420 = ~a3418 & ~a3416;
assign a3422 = ~a3420 & ~a3400;
assign a3424 = a3420 & a3400;
assign a3426 = ~a3424 & ~a3422;
assign a3428 = a3426 & a2702;
assign a3430 = ~a3428 & ~a3412;
assign a3432 = ~a3426 & ~a2702;
assign a3434 = ~a3432 & ~a3430;
assign a3436 = ~a3418 & ~a3400;
assign a3438 = ~a3436 & ~a3416;
assign a3440 = ~a3396 & a2702;
assign a3442 = ~a3440 & ~a3290;
assign a3444 = a3440 & a3290;
assign a3446 = ~a3444 & ~a3442;
assign a3448 = ~a3446 & ~a3438;
assign a3450 = a3446 & a3438;
assign a3452 = ~a3450 & ~a3448;
assign a3454 = a3452 & a2688;
assign a3456 = ~a3454 & ~a3434;
assign a3458 = ~a3452 & ~a2688;
assign a3460 = ~a3458 & ~a3456;
assign a3462 = ~a3444 & ~a3438;
assign a3464 = ~a3462 & ~a3442;
assign a3466 = ~a3396 & a2688;
assign a3468 = ~a3466 & ~a3316;
assign a3470 = a3466 & a3316;
assign a3472 = ~a3470 & ~a3468;
assign a3474 = ~a3472 & ~a3464;
assign a3476 = a3472 & a3464;
assign a3478 = ~a3476 & ~a3474;
assign a3480 = a3478 & a2672;
assign a3482 = ~a3480 & ~a3460;
assign a3484 = ~a3478 & ~a2672;
assign a3486 = ~a3484 & ~a3482;
assign a3488 = ~a3470 & ~a3464;
assign a3490 = ~a3488 & ~a3468;
assign a3492 = ~a3396 & a2672;
assign a3494 = ~a3492 & ~a3342;
assign a3496 = a3492 & a3342;
assign a3498 = ~a3496 & ~a3494;
assign a3500 = ~a3498 & ~a3490;
assign a3502 = a3498 & a3490;
assign a3504 = ~a3502 & ~a3500;
assign a3506 = a3504 & a2978;
assign a3508 = ~a3506 & ~a3486;
assign a3510 = ~a3396 & a2978;
assign a3512 = a3510 & a3368;
assign a3514 = ~a3510 & ~a3368;
assign a3516 = ~a3514 & ~a3512;
assign a3518 = ~a3496 & ~a3490;
assign a3520 = ~a3518 & ~a3494;
assign a3522 = ~a3520 & ~a3516;
assign a3524 = a3520 & a3516;
assign a3526 = ~a3524 & ~a3522;
assign a3528 = ~a3504 & ~a2978;
assign a3530 = ~a3528 & a3526;
assign a3532 = a3530 & ~a3508;
assign a3534 = ~a3532 & a2598;
assign a3536 = a3534 & ~a2610;
assign a3538 = ~a3534 & a2610;
assign a3540 = ~a3538 & ~a3536;
assign a3542 = a3540 & a2602;
assign a3544 = ~a3542 & ~a2600;
assign a3546 = ~a3540 & ~a2602;
assign a3548 = ~a3546 & ~a3544;
assign a3550 = ~a3532 & a2602;
assign a3552 = ~a3550 & ~a3404;
assign a3554 = a3550 & a3404;
assign a3556 = ~a3554 & ~a3552;
assign a3558 = ~a3556 & ~a3536;
assign a3560 = a3556 & a3536;
assign a3562 = ~a3560 & ~a3558;
assign a3564 = a3562 & a2702;
assign a3566 = ~a3564 & ~a3548;
assign a3568 = ~a3562 & ~a2702;
assign a3570 = ~a3568 & ~a3566;
assign a3572 = ~a3554 & ~a3536;
assign a3574 = ~a3572 & ~a3552;
assign a3576 = ~a3532 & a2702;
assign a3578 = ~a3576 & ~a3426;
assign a3580 = a3576 & a3426;
assign a3582 = ~a3580 & ~a3578;
assign a3584 = ~a3582 & ~a3574;
assign a3586 = a3582 & a3574;
assign a3588 = ~a3586 & ~a3584;
assign a3590 = a3588 & a2688;
assign a3592 = ~a3590 & ~a3570;
assign a3594 = ~a3588 & ~a2688;
assign a3596 = ~a3594 & ~a3592;
assign a3598 = ~a3580 & ~a3574;
assign a3600 = ~a3598 & ~a3578;
assign a3602 = ~a3532 & a2688;
assign a3604 = ~a3602 & ~a3452;
assign a3606 = a3602 & a3452;
assign a3608 = ~a3606 & ~a3604;
assign a3610 = ~a3608 & ~a3600;
assign a3612 = a3608 & a3600;
assign a3614 = ~a3612 & ~a3610;
assign a3616 = a3614 & a2672;
assign a3618 = ~a3616 & ~a3596;
assign a3620 = ~a3614 & ~a2672;
assign a3622 = ~a3620 & ~a3618;
assign a3624 = ~a3606 & ~a3600;
assign a3626 = ~a3624 & ~a3604;
assign a3628 = ~a3532 & a2672;
assign a3630 = ~a3628 & ~a3478;
assign a3632 = a3628 & a3478;
assign a3634 = ~a3632 & ~a3630;
assign a3636 = ~a3634 & ~a3626;
assign a3638 = a3634 & a3626;
assign a3640 = ~a3638 & ~a3636;
assign a3642 = a3640 & a2978;
assign a3644 = ~a3642 & ~a3622;
assign a3646 = ~a3632 & ~a3626;
assign a3648 = ~a3646 & ~a3630;
assign a3650 = ~a3532 & a2978;
assign a3652 = ~a3650 & ~a3504;
assign a3654 = a3650 & a3504;
assign a3656 = ~a3654 & ~a3652;
assign a3658 = ~a3656 & ~a3648;
assign a3660 = a3656 & a3648;
assign a3662 = ~a3660 & ~a3658;
assign a3664 = ~a3640 & ~a2978;
assign a3666 = ~a3664 & a3662;
assign a3668 = a3666 & ~a3644;
assign a3670 = ~a3668 & a2598;
assign a3672 = a3670 & ~a2580;
assign a3674 = ~a3670 & a2580;
assign a3676 = ~a3674 & ~a3672;
assign a3678 = ~a3668 & a2602;
assign a3680 = ~a3678 & ~a3540;
assign a3682 = a3678 & a3540;
assign a3684 = ~a3682 & ~a3680;
assign a3686 = ~a3684 & ~a3672;
assign a3688 = a3684 & a3672;
assign a3690 = ~a3688 & ~a3686;
assign a3692 = ~a3690 & ~a3676;
assign a3694 = ~a3682 & ~a3672;
assign a3696 = ~a3694 & ~a3680;
assign a3698 = ~a3668 & a2702;
assign a3700 = ~a3698 & ~a3562;
assign a3702 = a3698 & a3562;
assign a3704 = ~a3702 & ~a3700;
assign a3706 = ~a3704 & ~a3696;
assign a3708 = a3704 & a3696;
assign a3710 = ~a3708 & ~a3706;
assign a3712 = ~a3710 & a3692;
assign a3714 = ~a3702 & ~a3696;
assign a3716 = ~a3714 & ~a3700;
assign a3718 = ~a3668 & a2688;
assign a3720 = ~a3718 & ~a3588;
assign a3722 = a3718 & a3588;
assign a3724 = ~a3722 & ~a3720;
assign a3726 = ~a3724 & ~a3716;
assign a3728 = a3724 & a3716;
assign a3730 = ~a3728 & ~a3726;
assign a3732 = ~a3730 & a3712;
assign a3734 = ~a3722 & ~a3716;
assign a3736 = ~a3734 & ~a3720;
assign a3738 = ~a3668 & a2672;
assign a3740 = ~a3738 & ~a3614;
assign a3742 = a3738 & a3614;
assign a3744 = ~a3742 & ~a3740;
assign a3746 = ~a3744 & ~a3736;
assign a3748 = a3744 & a3736;
assign a3750 = ~a3748 & ~a3746;
assign a3752 = ~a3750 & a3732;
assign a3754 = a3750 & ~a3732;
assign a3756 = ~a3754 & ~a3752;
assign a3758 = a3756 & a1712;
assign a3760 = a3676 & a1712;
assign a3762 = i134 & ~i132;
assign a3764 = i140 & i138;
assign a3766 = a3764 & i136;
assign a3768 = a3766 & a3762;
assign a3770 = ~a3768 & i130;
assign a3772 = ~a1802 & i8;
assign a3774 = i104 & ~i8;
assign a3776 = ~a3774 & ~a3772;
assign a3778 = ~a1710 & i8;
assign a3780 = a3778 & ~a3776;
assign a3782 = ~a3780 & ~a1842;
assign a3784 = a2596 & a1790;
assign a3786 = a1860 & i84;
assign a3788 = ~a3786 & ~a3784;
assign a3790 = ~a1860 & ~i84;
assign a3792 = ~a3790 & ~a3788;
assign a3794 = a1946 & i86;
assign a3796 = ~a3794 & ~a3792;
assign a3798 = ~a1946 & ~i86;
assign a3800 = ~a3798 & ~a3796;
assign a3802 = a2028 & i92;
assign a3804 = ~a3802 & ~a3800;
assign a3806 = ~a2028 & ~i92;
assign a3808 = ~a3806 & ~a3804;
assign a3810 = a2110 & i88;
assign a3812 = ~a3810 & ~a3808;
assign a3814 = ~a2110 & ~i88;
assign a3816 = ~a3814 & ~a3812;
assign a3818 = a2174 & i90;
assign a3820 = ~a3818 & ~a3816;
assign a3822 = ~a2174 & ~i90;
assign a3824 = ~a3822 & ~a3820;
assign a3826 = a1700 & i142;
assign a3828 = a3826 & ~a3824;
assign a3830 = a3828 & ~a3782;
assign a3832 = ~a3830 & a3770;
assign a3834 = ~a3832 & a1698;
assign a3836 = ~i146 & i144;
assign a3838 = a3836 & a3824;
assign a3840 = a3838 & ~a3770;
assign a3842 = ~a3840 & a2596;
assign a3844 = ~a3770 & ~a2596;
assign a3846 = a3844 & a3838;
assign a3848 = ~a3846 & ~a1698;
assign a3850 = a3848 & ~a3842;
assign a3852 = ~a3850 & ~a3834;
assign a3854 = a1738 & ~a1716;
assign a3856 = a3854 & ~a3838;
assign a3858 = a3856 & ~a3852;
assign a3860 = a3838 & ~a2596;
assign a3862 = ~a3860 & ~a3830;
assign a3864 = a3862 & ~a3858;
assign a3866 = ~a1814 & ~a1700;
assign a3868 = ~a3866 & ~a1842;
assign a3870 = ~a3868 & a3864;
assign a3872 = a3830 & ~a3770;
assign a3874 = ~a1886 & i8;
assign a3876 = i106 & ~i8;
assign a3878 = ~a3876 & ~a3874;
assign a3880 = ~a3878 & a3778;
assign a3882 = a1858 & a1700;
assign a3884 = ~a3882 & ~a3880;
assign a3886 = ~a3884 & a3828;
assign a3888 = ~a3886 & i136;
assign a3890 = a3886 & ~i136;
assign a3892 = ~a3890 & ~a3888;
assign a3894 = a3892 & ~a3872;
assign a3896 = ~a3892 & a3872;
assign a3898 = ~a3896 & ~a3894;
assign a3900 = ~a3898 & a1698;
assign a3902 = ~i136 & ~i84;
assign a3904 = i136 & i84;
assign a3906 = ~a3904 & ~a3902;
assign a3908 = a3906 & a3844;
assign a3910 = ~a3906 & ~a3844;
assign a3912 = ~a3910 & ~a3908;
assign a3914 = a3912 & a3838;
assign a3916 = ~a3838 & ~i84;
assign a3918 = ~a3916 & ~a3914;
assign a3920 = ~a3918 & ~a1698;
assign a3922 = ~a3920 & ~a3900;
assign a3924 = ~a3922 & a3856;
assign a3926 = a3838 & ~i84;
assign a3928 = ~a3926 & ~a3886;
assign a3930 = a3928 & ~a3924;
assign a3932 = ~a1912 & ~a1700;
assign a3934 = ~a3932 & ~a3882;
assign a3936 = ~a3934 & a3930;
assign a3938 = ~a3936 & ~a3870;
assign a3940 = a3934 & ~a3930;
assign a3942 = ~a3940 & ~a3938;
assign a3944 = ~a3890 & ~a3872;
assign a3946 = ~a3944 & ~a3888;
assign a3948 = ~a1970 & i8;
assign a3950 = i108 & ~i8;
assign a3952 = ~a3950 & ~a3948;
assign a3954 = ~a3952 & a3778;
assign a3956 = a1944 & a1700;
assign a3958 = ~a3956 & ~a3954;
assign a3960 = ~a3958 & a3828;
assign a3962 = ~a3960 & i134;
assign a3964 = a3960 & ~i134;
assign a3966 = ~a3964 & ~a3962;
assign a3968 = a3966 & ~a3946;
assign a3970 = ~a3966 & a3946;
assign a3972 = ~a3970 & ~a3968;
assign a3974 = ~a3972 & a1698;
assign a3976 = ~a3902 & ~a3844;
assign a3978 = ~a3976 & ~a3904;
assign a3980 = ~i134 & ~i86;
assign a3982 = i134 & i86;
assign a3984 = ~a3982 & ~a3980;
assign a3986 = a3984 & a3978;
assign a3988 = ~a3984 & ~a3978;
assign a3990 = ~a3988 & ~a3986;
assign a3992 = a3990 & a3838;
assign a3994 = ~a3838 & ~i86;
assign a3996 = ~a3994 & ~a3992;
assign a3998 = ~a3996 & ~a1698;
assign a4000 = ~a3998 & ~a3974;
assign a4002 = ~a4000 & a3856;
assign a4004 = a3838 & ~i86;
assign a4006 = ~a4004 & ~a3960;
assign a4008 = a4006 & ~a4002;
assign a4010 = ~a1994 & ~a1700;
assign a4012 = ~a4010 & ~a3956;
assign a4014 = ~a4012 & a4008;
assign a4016 = ~a4014 & ~a3942;
assign a4018 = a4012 & ~a4008;
assign a4020 = ~a4018 & ~a4016;
assign a4022 = ~a3964 & ~a3946;
assign a4024 = ~a4022 & ~a3962;
assign a4026 = ~a2052 & i8;
assign a4028 = i110 & ~i8;
assign a4030 = ~a4028 & ~a4026;
assign a4032 = ~a4030 & a3778;
assign a4034 = a2026 & a1700;
assign a4036 = ~a4034 & ~a4032;
assign a4038 = ~a4036 & a3828;
assign a4040 = ~a4038 & i138;
assign a4042 = a4038 & ~i138;
assign a4044 = ~a4042 & ~a4040;
assign a4046 = a4044 & ~a4024;
assign a4048 = ~a4044 & a4024;
assign a4050 = ~a4048 & ~a4046;
assign a4052 = ~a4050 & a1698;
assign a4054 = ~a3980 & ~a3978;
assign a4056 = ~a4054 & ~a3982;
assign a4058 = ~i138 & ~i92;
assign a4060 = i138 & i92;
assign a4062 = ~a4060 & ~a4058;
assign a4064 = a4062 & a4056;
assign a4066 = ~a4062 & ~a4056;
assign a4068 = ~a4066 & ~a4064;
assign a4070 = a4068 & a3838;
assign a4072 = ~a3838 & ~i92;
assign a4074 = ~a4072 & ~a4070;
assign a4076 = ~a4074 & ~a1698;
assign a4078 = ~a4076 & ~a4052;
assign a4080 = ~a4078 & a3856;
assign a4082 = a3838 & ~i92;
assign a4084 = ~a4082 & ~a4038;
assign a4086 = a4084 & ~a4080;
assign a4088 = ~a2076 & ~a1700;
assign a4090 = ~a4088 & ~a4034;
assign a4092 = ~a4090 & a4086;
assign a4094 = ~a4092 & ~a4020;
assign a4096 = a4090 & ~a4086;
assign a4098 = ~a4096 & ~a4094;
assign a4100 = ~a4042 & ~a4024;
assign a4102 = ~a4100 & ~a4040;
assign a4104 = ~a2134 & i8;
assign a4106 = i112 & ~i8;
assign a4108 = ~a4106 & ~a4104;
assign a4110 = ~a4108 & a3778;
assign a4112 = a2108 & a1700;
assign a4114 = ~a4112 & ~a4110;
assign a4116 = ~a4114 & a3828;
assign a4118 = ~a4116 & i140;
assign a4120 = a4116 & ~i140;
assign a4122 = ~a4120 & ~a4118;
assign a4124 = a4122 & ~a4102;
assign a4126 = ~a4122 & a4102;
assign a4128 = ~a4126 & ~a4124;
assign a4130 = ~a4128 & a1698;
assign a4132 = ~a4058 & ~a4056;
assign a4134 = ~a4132 & ~a4060;
assign a4136 = ~i140 & ~i88;
assign a4138 = i140 & i88;
assign a4140 = ~a4138 & ~a4136;
assign a4142 = a4140 & a4134;
assign a4144 = ~a4140 & ~a4134;
assign a4146 = ~a4144 & ~a4142;
assign a4148 = a4146 & a3838;
assign a4150 = ~a3838 & ~i88;
assign a4152 = ~a4150 & ~a4148;
assign a4154 = ~a4152 & ~a1698;
assign a4156 = ~a4154 & ~a4130;
assign a4158 = ~a4156 & a3856;
assign a4160 = a3838 & ~i88;
assign a4162 = ~a4160 & ~a4116;
assign a4164 = a4162 & ~a4158;
assign a4166 = ~a2158 & ~a1700;
assign a4168 = ~a4166 & ~a4112;
assign a4170 = ~a4168 & a4164;
assign a4172 = ~a4170 & ~a4098;
assign a4174 = a4168 & ~a4164;
assign a4176 = ~a4174 & ~a4172;
assign a4178 = a2192 & i8;
assign a4180 = i114 & ~i8;
assign a4182 = ~a4180 & ~a4178;
assign a4184 = ~a4182 & a3778;
assign a4186 = a2104 & a1700;
assign a4188 = ~a4186 & ~a4184;
assign a4190 = ~a4188 & a3828;
assign a4192 = ~a4120 & ~a4102;
assign a4194 = ~a4192 & ~a4118;
assign a4196 = a4190 & ~i132;
assign a4198 = ~a4190 & i132;
assign a4200 = ~a4198 & ~a4196;
assign a4202 = ~a4200 & ~a4194;
assign a4204 = a4200 & a4194;
assign a4206 = ~a4204 & ~a4202;
assign a4208 = ~a4206 & a1698;
assign a4210 = ~a4136 & ~a4134;
assign a4212 = ~a4210 & ~a4138;
assign a4214 = a4212 & ~i132;
assign a4216 = ~a4212 & i132;
assign a4218 = ~a4216 & ~a4214;
assign a4220 = ~a4218 & a3838;
assign a4222 = ~a4220 & i90;
assign a4224 = ~a4222 & ~a1698;
assign a4226 = ~a4224 & ~a4208;
assign a4228 = ~a4226 & a3856;
assign a4230 = ~a4228 & ~a4190;
assign a4232 = ~a2214 & ~a1700;
assign a4234 = ~a4232 & ~a4186;
assign a4236 = ~a4234 & a4230;
assign a4238 = ~a4236 & ~a4176;
assign a4240 = a4234 & ~a4230;
assign a4242 = ~a4240 & ~a4238;
assign a4244 = ~a2232 & ~a1700;
assign a4246 = ~a4244 & ~a4242;
assign a4248 = ~a4246 & ~a3864;
assign a4250 = a4246 & a3868;
assign a4252 = ~a4250 & ~a4248;
assign a4254 = a4252 & a3760;
assign a4256 = a3690 & a3676;
assign a4258 = ~a4256 & ~a3692;
assign a4260 = a4258 & a1712;
assign a4262 = ~a4246 & ~a3930;
assign a4264 = a3934 & a3868;
assign a4266 = ~a3934 & ~a3868;
assign a4268 = ~a4266 & ~a4264;
assign a4270 = ~a4268 & a4246;
assign a4272 = ~a4270 & ~a4262;
assign a4274 = a4272 & a4260;
assign a4276 = ~a4274 & ~a4254;
assign a4278 = ~a4272 & ~a4260;
assign a4280 = ~a4278 & ~a4276;
assign a4282 = a3710 & ~a3692;
assign a4284 = ~a4282 & ~a3712;
assign a4286 = a4284 & a1712;
assign a4288 = ~a4246 & ~a4008;
assign a4290 = a4264 & a4012;
assign a4292 = ~a4264 & ~a4012;
assign a4294 = ~a4292 & ~a4290;
assign a4296 = ~a4294 & a4246;
assign a4298 = ~a4296 & ~a4288;
assign a4300 = a4298 & a4286;
assign a4302 = ~a4300 & ~a4280;
assign a4304 = ~a4298 & ~a4286;
assign a4306 = ~a4304 & ~a4302;
assign a4308 = a3730 & ~a3712;
assign a4310 = ~a4308 & ~a3732;
assign a4312 = a4310 & a1712;
assign a4314 = ~a4246 & ~a4086;
assign a4316 = a4290 & a4090;
assign a4318 = ~a4290 & ~a4090;
assign a4320 = ~a4318 & ~a4316;
assign a4322 = ~a4320 & a4246;
assign a4324 = ~a4322 & ~a4314;
assign a4326 = a4324 & a4312;
assign a4328 = ~a4326 & ~a4306;
assign a4330 = ~a4324 & ~a4312;
assign a4332 = ~a4330 & ~a4328;
assign a4334 = ~a4246 & ~a4164;
assign a4336 = a4316 & a4168;
assign a4338 = ~a4316 & ~a4168;
assign a4340 = ~a4338 & ~a4336;
assign a4342 = ~a4340 & a4246;
assign a4344 = ~a4342 & ~a4334;
assign a4346 = a4344 & a3758;
assign a4348 = ~a4346 & ~a4332;
assign a4350 = ~a4344 & ~a3758;
assign a4352 = ~a4350 & ~a4348;
assign a4354 = ~a3742 & ~a3736;
assign a4356 = ~a4354 & ~a3740;
assign a4358 = ~a3668 & a2978;
assign a4360 = ~a4358 & ~a3640;
assign a4362 = a4358 & a3640;
assign a4364 = ~a4362 & ~a4360;
assign a4366 = ~a4364 & ~a4356;
assign a4368 = a4364 & a4356;
assign a4370 = ~a4368 & ~a4366;
assign a4372 = ~a4370 & ~a3752;
assign a4374 = a4370 & a3752;
assign a4376 = ~a4374 & ~a4372;
assign a4378 = ~a4376 & a1712;
assign a4380 = a1766 & i148;
assign a4382 = a4380 & ~a4378;
assign a4384 = a4382 & ~a4352;
assign a4386 = ~i152 & ~i150;
assign a4388 = a4386 & a3838;
assign a4390 = a4388 & a4384;
assign a4392 = a4390 & a3758;
assign a4394 = ~a4392 & ~l1686;
assign a4396 = l1686 & l594;
assign a4398 = ~a4396 & ~a4394;
assign a4400 = a4398 & ~a2566;
assign a4402 = a4400 & ~a2564;
assign a4404 = l1686 & ~l540;
assign a4406 = ~a4404 & ~a2560;
assign a4408 = ~a2526 & ~a2524;
assign a4410 = a2554 & a2526;
assign a4412 = ~a4410 & ~a4408;
assign a4414 = a4412 & a4404;
assign a4416 = ~a4414 & ~a4406;
assign a4418 = ~a4416 & ~a2542;
assign a4420 = ~a2560 & a2542;
assign a4422 = ~a4420 & ~a4418;
assign a4424 = a4422 & ~a4400;
assign a4426 = ~a4424 & ~a4402;
assign a4428 = l1686 & ~l544;
assign a4430 = a4390 & a4312;
assign a4432 = ~a4430 & ~l1686;
assign a4434 = l1686 & l592;
assign a4436 = ~a4434 & ~a4432;
assign a4438 = a4436 & ~a4428;
assign a4440 = a4438 & ~a4426;
assign a4442 = ~a4422 & ~a2566;
assign a4444 = ~a4412 & ~a2542;
assign a4446 = a4416 & a2542;
assign a4448 = ~a4446 & ~a4444;
assign a4450 = a4448 & a2566;
assign a4452 = ~a4450 & ~a4442;
assign a4454 = ~a4452 & ~a4398;
assign a4456 = ~a4422 & a4398;
assign a4458 = ~a4456 & ~a4454;
assign a4460 = a4458 & ~a4438;
assign a4462 = ~a4460 & ~a4440;
assign a4464 = l1686 & ~l546;
assign a4466 = a4390 & a4286;
assign a4468 = ~a4466 & ~l1686;
assign a4470 = l1686 & l590;
assign a4472 = ~a4470 & ~a4468;
assign a4474 = a4472 & ~a4464;
assign a4476 = a4474 & ~a4462;
assign a4478 = ~a4458 & ~a4428;
assign a4480 = ~a4448 & ~a4398;
assign a4482 = a4452 & a4398;
assign a4484 = ~a4482 & ~a4480;
assign a4486 = a4484 & a4428;
assign a4488 = ~a4486 & ~a4478;
assign a4490 = ~a4488 & ~a4436;
assign a4492 = ~a4458 & a4436;
assign a4494 = ~a4492 & ~a4490;
assign a4496 = a4494 & ~a4474;
assign a4498 = ~a4496 & ~a4476;
assign a4500 = l1686 & ~l520;
assign a4502 = a4390 & a4260;
assign a4504 = ~a4502 & ~l1686;
assign a4506 = l1686 & l588;
assign a4508 = ~a4506 & ~a4504;
assign a4510 = a4508 & ~a4500;
assign a4512 = a4510 & ~a4498;
assign a4514 = ~a4494 & ~a4464;
assign a4516 = ~a4484 & ~a4436;
assign a4518 = a4488 & a4436;
assign a4520 = ~a4518 & ~a4516;
assign a4522 = a4520 & a4464;
assign a4524 = ~a4522 & ~a4514;
assign a4526 = ~a4524 & ~a4472;
assign a4528 = ~a4494 & a4472;
assign a4530 = ~a4528 & ~a4526;
assign a4532 = a4530 & ~a4510;
assign a4534 = ~a4532 & ~a4512;
assign a4536 = l1686 & ~l548;
assign a4538 = a4390 & a3760;
assign a4540 = ~a4538 & ~l1686;
assign a4542 = l1686 & l640;
assign a4544 = ~a4542 & ~a4540;
assign a4546 = a4544 & ~a4536;
assign a4548 = a4546 & ~a4534;
assign a4550 = ~a4520 & ~a4472;
assign a4552 = a4524 & a4472;
assign a4554 = ~a4552 & ~a4550;
assign a4556 = ~a4508 & a4500;
assign a4558 = a4556 & ~a4554;
assign a4560 = ~a4556 & a4530;
assign a4562 = ~a4560 & ~a4558;
assign a4564 = ~a4562 & ~a4546;
assign a4566 = ~a4564 & ~a4548;
assign a4568 = a4566 & a1690;
assign a4570 = a2338 & ~a1694;
assign a4572 = a2350 & a1694;
assign a4574 = ~a4572 & ~a4570;
assign a4576 = ~a4574 & ~a1726;
assign a4578 = ~a2342 & ~a1694;
assign a4580 = ~a2354 & a1694;
assign a4582 = ~a4580 & ~a4578;
assign a4584 = a4582 & a1726;
assign a4586 = ~a4584 & ~a4576;
assign a4588 = ~a4586 & ~a1746;
assign a4590 = ~a2366 & ~a1694;
assign a4592 = ~a2380 & a1694;
assign a4594 = ~a4592 & ~a4590;
assign a4596 = ~a4594 & ~a1726;
assign a4598 = ~a2370 & ~a1694;
assign a4600 = ~a2384 & a1694;
assign a4602 = ~a4600 & ~a4598;
assign a4604 = ~a4602 & a1726;
assign a4606 = ~a4604 & ~a4596;
assign a4608 = a4606 & a1746;
assign a4610 = ~a4608 & ~a4588;
assign a4612 = ~a4610 & a2270;
assign a4614 = ~a4612 & ~a1736;
assign a4616 = ~a2338 & a1694;
assign a4618 = ~a4616 & ~a4590;
assign a4620 = ~a4618 & ~a1726;
assign a4622 = ~a4620 & ~a4604;
assign a4624 = ~a4622 & ~a1746;
assign a4626 = ~a4582 & ~a1726;
assign a4628 = ~a2350 & ~a1694;
assign a4630 = ~a4628 & ~a4616;
assign a4632 = ~a4630 & a1726;
assign a4634 = ~a4632 & ~a4626;
assign a4636 = ~a4634 & a1746;
assign a4638 = ~a4636 & ~a4624;
assign a4640 = a4638 & ~a2270;
assign a4642 = ~a4640 & a1736;
assign a4644 = ~a4642 & ~a4614;
assign a4646 = ~a1928 & i62;
assign a4648 = ~a1814 & ~i62;
assign a4650 = ~a4648 & ~a4646;
assign a4652 = a4650 & ~l1686;
assign a4654 = l1686 & l550;
assign a4656 = ~a4654 & ~a4652;
assign a4658 = ~a1928 & a1924;
assign a4660 = ~a1930 & i62;
assign a4662 = a4660 & ~a4658;
assign a4664 = ~a1912 & ~i62;
assign a4666 = ~a4664 & ~a4662;
assign a4668 = a4666 & ~l1686;
assign a4670 = l1686 & l522;
assign a4672 = ~a4670 & ~a4668;
assign a4674 = ~a4672 & a4500;
assign a4676 = a2006 & ~a1930;
assign a4678 = ~a2008 & i62;
assign a4680 = a4678 & ~a4676;
assign a4682 = ~a1994 & ~i62;
assign a4684 = ~a4682 & ~a4680;
assign a4686 = a4684 & ~l1686;
assign a4688 = l1686 & l524;
assign a4690 = ~a4688 & ~a4686;
assign a4692 = a2088 & ~a2008;
assign a4694 = ~a2090 & i62;
assign a4696 = a4694 & ~a4692;
assign a4698 = ~a2076 & ~i62;
assign a4700 = ~a4698 & ~a4696;
assign a4702 = a4700 & ~l1686;
assign a4704 = l1686 & l526;
assign a4706 = ~a4704 & ~a4702;
assign a4708 = a2170 & ~a2090;
assign a4710 = ~a2172 & i62;
assign a4712 = a4710 & ~a4708;
assign a4714 = ~a2158 & ~i62;
assign a4716 = ~a4714 & ~a4712;
assign a4718 = a4716 & ~l1686;
assign a4720 = l1686 & l528;
assign a4722 = ~a4720 & ~a4718;
assign a4724 = ~a2224 & ~a2172;
assign a4726 = ~a2226 & i62;
assign a4728 = a4726 & ~a4724;
assign a4730 = ~a2214 & ~i62;
assign a4732 = ~a4730 & ~a4728;
assign a4734 = a4732 & ~l1686;
assign a4736 = l1686 & l530;
assign a4738 = ~a4736 & ~a4734;
assign a4740 = a2232 & ~i62;
assign a4742 = a2234 & ~a2226;
assign a4744 = ~a4742 & ~a4740;
assign a4746 = a4744 & ~a2238;
assign a4748 = ~a4746 & ~l1686;
assign a4750 = l1686 & l536;
assign a4752 = ~a4750 & ~a4748;
assign a4754 = a4752 & ~a2548;
assign a4756 = ~a2238 & ~l1686;
assign a4758 = l1686 & l534;
assign a4760 = ~a4758 & ~a4756;
assign a4762 = ~a4760 & ~a2268;
assign a4764 = a4760 & a2268;
assign a4766 = ~a4764 & ~a4762;
assign a4768 = a4766 & a4754;
assign a4770 = ~a4752 & a2548;
assign a4772 = a4770 & ~a4766;
assign a4774 = ~a4772 & ~a4768;
assign a4776 = a4774 & a4404;
assign a4778 = ~a4770 & a4766;
assign a4780 = ~a4778 & ~a4772;
assign a4782 = a4780 & ~a4404;
assign a4784 = ~a4782 & ~a4776;
assign a4786 = ~a4784 & ~a4738;
assign a4788 = a4778 & ~a4754;
assign a4790 = ~a4788 & ~a4404;
assign a4792 = ~a4790 & ~a4780;
assign a4794 = ~a4792 & a4738;
assign a4796 = ~a4794 & ~a4786;
assign a4798 = ~a4796 & ~a2566;
assign a4800 = a4774 & ~a4404;
assign a4802 = ~a4766 & ~a4754;
assign a4804 = ~a4802 & ~a4768;
assign a4806 = a4804 & a4404;
assign a4808 = ~a4806 & ~a4800;
assign a4810 = ~a4808 & ~a4738;
assign a4812 = ~a4784 & a4738;
assign a4814 = ~a4812 & ~a4810;
assign a4816 = ~a4814 & a2566;
assign a4818 = ~a4816 & ~a4798;
assign a4820 = ~a4818 & ~a4722;
assign a4822 = ~a4796 & a4722;
assign a4824 = ~a4822 & ~a4820;
assign a4826 = ~a4824 & ~a4428;
assign a4828 = ~a4814 & ~a4722;
assign a4830 = ~a4818 & a4722;
assign a4832 = ~a4830 & ~a4828;
assign a4834 = ~a4832 & a4428;
assign a4836 = ~a4834 & ~a4826;
assign a4838 = ~a4836 & ~a4706;
assign a4840 = ~a4824 & a4706;
assign a4842 = ~a4840 & ~a4838;
assign a4844 = ~a4842 & ~a4464;
assign a4846 = ~a4832 & ~a4706;
assign a4848 = ~a4836 & a4706;
assign a4850 = ~a4848 & ~a4846;
assign a4852 = ~a4850 & a4464;
assign a4854 = ~a4852 & ~a4844;
assign a4856 = ~a4854 & ~a4690;
assign a4858 = ~a4842 & a4690;
assign a4860 = ~a4858 & ~a4856;
assign a4862 = ~a4860 & ~a4674;
assign a4864 = ~a4850 & ~a4690;
assign a4866 = ~a4854 & a4690;
assign a4868 = ~a4866 & ~a4864;
assign a4870 = ~a4868 & ~a4672;
assign a4872 = a4870 & a4500;
assign a4874 = ~a4872 & ~a4862;
assign a4876 = ~a4874 & ~a4656;
assign a4878 = ~a4860 & ~a4672;
assign a4880 = ~a4806 & ~a4782;
assign a4882 = ~a4880 & ~a4738;
assign a4884 = a4780 & a4738;
assign a4886 = ~a4884 & ~a4882;
assign a4888 = ~a4886 & ~a2566;
assign a4890 = ~a4888 & ~a4816;
assign a4892 = ~a4890 & ~a4722;
assign a4894 = ~a4886 & a2566;
assign a4896 = ~a4894 & ~a4798;
assign a4898 = ~a4896 & a4722;
assign a4900 = ~a4898 & ~a4892;
assign a4902 = ~a4900 & ~a4428;
assign a4904 = ~a4902 & ~a4834;
assign a4906 = ~a4904 & ~a4706;
assign a4908 = ~a4900 & a4428;
assign a4910 = ~a4908 & ~a4826;
assign a4912 = ~a4910 & a4706;
assign a4914 = ~a4912 & ~a4906;
assign a4916 = ~a4914 & a4464;
assign a4918 = ~a4916 & ~a4844;
assign a4920 = ~a4918 & ~a4690;
assign a4922 = ~a4910 & ~a4706;
assign a4924 = ~a4896 & ~a4722;
assign a4926 = a4738 & ~a4404;
assign a4928 = a4926 & ~a4804;
assign a4930 = ~a4926 & a4780;
assign a4932 = ~a4930 & ~a4928;
assign a4934 = ~a4932 & ~a2566;
assign a4936 = ~a4796 & a2566;
assign a4938 = ~a4936 & ~a4934;
assign a4940 = ~a4938 & a4722;
assign a4942 = ~a4940 & ~a4924;
assign a4944 = ~a4942 & ~a4428;
assign a4946 = ~a4824 & a4428;
assign a4948 = ~a4946 & ~a4944;
assign a4950 = ~a4948 & a4706;
assign a4952 = ~a4950 & ~a4922;
assign a4954 = ~a4952 & ~a4464;
assign a4956 = ~a4842 & a4464;
assign a4958 = ~a4956 & ~a4954;
assign a4960 = ~a4958 & a4690;
assign a4962 = ~a4960 & ~a4920;
assign a4964 = ~a4962 & a4672;
assign a4966 = ~a4964 & ~a4878;
assign a4968 = ~a4966 & ~a4500;
assign a4970 = ~a4914 & ~a4464;
assign a4972 = ~a4970 & ~a4852;
assign a4974 = ~a4972 & ~a4690;
assign a4976 = ~a4918 & a4690;
assign a4978 = ~a4976 & ~a4974;
assign a4980 = ~a4978 & ~a4672;
assign a4982 = ~a4860 & a4672;
assign a4984 = ~a4982 & ~a4980;
assign a4986 = ~a4984 & a4500;
assign a4988 = ~a4986 & ~a4968;
assign a4990 = ~a4988 & a4656;
assign a4992 = ~a4990 & ~a4876;
assign a4994 = ~a4992 & ~a4536;
assign a4996 = ~a4984 & ~a4500;
assign a4998 = ~a4978 & a4672;
assign a5000 = ~a4998 & ~a4870;
assign a5002 = ~a5000 & a4500;
assign a5004 = ~a5002 & ~a4996;
assign a5006 = ~a5004 & ~a4656;
assign a5008 = ~a4874 & a4656;
assign a5010 = ~a5008 & ~a5006;
assign a5012 = ~a5010 & a4536;
assign a5014 = ~a5012 & ~a4994;
assign a5016 = ~a5014 & ~a2246;
assign a5018 = a5016 & ~a4644;
assign a5020 = ~a4610 & ~a2270;
assign a5022 = a5020 & ~a1736;
assign a5024 = a4612 & a1736;
assign a5026 = ~a5024 & ~a5022;
assign a5028 = ~a4804 & ~a4738;
assign a5030 = a4880 & a4738;
assign a5032 = ~a5030 & ~a5028;
assign a5034 = ~a5032 & ~a4722;
assign a5036 = a5032 & a2566;
assign a5038 = ~a5036 & ~a4888;
assign a5040 = a5038 & a4722;
assign a5042 = ~a5040 & ~a5034;
assign a5044 = ~a5042 & ~a4706;
assign a5046 = ~a5038 & ~a4722;
assign a5048 = ~a4886 & a4722;
assign a5050 = ~a5048 & ~a5046;
assign a5052 = ~a5050 & ~a4428;
assign a5054 = a5042 & a4428;
assign a5056 = ~a5054 & ~a5052;
assign a5058 = a5056 & a4706;
assign a5060 = ~a5058 & ~a5044;
assign a5062 = ~a5060 & ~a4690;
assign a5064 = ~a5056 & ~a4706;
assign a5066 = ~a5050 & a4706;
assign a5068 = ~a5066 & ~a5064;
assign a5070 = ~a5068 & ~a4464;
assign a5072 = a5060 & a4464;
assign a5074 = ~a5072 & ~a5070;
assign a5076 = a5074 & a4690;
assign a5078 = ~a5076 & ~a5062;
assign a5080 = ~a5078 & ~a4672;
assign a5082 = ~a5074 & ~a4690;
assign a5084 = ~a5068 & a4690;
assign a5086 = ~a5084 & ~a5082;
assign a5088 = a5086 & a4672;
assign a5090 = ~a5088 & ~a5080;
assign a5092 = ~a5090 & ~a4500;
assign a5094 = ~a5078 & a4500;
assign a5096 = ~a5094 & ~a5092;
assign a5098 = ~a4656 & a4536;
assign a5100 = a5098 & ~a5096;
assign a5102 = ~a5086 & ~a4500;
assign a5104 = ~a5102 & ~a5098;
assign a5106 = a5090 & a4500;
assign a5108 = ~a5106 & a5104;
assign a5110 = ~a5108 & ~a5100;
assign a5112 = a5110 & a2246;
assign a5114 = a5112 & a5026;
assign a5116 = ~a5114 & ~a5018;
assign a5118 = ~a5116 & ~a1690;
assign a5120 = ~a5118 & ~a4568;
assign a5122 = ~a5120 & ~l494;
assign a5124 = l1686 & ~l500;
assign a5126 = l1686 & ~l498;
assign a5128 = l1686 & ~l502;
assign a5130 = l1686 & ~l496;
assign a5132 = ~a5130 & a2338;
assign a5134 = a5130 & a2342;
assign a5136 = ~a5134 & ~a5132;
assign a5138 = ~a5136 & ~a5128;
assign a5140 = ~a5130 & ~a2350;
assign a5142 = a5130 & ~a2354;
assign a5144 = ~a5142 & ~a5140;
assign a5146 = a5144 & a5128;
assign a5148 = ~a5146 & ~a5138;
assign a5150 = ~a5148 & ~a5126;
assign a5152 = ~a5130 & ~a2380;
assign a5154 = a5130 & ~a2384;
assign a5156 = ~a5154 & ~a5152;
assign a5158 = ~a5156 & a5128;
assign a5160 = ~a5130 & ~a2366;
assign a5162 = a5130 & ~a2370;
assign a5164 = ~a5162 & ~a5160;
assign a5166 = ~a5164 & ~a5128;
assign a5168 = ~a5166 & ~a5158;
assign a5170 = a5168 & a5126;
assign a5172 = ~a5170 & ~a5150;
assign a5174 = ~a5172 & a2270;
assign a5176 = ~a5174 & ~a5124;
assign a5178 = a5136 & a5128;
assign a5180 = ~a5178 & ~a5166;
assign a5182 = ~a5180 & ~a5126;
assign a5184 = ~a5130 & ~a2342;
assign a5186 = a5130 & ~a2350;
assign a5188 = ~a5186 & ~a5184;
assign a5190 = ~a5188 & a5126;
assign a5192 = ~a5190 & ~a5182;
assign a5194 = a5192 & ~a2270;
assign a5196 = ~a5194 & a5124;
assign a5198 = ~a5196 & ~a5176;
assign a5200 = ~a1814 & ~a1704;
assign a5202 = ~a5200 & a3782;
assign a5204 = a5202 & a3760;
assign a5206 = ~a1912 & ~a1704;
assign a5208 = ~a5206 & a3884;
assign a5210 = a5208 & a4260;
assign a5212 = ~a5210 & ~a5204;
assign a5214 = ~a5208 & ~a4260;
assign a5216 = ~a5214 & ~a5212;
assign a5218 = ~a1994 & ~a1704;
assign a5220 = ~a5218 & a3958;
assign a5222 = a5220 & a4286;
assign a5224 = ~a5222 & ~a5216;
assign a5226 = ~a5220 & ~a4286;
assign a5228 = ~a5226 & ~a5224;
assign a5230 = ~a2076 & ~a1704;
assign a5232 = ~a5230 & a4036;
assign a5234 = a5232 & a4312;
assign a5236 = ~a5234 & ~a5228;
assign a5238 = ~a5232 & ~a4312;
assign a5240 = ~a5238 & ~a5236;
assign a5242 = ~a2158 & ~a1704;
assign a5244 = ~a5242 & a4114;
assign a5246 = a5244 & a3758;
assign a5248 = ~a5246 & ~a5240;
assign a5250 = ~a5244 & ~a3758;
assign a5252 = ~a5250 & ~a5248;
assign a5254 = ~a2214 & ~a1704;
assign a5256 = ~a5254 & a4188;
assign a5258 = a5256 & a4378;
assign a5260 = ~a5258 & ~a5252;
assign a5262 = ~a5256 & ~a4378;
assign a5264 = ~a5262 & ~a5260;
assign a5266 = ~a5264 & a3760;
assign a5268 = a5264 & ~a5202;
assign a5270 = ~a5268 & ~a5266;
assign a5272 = ~a5270 & ~i66;
assign a5274 = ~a5264 & a1712;
assign a5276 = a5274 & a4258;
assign a5278 = a5264 & ~a5208;
assign a5280 = ~a5278 & ~a5276;
assign a5282 = ~a5280 & ~i64;
assign a5284 = ~a5282 & ~a5272;
assign a5286 = a5280 & i64;
assign a5288 = ~a5286 & ~a5284;
assign a5290 = a5274 & a4284;
assign a5292 = a5264 & ~a5220;
assign a5294 = ~a5292 & ~a5290;
assign a5296 = ~a5294 & ~i116;
assign a5298 = ~a5296 & ~a5288;
assign a5300 = a5294 & i116;
assign a5302 = ~a5300 & ~a5298;
assign a5304 = a5274 & a4310;
assign a5306 = a5264 & ~a5232;
assign a5308 = ~a5306 & ~a5304;
assign a5310 = ~a5308 & ~i118;
assign a5312 = ~a5310 & ~a5302;
assign a5314 = a5308 & i118;
assign a5316 = ~a5314 & ~a5312;
assign a5318 = a5274 & a3756;
assign a5320 = a5264 & ~a5244;
assign a5322 = ~a5320 & ~a5318;
assign a5324 = ~a5322 & ~i120;
assign a5326 = ~a5324 & ~a5316;
assign a5328 = a5322 & i120;
assign a5330 = ~a5328 & ~a5326;
assign a5332 = ~a5256 & a4378;
assign a5334 = a5332 & ~i122;
assign a5336 = ~a5334 & ~a5330;
assign a5338 = ~a5332 & i122;
assign a5340 = ~i120 & ~i116;
assign a5342 = ~i66 & ~i64;
assign a5344 = ~i122 & ~i118;
assign a5346 = a5344 & a5342;
assign a5348 = a5346 & a5340;
assign a5350 = i124 & i14;
assign a5352 = ~i128 & ~i126;
assign a5354 = a5352 & a5350;
assign a5356 = a5354 & ~a5348;
assign a5358 = a5356 & ~a5338;
assign a5360 = a5358 & ~a5336;
assign a5362 = a5360 & i64;
assign a5364 = ~a5362 & ~l1686;
assign a5366 = l1686 & l552;
assign a5368 = ~a5366 & ~a5364;
assign a5370 = a5360 & i116;
assign a5372 = ~a5370 & ~l1686;
assign a5374 = l1686 & l554;
assign a5376 = ~a5374 & ~a5372;
assign a5378 = a5360 & i118;
assign a5380 = ~a5378 & ~l1686;
assign a5382 = l1686 & l556;
assign a5384 = ~a5382 & ~a5380;
assign a5386 = a5360 & i120;
assign a5388 = ~a5386 & ~l1686;
assign a5390 = l1686 & l558;
assign a5392 = ~a5390 & ~a5388;
assign a5394 = l1686 & ~l560;
assign a5396 = l1686 & ~l562;
assign a5398 = l1686 & ~l564;
assign a5400 = ~a5398 & ~a2268;
assign a5402 = a5398 & a2268;
assign a5404 = ~a5402 & ~a5400;
assign a5406 = ~a5404 & ~a5396;
assign a5408 = a5404 & a5396;
assign a5410 = ~a5408 & ~a5406;
assign a5412 = ~a5410 & ~a2548;
assign a5414 = ~a5404 & a2548;
assign a5416 = ~a5414 & ~a5412;
assign a5418 = ~a5416 & ~a5394;
assign a5420 = ~a5404 & ~a2548;
assign a5422 = a5410 & a2548;
assign a5424 = ~a5422 & ~a5420;
assign a5426 = a5424 & a5394;
assign a5428 = ~a5426 & ~a5418;
assign a5430 = ~a5428 & ~a4404;
assign a5432 = ~a5416 & a4404;
assign a5434 = ~a5432 & ~a5430;
assign a5436 = ~a5434 & ~a5392;
assign a5438 = ~a5424 & ~a4404;
assign a5440 = a5428 & a4404;
assign a5442 = ~a5440 & ~a5438;
assign a5444 = a5442 & a5392;
assign a5446 = ~a5444 & ~a5436;
assign a5448 = ~a5446 & ~a2566;
assign a5450 = ~a5434 & a2566;
assign a5452 = ~a5450 & ~a5448;
assign a5454 = ~a5452 & ~a5384;
assign a5456 = ~a5442 & ~a2566;
assign a5458 = a5446 & a2566;
assign a5460 = ~a5458 & ~a5456;
assign a5462 = a5460 & a5384;
assign a5464 = ~a5462 & ~a5454;
assign a5466 = ~a5464 & ~a4428;
assign a5468 = ~a5452 & a4428;
assign a5470 = ~a5468 & ~a5466;
assign a5472 = ~a5470 & ~a5376;
assign a5474 = ~a5460 & ~a4428;
assign a5476 = a5464 & a4428;
assign a5478 = ~a5476 & ~a5474;
assign a5480 = a5478 & a5376;
assign a5482 = ~a5480 & ~a5472;
assign a5484 = ~a5482 & ~a4464;
assign a5486 = ~a5470 & a4464;
assign a5488 = ~a5486 & ~a5484;
assign a5490 = ~a5488 & ~a5368;
assign a5492 = ~a5478 & ~a4464;
assign a5494 = a5482 & a4464;
assign a5496 = ~a5494 & ~a5492;
assign a5498 = a5496 & a5368;
assign a5500 = ~a5498 & ~a5490;
assign a5502 = ~a5500 & ~a4500;
assign a5504 = ~a5488 & a4500;
assign a5506 = ~a5504 & ~a5502;
assign a5508 = a5360 & i66;
assign a5510 = ~a5508 & ~l1686;
assign a5512 = l1686 & l566;
assign a5514 = ~a5512 & ~a5510;
assign a5516 = ~a5514 & a4536;
assign a5518 = a5516 & ~a5506;
assign a5520 = ~a5496 & ~a4500;
assign a5522 = ~a5520 & ~a5516;
assign a5524 = a5500 & a4500;
assign a5526 = ~a5524 & a5522;
assign a5528 = ~a5526 & ~a5518;
assign a5530 = a5528 & l494;
assign a5532 = a5530 & ~a5198;
assign a5534 = ~a5532 & ~a5122;
assign a5536 = a1728 & ~a1704;
assign a5538 = ~a5536 & ~l1686;
assign a5540 = l1686 & l568;
assign a5542 = ~a5540 & ~a5538;
assign a5544 = ~a1738 & ~l1686;
assign a5546 = l1686 & l570;
assign a5548 = ~a5546 & ~a5544;
assign a5550 = ~a1728 & a1704;
assign a5552 = a5550 & ~l1686;
assign a5554 = l1686 & l572;
assign a5556 = ~a5554 & ~a5552;
assign a5558 = ~l586 & ~l584;
assign a5560 = a5558 & ~l582;
assign a5562 = a5560 & ~l580;
assign a5564 = a5562 & ~l578;
assign a5566 = a5564 & ~l576;
assign a5568 = a1720 & ~l1686;
assign a5570 = l1686 & l574;
assign a5572 = ~a5570 & ~a5568;
assign a5574 = a5572 & a5566;
assign a5576 = a5574 & a5556;
assign a5578 = a5576 & a5548;
assign a5580 = a5578 & a5542;
assign a5582 = ~a5580 & ~a5534;
assign a5584 = ~a5112 & ~a5016;
assign a5586 = ~a5584 & ~l494;
assign a5588 = ~a5586 & ~a5530;
assign a5590 = ~a5588 & a5580;
assign a5592 = ~a5590 & ~a5582;
assign a5594 = l1686 & ~l632;
assign a5596 = l1686 & ~l634;
assign a5598 = l1686 & ~l638;
assign a5600 = l1686 & ~l636;
assign a5602 = a2306 & ~a2292;
assign a5604 = a5602 & ~a2280;
assign a5606 = a5604 & ~a5600;
assign a5608 = a2318 & a2292;
assign a5610 = a5608 & ~a2280;
assign a5612 = a5610 & a5600;
assign a5614 = ~a5612 & ~a5606;
assign a5616 = ~a5614 & ~a2284;
assign a5618 = a5616 & ~a5598;
assign a5620 = a2300 & ~a2292;
assign a5622 = a5620 & ~a2280;
assign a5624 = ~a5622 & ~a5600;
assign a5626 = a2314 & a2292;
assign a5628 = a5626 & ~a2280;
assign a5630 = ~a5628 & a5600;
assign a5632 = ~a5630 & ~a5624;
assign a5634 = a5632 & ~a2284;
assign a5636 = a5634 & a5598;
assign a5638 = ~a5636 & ~a5618;
assign a5640 = ~a5638 & ~a5596;
assign a5642 = a5620 & a2280;
assign a5644 = ~a5642 & ~a5600;
assign a5646 = a5626 & a2280;
assign a5648 = ~a5646 & a5600;
assign a5650 = ~a5648 & ~a5644;
assign a5652 = a5650 & a2284;
assign a5654 = ~a5652 & a5598;
assign a5656 = a5602 & a2280;
assign a5658 = ~a5656 & ~a5600;
assign a5660 = a5608 & a2280;
assign a5662 = ~a5660 & a5600;
assign a5664 = ~a5662 & ~a5658;
assign a5666 = a5664 & a2284;
assign a5668 = ~a5666 & ~a5598;
assign a5670 = ~a5668 & ~a5654;
assign a5672 = a5670 & a5596;
assign a5674 = ~a5672 & ~a5640;
assign a5676 = ~a5674 & a2270;
assign a5678 = a5676 & a2274;
assign a5680 = ~a5678 & ~a5594;
assign a5682 = ~a5616 & a5598;
assign a5684 = ~a5682 & ~a5668;
assign a5686 = ~a5684 & ~a5596;
assign a5688 = ~a5610 & ~a5600;
assign a5690 = ~a5622 & a5600;
assign a5692 = ~a5690 & ~a5688;
assign a5694 = a5692 & ~a2284;
assign a5696 = ~a5694 & a5596;
assign a5698 = ~a5696 & ~a5686;
assign a5700 = a5698 & ~a2270;
assign a5702 = a5700 & ~a2274;
assign a5704 = ~a5702 & a5594;
assign a5706 = ~a5704 & ~a5680;
assign a5708 = ~a5706 & ~l506;
assign a5710 = a5604 & ~a2336;
assign a5712 = a5610 & a2336;
assign a5714 = ~a5712 & ~a5710;
assign a5716 = ~a5714 & ~a2284;
assign a5718 = a5716 & ~a2334;
assign a5720 = ~a5622 & ~a2336;
assign a5722 = ~a5628 & a2336;
assign a5724 = ~a5722 & ~a5720;
assign a5726 = a5724 & ~a2284;
assign a5728 = a5726 & a2334;
assign a5730 = ~a5728 & ~a5718;
assign a5732 = ~a5730 & ~a2332;
assign a5734 = ~a5656 & ~a2336;
assign a5736 = ~a5660 & a2336;
assign a5738 = ~a5736 & ~a5734;
assign a5740 = a5738 & a2284;
assign a5742 = ~a5740 & ~a2334;
assign a5744 = ~a5742 & a2332;
assign a5746 = ~a5642 & ~a2336;
assign a5748 = ~a5646 & a2336;
assign a5750 = ~a5748 & ~a5746;
assign a5752 = a5750 & a2284;
assign a5754 = ~a5752 & a2334;
assign a5756 = ~a5754 & a5744;
assign a5758 = ~a5756 & ~a5732;
assign a5760 = ~a5758 & a2270;
assign a5762 = a5760 & a2274;
assign a5764 = ~a5762 & ~a2330;
assign a5766 = ~a5716 & a2334;
assign a5768 = ~a5766 & ~a5742;
assign a5770 = ~a5768 & ~a2332;
assign a5772 = ~a5610 & ~a2336;
assign a5774 = ~a5622 & a2336;
assign a5776 = ~a5774 & ~a5772;
assign a5778 = a5776 & ~a2284;
assign a5780 = ~a5778 & a2332;
assign a5782 = ~a5780 & ~a5770;
assign a5784 = a5782 & ~a2270;
assign a5786 = a5784 & ~a2274;
assign a5788 = ~a5786 & a2330;
assign a5790 = ~a5788 & ~a5764;
assign a5792 = ~a5790 & l506;
assign a5794 = a5792 & ~l508;
assign a5796 = ~a5794 & ~a2424;
assign a5798 = a5796 & ~a5708;
assign a5800 = ~a5798 & ~l512;
assign a5802 = ~a5800 & ~a2512;
assign a5804 = a5604 & ~a2436;
assign a5806 = a5610 & a2436;
assign a5808 = ~a5806 & ~a5804;
assign a5810 = ~a5808 & ~a2284;
assign a5812 = a5810 & ~a2434;
assign a5814 = ~a5622 & ~a2436;
assign a5816 = ~a5628 & a2436;
assign a5818 = ~a5816 & ~a5814;
assign a5820 = a5818 & ~a2284;
assign a5822 = a5820 & a2434;
assign a5824 = ~a5822 & ~a5812;
assign a5826 = ~a5824 & ~a2432;
assign a5828 = ~a5642 & ~a2436;
assign a5830 = ~a5646 & a2436;
assign a5832 = ~a5830 & ~a5828;
assign a5834 = a5832 & a2284;
assign a5836 = ~a5834 & a2434;
assign a5838 = ~a5656 & ~a2436;
assign a5840 = ~a5660 & a2436;
assign a5842 = ~a5840 & ~a5838;
assign a5844 = a5842 & a2284;
assign a5846 = ~a5844 & ~a2434;
assign a5848 = ~a5846 & ~a5836;
assign a5850 = a5848 & a2432;
assign a5852 = ~a5850 & ~a5826;
assign a5854 = ~a5852 & a2270;
assign a5856 = a5854 & a2274;
assign a5858 = ~a5856 & ~a2430;
assign a5860 = ~a5810 & a2434;
assign a5862 = ~a5860 & ~a5846;
assign a5864 = ~a5862 & ~a2432;
assign a5866 = ~a5610 & ~a2436;
assign a5868 = ~a5622 & a2436;
assign a5870 = ~a5868 & ~a5866;
assign a5872 = a5870 & ~a2284;
assign a5874 = ~a5872 & a2432;
assign a5876 = ~a5874 & ~a5864;
assign a5878 = a5876 & ~a2270;
assign a5880 = a5878 & ~a2274;
assign a5882 = ~a5880 & a2430;
assign a5884 = ~a5882 & ~a5858;
assign a5886 = ~a5884 & ~l506;
assign a5888 = ~a5886 & a5796;
assign a5890 = ~a5888 & l512;
assign a5892 = a5890 & ~l510;
assign a5894 = ~a5892 & a5802;
assign a5896 = ~a5894 & l516;
assign a5898 = ~a2514 & ~l516;
assign a5900 = ~a5898 & ~a5896;
assign a5902 = ~a5900 & l514;
assign a5904 = ~a2514 & ~l514;
assign a5906 = ~a5904 & ~a5902;
assign a5908 = ~a5906 & a2268;
assign a5910 = ~a5908 & ~a2266;
assign a5912 = ~a5906 & ~a2268;
assign a5914 = ~a5912 & a2266;
assign a5916 = ~a5914 & ~a5910;
assign a5918 = ~a5916 & a2528;
assign a5920 = a5912 & ~a2266;
assign a5922 = a5908 & a2266;
assign a5924 = ~a5922 & ~a5920;
assign a5926 = a5924 & ~a2528;
assign a5928 = ~a5926 & ~a5918;
assign a5930 = ~a5928 & a2544;
assign a5932 = ~a5924 & ~a2548;
assign a5934 = a5916 & a2548;
assign a5936 = ~a5934 & ~a5932;
assign a5938 = ~a5936 & ~a2526;
assign a5940 = ~a5924 & a2526;
assign a5942 = ~a5940 & ~a5938;
assign a5944 = a5942 & ~a2544;
assign a5946 = ~a5944 & ~a5930;
assign a5948 = ~a5946 & a4400;
assign a5950 = ~a5942 & ~a4404;
assign a5952 = ~a5916 & ~a2526;
assign a5954 = a5936 & a2526;
assign a5956 = ~a5954 & ~a5952;
assign a5958 = a5956 & a4404;
assign a5960 = ~a5958 & ~a5950;
assign a5962 = ~a5960 & ~a2542;
assign a5964 = ~a5942 & a2542;
assign a5966 = ~a5964 & ~a5962;
assign a5968 = a5966 & ~a4400;
assign a5970 = ~a5968 & ~a5948;
assign a5972 = ~a5970 & a4438;
assign a5974 = ~a5966 & ~a2566;
assign a5976 = ~a5956 & ~a2542;
assign a5978 = a5960 & a2542;
assign a5980 = ~a5978 & ~a5976;
assign a5982 = a5980 & a2566;
assign a5984 = ~a5982 & ~a5974;
assign a5986 = ~a5984 & ~a4398;
assign a5988 = ~a5966 & a4398;
assign a5990 = ~a5988 & ~a5986;
assign a5992 = a5990 & ~a4438;
assign a5994 = ~a5992 & ~a5972;
assign a5996 = ~a5994 & a4474;
assign a5998 = ~a5990 & ~a4428;
assign a6000 = ~a5980 & ~a4398;
assign a6002 = a5984 & a4398;
assign a6004 = ~a6002 & ~a6000;
assign a6006 = a6004 & a4428;
assign a6008 = ~a6006 & ~a5998;
assign a6010 = ~a6008 & ~a4436;
assign a6012 = ~a5990 & a4436;
assign a6014 = ~a6012 & ~a6010;
assign a6016 = a6014 & ~a4474;
assign a6018 = ~a6016 & ~a5996;
assign a6020 = ~a6018 & a4510;
assign a6022 = ~a6014 & ~a4464;
assign a6024 = ~a6004 & ~a4436;
assign a6026 = a6008 & a4436;
assign a6028 = ~a6026 & ~a6024;
assign a6030 = a6028 & a4464;
assign a6032 = ~a6030 & ~a6022;
assign a6034 = ~a6032 & ~a4472;
assign a6036 = ~a6014 & a4472;
assign a6038 = ~a6036 & ~a6034;
assign a6040 = a6038 & ~a4510;
assign a6042 = ~a6040 & ~a6020;
assign a6044 = ~a6042 & a4546;
assign a6046 = ~a6028 & ~a4472;
assign a6048 = a6032 & a4472;
assign a6050 = ~a6048 & ~a6046;
assign a6052 = ~a6050 & a4556;
assign a6054 = a6038 & ~a4556;
assign a6056 = ~a6054 & ~a6052;
assign a6058 = ~a6056 & ~a4546;
assign a6060 = ~a6058 & ~a6044;
assign a6062 = a6060 & a1690;
assign a6064 = ~a6062 & ~a5118;
assign a6066 = ~a6064 & ~l494;
assign a6068 = ~a6066 & ~a5532;
assign a6070 = ~a6068 & ~a5580;
assign a6072 = ~a6070 & ~a5590;
assign a6076 = a6074 & a5592;
assign a6078 = ~a6076 & i154;
assign a6080 = ~a5600 & a2338;
assign a6082 = a5600 & a2342;
assign a6084 = ~a6082 & ~a6080;
assign a6086 = ~a6084 & ~a5598;
assign a6088 = ~a5600 & ~a2350;
assign a6090 = a5600 & ~a2354;
assign a6092 = ~a6090 & ~a6088;
assign a6094 = a6092 & a5598;
assign a6096 = ~a6094 & ~a6086;
assign a6098 = ~a6096 & ~a5596;
assign a6100 = ~a5600 & ~a2380;
assign a6102 = a5600 & ~a2384;
assign a6104 = ~a6102 & ~a6100;
assign a6106 = ~a6104 & a5598;
assign a6108 = ~a5600 & ~a2366;
assign a6110 = a5600 & ~a2370;
assign a6112 = ~a6110 & ~a6108;
assign a6114 = ~a6112 & ~a5598;
assign a6116 = ~a6114 & ~a6106;
assign a6118 = a6116 & a5596;
assign a6120 = ~a6118 & ~a6098;
assign a6122 = ~a6120 & a2270;
assign a6124 = ~a6122 & ~a5594;
assign a6126 = a6084 & a5598;
assign a6128 = ~a6126 & ~a6114;
assign a6130 = ~a6128 & ~a5596;
assign a6132 = ~a5600 & ~a2342;
assign a6134 = a5600 & ~a2350;
assign a6136 = ~a6134 & ~a6132;
assign a6138 = ~a6136 & a5596;
assign a6140 = ~a6138 & ~a6130;
assign a6142 = a6140 & ~a2270;
assign a6144 = ~a6142 & a5594;
assign a6146 = ~a6144 & ~a6124;
assign a6148 = ~a6146 & ~l506;
assign a6150 = ~a6148 & ~a2422;
assign a6152 = ~a6150 & ~l512;
assign a6154 = ~a6152 & ~a2510;
assign a6156 = ~a6154 & l516;
assign a6158 = ~a6156 & ~a5898;
assign a6160 = ~a6158 & l514;
assign a6162 = ~a6160 & ~a5904;
assign a6164 = ~a6162 & a2268;
assign a6166 = ~a6164 & ~a2266;
assign a6168 = ~a6162 & ~a2268;
assign a6170 = ~a6168 & a2266;
assign a6172 = ~a6170 & ~a6166;
assign a6174 = ~a6172 & a2528;
assign a6176 = a6168 & ~a2266;
assign a6178 = a6164 & a2266;
assign a6180 = ~a6178 & ~a6176;
assign a6182 = a6180 & ~a2528;
assign a6184 = ~a6182 & ~a6174;
assign a6186 = ~a6184 & a2544;
assign a6188 = ~a6180 & ~a2548;
assign a6190 = a6172 & a2548;
assign a6192 = ~a6190 & ~a6188;
assign a6194 = ~a6192 & ~a2526;
assign a6196 = ~a6180 & a2526;
assign a6198 = ~a6196 & ~a6194;
assign a6200 = a6198 & ~a2544;
assign a6202 = ~a6200 & ~a6186;
assign a6204 = ~a6202 & a4400;
assign a6206 = ~a6198 & ~a4404;
assign a6208 = ~a6172 & ~a2526;
assign a6210 = a6192 & a2526;
assign a6212 = ~a6210 & ~a6208;
assign a6214 = a6212 & a4404;
assign a6216 = ~a6214 & ~a6206;
assign a6218 = ~a6216 & ~a2542;
assign a6220 = ~a6198 & a2542;
assign a6222 = ~a6220 & ~a6218;
assign a6224 = a6222 & ~a4400;
assign a6226 = ~a6224 & ~a6204;
assign a6228 = ~a6226 & a4438;
assign a6230 = ~a6222 & ~a2566;
assign a6232 = ~a6212 & ~a2542;
assign a6234 = a6216 & a2542;
assign a6236 = ~a6234 & ~a6232;
assign a6238 = a6236 & a2566;
assign a6240 = ~a6238 & ~a6230;
assign a6242 = ~a6240 & ~a4398;
assign a6244 = ~a6222 & a4398;
assign a6246 = ~a6244 & ~a6242;
assign a6248 = a6246 & ~a4438;
assign a6250 = ~a6248 & ~a6228;
assign a6252 = ~a6250 & a4474;
assign a6254 = ~a6246 & ~a4428;
assign a6256 = ~a6236 & ~a4398;
assign a6258 = a6240 & a4398;
assign a6260 = ~a6258 & ~a6256;
assign a6262 = a6260 & a4428;
assign a6264 = ~a6262 & ~a6254;
assign a6266 = ~a6264 & ~a4436;
assign a6268 = ~a6246 & a4436;
assign a6270 = ~a6268 & ~a6266;
assign a6272 = a6270 & ~a4474;
assign a6274 = ~a6272 & ~a6252;
assign a6276 = ~a6274 & a4510;
assign a6278 = ~a6270 & ~a4464;
assign a6280 = ~a6260 & ~a4436;
assign a6282 = a6264 & a4436;
assign a6284 = ~a6282 & ~a6280;
assign a6286 = a6284 & a4464;
assign a6288 = ~a6286 & ~a6278;
assign a6290 = ~a6288 & ~a4472;
assign a6292 = ~a6270 & a4472;
assign a6294 = ~a6292 & ~a6290;
assign a6296 = a6294 & ~a4510;
assign a6298 = ~a6296 & ~a6276;
assign a6300 = ~a6298 & a4546;
assign a6302 = ~a6284 & ~a4472;
assign a6304 = a6288 & a4472;
assign a6306 = ~a6304 & ~a6302;
assign a6308 = ~a6306 & a4556;
assign a6310 = a6294 & ~a4556;
assign a6312 = ~a6310 & ~a6308;
assign a6314 = ~a6312 & ~a4546;
assign a6316 = ~a6314 & ~a6300;
assign a6318 = a6316 & a1690;
assign a6320 = ~a6318 & ~a5118;
assign a6322 = ~a6320 & ~l494;
assign a6324 = ~a6322 & ~a5532;
assign a6326 = ~a6324 & ~a5580;
assign a6328 = ~a6326 & ~a5590;
assign a6330 = ~a6076 & i2;
assign a6332 = ~a6330 & a6074;
assign a6334 = a6332 & a6328;
assign a6336 = ~a6334 & ~a6078;
assign a6338 = ~a6330 & l516;
assign a6340 = a6338 & a6336;
assign a6342 = a6340 & l514;
assign a6344 = ~a6342 & ~a2264;
assign a6348 = a6346 & a2260;
assign a6350 = a2334 & l506;
assign a6352 = l512 & ~l506;
assign a6354 = a6352 & a2434;
assign a6356 = ~a6354 & ~a6350;
assign a6358 = ~l512 & ~l506;
assign a6360 = a6358 & a5598;
assign a6364 = a2336 & l506;
assign a6366 = a6352 & a2436;
assign a6368 = ~a6366 & ~a6364;
assign a6370 = a6358 & a5600;
assign a6374 = a6372 & ~a6362;
assign a6376 = a2332 & l506;
assign a6378 = a6352 & a2432;
assign a6380 = ~a6378 & ~a6376;
assign a6382 = a6358 & a5596;
assign a6386 = a2330 & l506;
assign a6388 = a6352 & a2430;
assign a6390 = ~a6388 & ~a6386;
assign a6392 = a6358 & a5594;
assign a6396 = ~a6394 & a6384;
assign a6398 = a6396 & a6374;
assign a6400 = l1686 & ~l656;
assign a6402 = a6400 & l506;
assign a6404 = l1686 & ~l654;
assign a6406 = a6404 & a6352;
assign a6408 = ~a6406 & ~a6402;
assign a6410 = l1686 & ~l652;
assign a6412 = a6410 & a6358;
assign a6414 = ~a6412 & a6408;
assign a6416 = a6414 & a6398;
assign a6418 = ~a6414 & ~a6398;
assign a6420 = ~a6418 & ~a6416;
assign a6422 = ~a6420 & ~a6346;
assign a6426 = ~a6424 & a1690;
assign a6428 = ~a6426 & ~a2258;
assign a6430 = ~a6428 & ~l494;
assign a6432 = l1686 & ~l650;
assign a6434 = a5128 & a5124;
assign a6436 = a6434 & ~a5130;
assign a6438 = a6436 & ~a5126;
assign a6440 = ~a6438 & a6432;
assign a6442 = a6438 & ~a6432;
assign a6444 = ~a6442 & ~a6440;
assign a6446 = ~a6444 & l494;
assign a6450 = ~a6448 & ~a1688;
assign a6452 = a6448 & a1688;
assign a6454 = ~a6452 & ~a6450;
assign a6456 = ~a2248 & a1750;
assign a6458 = ~a6456 & ~a1694;
assign a6460 = ~a6458 & ~a2250;
assign a6462 = a6460 & ~a1690;
assign a6464 = a6346 & a2294;
assign a6466 = a6394 & ~a6362;
assign a6468 = ~a6394 & ~a6384;
assign a6470 = a6468 & ~a6372;
assign a6472 = ~a6470 & ~a6466;
assign a6474 = ~a6472 & ~a6346;
assign a6478 = ~a6476 & a1690;
assign a6480 = ~a6478 & ~a6462;
assign a6482 = ~a6480 & ~l494;
assign a6484 = a5128 & l500;
assign a6486 = a5126 & a5124;
assign a6488 = a6486 & a5130;
assign a6490 = ~a6488 & ~a6484;
assign a6492 = ~a6490 & l494;
assign a6496 = a6494 & a2296;
assign a6498 = ~a6496 & ~a6454;
assign a6500 = a2246 & ~a1736;
assign a6502 = ~a2246 & a1736;
assign a6504 = ~a6502 & ~a6500;
assign a6506 = a6504 & ~a1690;
assign a6508 = a6346 & a2274;
assign a6510 = a6394 & ~a6346;
assign a6514 = ~a6512 & a1690;
assign a6516 = ~a6514 & ~a6506;
assign a6518 = ~a6516 & ~l494;
assign a6520 = ~a5124 & l494;
assign a6524 = ~a6522 & ~a2270;
assign a6526 = ~a1758 & ~a1748;
assign a6528 = ~a6526 & ~a2248;
assign a6530 = ~a2248 & a1736;
assign a6532 = ~a6530 & ~a1746;
assign a6534 = ~a6532 & ~a6528;
assign a6536 = a6534 & ~a1690;
assign a6538 = a6346 & a2284;
assign a6540 = a6394 & ~a6384;
assign a6542 = a6396 & a6362;
assign a6544 = ~a6542 & ~a6540;
assign a6546 = ~a6544 & ~a6346;
assign a6550 = ~a6548 & a1690;
assign a6552 = ~a6550 & ~a6536;
assign a6554 = ~a6552 & ~l494;
assign a6556 = a5126 & l500;
assign a6558 = ~a5128 & ~a5126;
assign a6560 = a6558 & a5124;
assign a6562 = ~a6560 & ~a6556;
assign a6564 = ~a6562 & l494;
assign a6568 = ~a6566 & ~a2280;
assign a6570 = ~a6568 & ~a6524;
assign a6572 = a6566 & a2280;
assign a6574 = ~a6572 & ~a6570;
assign a6576 = ~a2248 & a1748;
assign a6578 = ~a6576 & ~a1726;
assign a6580 = ~a6578 & ~a6456;
assign a6582 = a6580 & ~a1690;
assign a6584 = a6346 & a2292;
assign a6586 = ~a6468 & a6372;
assign a6588 = ~a6586 & ~a6470;
assign a6590 = a6588 & ~a6346;
assign a6594 = ~a6592 & a1690;
assign a6596 = ~a6594 & ~a6582;
assign a6598 = ~a6596 & ~l494;
assign a6600 = ~a6486 & a5130;
assign a6602 = a6486 & ~a5130;
assign a6604 = ~a6602 & ~a6600;
assign a6606 = ~a6604 & l494;
assign a6610 = ~a6608 & ~a2302;
assign a6612 = ~a6610 & ~a6574;
assign a6614 = a6608 & a2302;
assign a6616 = ~a6614 & ~a6612;
assign a6618 = ~a6494 & ~a2296;
assign a6620 = ~a6618 & ~a6616;
assign a6622 = ~a6620 & a6498;
assign a6624 = ~a6618 & a6454;
assign a6626 = a6522 & a2270;
assign a6628 = ~a6626 & ~a6572;
assign a6630 = ~a6628 & ~a6568;
assign a6632 = ~a6630 & ~a6614;
assign a6634 = ~a6632 & ~a6610;
assign a6636 = ~a6634 & ~a6496;
assign a6638 = ~a6636 & a6624;
assign a6640 = ~a6638 & ~a6622;
assign a6642 = ~l666 & ~l664;
assign a6644 = a6642 & a2296;
assign a6646 = l666 & ~l664;
assign a6648 = a2296 & l604;
assign a6650 = a2280 & a2270;
assign a6652 = a6650 & a2302;
assign a6654 = ~a6652 & ~a6648;
assign a6656 = ~a6654 & a6646;
assign a6658 = ~a6656 & ~a6644;
assign a6660 = ~a6490 & l664;
assign a6664 = ~a1696 & i204;
assign a6666 = ~a5360 & ~a4384;
assign a6668 = a6666 & a6664;
assign a6670 = a6668 & ~l1686;
assign a6672 = l1686 & l940;
assign a6674 = ~a6672 & ~a6670;
assign a6676 = a1698 & ~l1686;
assign a6678 = l1686 & l942;
assign a6680 = ~a6678 & ~a6676;
assign a6684 = l1686 & ~l1650;
assign a6686 = l1686 & ~l1648;
assign a6688 = a6686 & ~a6604;
assign a6692 = l1686 & ~l1656;
assign a6694 = a6686 & ~a6562;
assign a6698 = l1686 & ~l1654;
assign a6700 = a6686 & l500;
assign a6704 = l1686 & ~l1652;
assign a6706 = a6686 & ~a6490;
assign a6710 = l1686 & ~l700;
assign a6714 = l1686 & ~l722;
assign a6716 = a6714 & l562;
assign a6718 = a5396 & l722;
assign a6720 = l1686 & ~l720;
assign a6722 = a6720 & l560;
assign a6724 = a5394 & l720;
assign a6726 = l1686 & ~l718;
assign a6728 = a6726 & ~a5392;
assign a6730 = ~a6726 & a5392;
assign a6732 = a1716 & ~a1704;
assign a6734 = i176 & i172;
assign a6736 = a6734 & i180;
assign a6738 = a6736 & ~a6732;
assign a6740 = ~a6738 & ~l1686;
assign a6742 = l1686 & l716;
assign a6744 = ~a6742 & ~a6740;
assign a6746 = a6744 & ~a5384;
assign a6748 = ~a6744 & a5384;
assign a6750 = a6732 & i62;
assign a6752 = ~a1912 & i62;
assign a6754 = i174 & ~i62;
assign a6756 = ~a6754 & ~a6752;
assign a6758 = a6756 & ~i176;
assign a6760 = ~a1814 & i62;
assign a6762 = i170 & ~i62;
assign a6764 = ~a6762 & ~a6760;
assign a6766 = ~a6764 & i172;
assign a6768 = ~a6756 & i176;
assign a6770 = ~a6768 & ~a6766;
assign a6772 = ~a6770 & ~a6758;
assign a6774 = ~a1994 & i62;
assign a6776 = i178 & ~i62;
assign a6778 = ~a6776 & ~a6774;
assign a6780 = ~a6778 & ~i180;
assign a6782 = a6778 & i180;
assign a6784 = ~a6782 & ~a6780;
assign a6786 = ~a6784 & ~a6772;
assign a6788 = a6784 & a6772;
assign a6790 = ~a6788 & ~a6786;
assign a6792 = ~a6790 & a6750;
assign a6794 = ~a6734 & ~i180;
assign a6796 = ~a6794 & ~a6736;
assign a6798 = a6796 & ~a6732;
assign a6800 = ~a6798 & ~a6792;
assign a6802 = a6800 & ~l1686;
assign a6804 = l1686 & l714;
assign a6806 = ~a6804 & ~a6802;
assign a6808 = a6806 & ~a5376;
assign a6810 = ~a6806 & a5376;
assign a6812 = a6770 & ~a6758;
assign a6814 = ~a6768 & ~a6758;
assign a6816 = ~a6814 & a6766;
assign a6818 = ~a6816 & ~a6812;
assign a6820 = ~a6818 & a6750;
assign a6822 = ~i176 & ~i172;
assign a6824 = ~a6822 & ~a6734;
assign a6826 = a6824 & ~a6732;
assign a6828 = ~a6826 & ~a6820;
assign a6830 = a6828 & ~l1686;
assign a6832 = l1686 & l712;
assign a6834 = ~a6832 & ~a6830;
assign a6836 = a6834 & ~a5368;
assign a6838 = ~a6834 & a5368;
assign a6840 = a6764 & ~i172;
assign a6842 = ~a6840 & a6750;
assign a6844 = ~a6732 & ~i172;
assign a6846 = ~a6844 & ~a6842;
assign a6848 = a6846 & ~l1686;
assign a6850 = l1686 & l710;
assign a6852 = ~a6850 & ~a6848;
assign a6854 = ~a6852 & a5514;
assign a6856 = ~a6854 & ~a6838;
assign a6858 = ~a6856 & ~a6836;
assign a6860 = ~a6858 & ~a6810;
assign a6862 = ~a6860 & ~a6808;
assign a6864 = ~a6862 & ~a6748;
assign a6866 = ~a6864 & ~a6746;
assign a6868 = ~a6866 & ~a6730;
assign a6870 = ~a6868 & ~a6728;
assign a6872 = ~a6870 & ~a6724;
assign a6874 = ~a6872 & ~a6722;
assign a6876 = ~a6874 & ~a6718;
assign a6878 = ~a6876 & ~a6716;
assign a6880 = a5398 & l708;
assign a6882 = l1686 & ~l708;
assign a6884 = a6882 & l564;
assign a6886 = ~a6884 & ~a6880;
assign a6888 = ~a6886 & ~a6878;
assign a6890 = a6886 & a6878;
assign a6892 = ~a6890 & ~a6888;
assign a6894 = ~a6732 & i168;
assign a6896 = a6894 & ~l1686;
assign a6898 = l1686 & l704;
assign a6900 = ~a6898 & ~a6896;
assign a6902 = l1686 & ~l706;
assign a6904 = a6902 & ~a6900;
assign a6906 = a6904 & ~l494;
assign a6908 = a6906 & ~a6892;
assign a6910 = ~a6908 & a4500;
assign a6912 = ~a6906 & i192;
assign a6914 = a6906 & a6834;
assign a6916 = ~a6914 & ~a6912;
assign a6918 = ~a6916 & a6908;
assign a6922 = a4672 & a2246;
assign a6924 = ~a4962 & ~a4500;
assign a6926 = ~a4980 & ~a4964;
assign a6928 = ~a6926 & a4500;
assign a6930 = ~a6928 & ~a6924;
assign a6932 = ~a6930 & ~a4644;
assign a6934 = ~a2246 & ~l494;
assign a6936 = a6074 & ~a5580;
assign a6938 = a6936 & a6934;
assign a6940 = a6938 & ~a1690;
assign a6942 = ~a4988 & ~a4536;
assign a6944 = ~a5006 & ~a4990;
assign a6946 = ~a6944 & a4536;
assign a6948 = ~a6946 & ~a6942;
assign a6950 = a6934 & a5580;
assign a6952 = a6950 & a6074;
assign a6954 = a6952 & a6948;
assign a6956 = ~a6954 & i482;
assign a6958 = ~a6948 & ~a4644;
assign a6960 = ~a6958 & a6940;
assign a6962 = ~a6960 & a6956;
assign a6964 = ~a6944 & ~a4536;
assign a6966 = ~a5004 & a4536;
assign a6968 = ~a6966 & ~a6964;
assign a6970 = a6968 & a6952;
assign a6972 = ~a6968 & ~a4644;
assign a6974 = ~a6972 & a6940;
assign a6976 = ~a6974 & ~a6970;
assign a6978 = a6976 & ~a6962;
assign a6980 = a6978 & a6940;
assign a6982 = a6980 & ~a4536;
assign a6984 = ~a6978 & a6940;
assign a6986 = a6984 & a4536;
assign a6988 = ~a6986 & ~a6982;
assign a6990 = ~a6988 & a4656;
assign a6992 = a6984 & ~a4536;
assign a6994 = ~a6992 & ~a6990;
assign a6996 = ~a6994 & ~a6932;
assign a6998 = ~a6996 & i484;
assign a7000 = a6980 & a4536;
assign a7002 = ~a6988 & ~a4656;
assign a7004 = ~a7002 & ~a7000;
assign a7006 = ~a6926 & ~a4500;
assign a7008 = ~a4978 & a4500;
assign a7010 = ~a7008 & ~a7006;
assign a7012 = ~a7010 & ~a4644;
assign a7014 = ~a7012 & ~a7004;
assign a7016 = ~a7014 & a6998;
assign a7018 = a6978 & a6952;
assign a7020 = a7018 & a4536;
assign a7022 = a7018 & ~a4536;
assign a7024 = ~a6978 & a6952;
assign a7026 = a7024 & a4536;
assign a7028 = ~a7026 & ~a7022;
assign a7030 = ~a7028 & ~a4656;
assign a7032 = ~a7030 & ~a7020;
assign a7034 = ~a7032 & a7010;
assign a7036 = ~a7028 & a4656;
assign a7038 = a7024 & ~a4536;
assign a7040 = ~a7038 & ~a7036;
assign a7042 = ~a7040 & a6930;
assign a7044 = ~a7042 & ~a7034;
assign a7046 = a7044 & a7016;
assign a7048 = ~a4850 & ~a4464;
assign a7050 = ~a4832 & ~a4428;
assign a7052 = ~a4814 & ~a2566;
assign a7054 = ~a7052 & ~a5036;
assign a7056 = ~a7054 & ~a4722;
assign a7058 = ~a4890 & a4722;
assign a7060 = ~a7058 & ~a7056;
assign a7062 = ~a7060 & a4428;
assign a7064 = ~a7062 & ~a7050;
assign a7066 = ~a7064 & ~a4706;
assign a7068 = ~a4904 & a4706;
assign a7070 = ~a7068 & ~a7066;
assign a7072 = ~a7070 & a4464;
assign a7074 = ~a7072 & ~a7048;
assign a7076 = ~a7074 & ~a4690;
assign a7078 = ~a4972 & a4690;
assign a7080 = ~a7078 & ~a7076;
assign a7082 = ~a7080 & a4674;
assign a7084 = ~a4978 & ~a4674;
assign a7086 = ~a7084 & ~a7082;
assign a7088 = ~a7086 & ~a4644;
assign a7090 = ~a7088 & ~a7004;
assign a7092 = ~a7012 & ~a6994;
assign a7094 = ~a7092 & ~a7090;
assign a7096 = ~a7040 & a7010;
assign a7098 = ~a7096 & a7094;
assign a7100 = a7086 & ~a7032;
assign a7102 = ~a7100 & a7098;
assign a7104 = a7102 & ~a7046;
assign a7106 = a7104 & ~a4672;
assign a7108 = ~a7104 & a4672;
assign a7110 = ~a7108 & ~a7106;
assign a7112 = ~a6978 & a4656;
assign a7114 = a7112 & ~a7110;
assign a7116 = ~a7112 & a7110;
assign a7118 = ~a7116 & ~a7114;
assign a7120 = a6978 & ~a4656;
assign a7122 = ~a7120 & ~a7112;
assign a7124 = ~a7122 & a7118;
assign a7126 = a7122 & ~a7118;
assign a7128 = ~a7126 & ~a7124;
assign a7130 = a7128 & ~a2246;
assign a7132 = ~a7130 & ~a6922;
assign a7134 = ~a5580 & a1690;
assign a7136 = ~a7134 & ~a7132;
assign a7138 = ~a4544 & ~a4508;
assign a7140 = a4544 & a4508;
assign a7142 = ~a7140 & ~a7138;
assign a7144 = a7142 & a7134;
assign a7146 = ~a7144 & ~a7136;
assign a7148 = ~a7146 & ~l494;
assign a7150 = a5368 & l494;
assign a7154 = a4690 & a2246;
assign a7156 = ~a7072 & ~a4970;
assign a7158 = ~a7156 & ~a4690;
assign a7160 = ~a4914 & a4690;
assign a7162 = ~a7160 & ~a7158;
assign a7164 = ~a7162 & ~a4644;
assign a7166 = a7104 & ~a7004;
assign a7168 = a7166 & a4674;
assign a7170 = a7168 & ~a7164;
assign a7172 = ~a7170 & i486;
assign a7174 = a7104 & ~a7032;
assign a7176 = a7174 & a4674;
assign a7178 = a7176 & a7162;
assign a7180 = ~a7178 & a7172;
assign a7182 = ~a4914 & ~a4690;
assign a7184 = ~a4954 & ~a4916;
assign a7186 = ~a7184 & a4690;
assign a7188 = ~a7186 & ~a7182;
assign a7190 = a7174 & ~a4674;
assign a7192 = ~a7104 & ~a7032;
assign a7194 = a7104 & ~a7040;
assign a7196 = ~a7194 & ~a7192;
assign a7198 = ~a7196 & a4500;
assign a7200 = ~a7198 & ~a7190;
assign a7202 = ~a7196 & ~a4500;
assign a7204 = ~a7104 & ~a7040;
assign a7206 = a7204 & a4500;
assign a7208 = ~a7206 & ~a7202;
assign a7210 = ~a7208 & ~a4672;
assign a7212 = ~a7210 & a7200;
assign a7214 = ~a7212 & a7188;
assign a7216 = ~a7214 & a7180;
assign a7218 = ~a7184 & ~a4690;
assign a7220 = ~a4952 & a4690;
assign a7222 = ~a7220 & ~a7218;
assign a7224 = ~a7222 & ~a4644;
assign a7226 = ~a7104 & ~a7004;
assign a7228 = a7104 & ~a6994;
assign a7230 = ~a7228 & ~a7226;
assign a7232 = ~a7230 & ~a4500;
assign a7234 = ~a7104 & ~a6994;
assign a7236 = a7234 & a4500;
assign a7238 = ~a7236 & ~a7232;
assign a7240 = ~a7238 & a4672;
assign a7242 = a7234 & ~a4500;
assign a7244 = ~a7242 & ~a7240;
assign a7246 = ~a7244 & ~a7224;
assign a7248 = ~a7246 & a7216;
assign a7250 = ~a7208 & a4672;
assign a7252 = a7204 & ~a4500;
assign a7254 = ~a7252 & ~a7250;
assign a7256 = ~a7254 & a7222;
assign a7258 = a7166 & ~a4674;
assign a7260 = ~a7230 & a4500;
assign a7262 = ~a7260 & ~a7258;
assign a7264 = ~a7238 & ~a4672;
assign a7266 = ~a7264 & a7262;
assign a7268 = ~a7188 & ~a4644;
assign a7270 = ~a7268 & ~a7266;
assign a7272 = ~a7270 & ~a7256;
assign a7274 = a7272 & a7248;
assign a7276 = ~a7266 & ~a7164;
assign a7278 = ~a7268 & ~a7244;
assign a7280 = ~a7278 & ~a7276;
assign a7282 = ~a7070 & ~a4690;
assign a7284 = ~a7156 & a4690;
assign a7286 = ~a7284 & ~a7282;
assign a7288 = ~a7286 & ~a4644;
assign a7290 = ~a7288 & a7168;
assign a7292 = ~a7290 & a7280;
assign a7294 = ~a7254 & a7188;
assign a7296 = ~a7294 & a7292;
assign a7298 = ~a7212 & a7162;
assign a7300 = ~a7298 & a7296;
assign a7302 = a7286 & a7176;
assign a7304 = ~a7302 & a7300;
assign a7306 = a7304 & ~a7274;
assign a7308 = ~a7306 & a4690;
assign a7310 = a7306 & ~a4690;
assign a7312 = ~a7310 & ~a7308;
assign a7314 = ~a7112 & ~a7108;
assign a7316 = ~a7314 & ~a7106;
assign a7318 = a7316 & ~a7312;
assign a7320 = ~a7316 & ~a7308;
assign a7322 = a7320 & ~a7310;
assign a7324 = ~a7322 & ~a7318;
assign a7326 = a7324 & ~a7126;
assign a7328 = ~a7324 & a7126;
assign a7330 = ~a7328 & ~a7326;
assign a7332 = a7330 & ~a2246;
assign a7334 = ~a7332 & ~a7154;
assign a7336 = ~a7334 & ~a7134;
assign a7338 = ~a7140 & ~a4472;
assign a7340 = a7140 & a4472;
assign a7342 = ~a7340 & ~a7338;
assign a7344 = a7342 & a7134;
assign a7346 = ~a7344 & ~a7336;
assign a7348 = ~a7346 & ~l494;
assign a7350 = a5376 & l494;
assign a7354 = a4706 & a2246;
assign a7356 = ~a7062 & ~a4902;
assign a7358 = ~a7356 & ~a4706;
assign a7360 = ~a4900 & a4706;
assign a7362 = ~a7360 & ~a7358;
assign a7364 = a7306 & a7176;
assign a7366 = a7364 & ~a4690;
assign a7368 = a7364 & a4690;
assign a7370 = ~a7306 & a7176;
assign a7372 = a7306 & ~a7212;
assign a7374 = ~a7372 & ~a7370;
assign a7376 = ~a7374 & ~a4690;
assign a7378 = ~a7376 & ~a7368;
assign a7380 = ~a7378 & a4464;
assign a7382 = ~a7380 & ~a7366;
assign a7384 = ~a7382 & a7362;
assign a7386 = ~a4900 & ~a4706;
assign a7388 = ~a4944 & ~a4908;
assign a7390 = ~a7388 & a4706;
assign a7392 = ~a7390 & ~a7386;
assign a7394 = ~a7374 & a4690;
assign a7396 = ~a7306 & ~a7212;
assign a7398 = a7306 & ~a7254;
assign a7400 = ~a7398 & ~a7396;
assign a7402 = ~a7400 & ~a4690;
assign a7404 = ~a7402 & ~a7394;
assign a7406 = ~a7378 & ~a4464;
assign a7408 = ~a7406 & a7404;
assign a7410 = ~a7400 & a4690;
assign a7412 = ~a7306 & ~a7254;
assign a7414 = a7412 & ~a4690;
assign a7416 = ~a7414 & ~a7410;
assign a7418 = ~a7416 & a4464;
assign a7420 = ~a7418 & a7408;
assign a7422 = ~a7420 & a7392;
assign a7424 = ~a7422 & ~a7384;
assign a7426 = ~a7388 & ~a4706;
assign a7428 = ~a4942 & a4706;
assign a7430 = ~a7428 & ~a7426;
assign a7432 = a7412 & a4690;
assign a7434 = ~a7416 & ~a4464;
assign a7436 = ~a7434 & ~a7432;
assign a7438 = ~a7436 & a7430;
assign a7440 = ~a7438 & i488;
assign a7442 = a7440 & a7424;
assign a7444 = ~a7362 & ~a4644;
assign a7446 = a7306 & a7168;
assign a7448 = a7446 & ~a4690;
assign a7450 = a7446 & a4690;
assign a7452 = ~a7306 & a7168;
assign a7454 = a7306 & ~a7266;
assign a7456 = ~a7454 & ~a7452;
assign a7458 = ~a7456 & ~a4690;
assign a7460 = ~a7458 & ~a7450;
assign a7462 = ~a7460 & a4464;
assign a7464 = ~a7462 & ~a7448;
assign a7466 = ~a7464 & ~a7444;
assign a7468 = ~a7430 & ~a4644;
assign a7470 = ~a7306 & ~a7244;
assign a7472 = a7470 & a4690;
assign a7474 = ~a7306 & ~a7266;
assign a7476 = a7306 & ~a7244;
assign a7478 = ~a7476 & ~a7474;
assign a7480 = ~a7478 & a4690;
assign a7482 = a7470 & ~a4690;
assign a7484 = ~a7482 & ~a7480;
assign a7486 = ~a7484 & ~a4464;
assign a7488 = ~a7486 & ~a7472;
assign a7490 = ~a7488 & ~a7468;
assign a7492 = ~a7490 & ~a7466;
assign a7494 = ~a7456 & a4690;
assign a7496 = ~a7478 & ~a4690;
assign a7498 = ~a7496 & ~a7494;
assign a7500 = ~a7460 & ~a4464;
assign a7502 = ~a7500 & a7498;
assign a7504 = ~a7484 & a4464;
assign a7506 = ~a7504 & a7502;
assign a7508 = ~a7392 & ~a4644;
assign a7510 = ~a7508 & ~a7506;
assign a7512 = ~a7510 & a7492;
assign a7514 = a7512 & a7442;
assign a7516 = ~a7506 & ~a7444;
assign a7518 = ~a7508 & ~a7488;
assign a7520 = ~a7518 & ~a7516;
assign a7522 = ~a7060 & ~a4706;
assign a7524 = ~a7356 & a4706;
assign a7526 = ~a7524 & ~a7522;
assign a7528 = ~a7526 & ~a4644;
assign a7530 = ~a7528 & ~a7464;
assign a7532 = ~a7530 & a7520;
assign a7534 = ~a7436 & a7392;
assign a7536 = ~a7534 & a7532;
assign a7538 = ~a7420 & a7362;
assign a7540 = ~a7538 & a7536;
assign a7542 = a7526 & ~a7382;
assign a7544 = ~a7542 & a7540;
assign a7546 = a7544 & ~a7514;
assign a7548 = ~a7546 & a4706;
assign a7550 = a7546 & ~a4706;
assign a7552 = ~a7550 & ~a7548;
assign a7554 = ~a7320 & ~a7310;
assign a7556 = a7554 & ~a7552;
assign a7558 = ~a7554 & ~a7548;
assign a7560 = a7558 & ~a7550;
assign a7562 = ~a7560 & ~a7556;
assign a7564 = a7562 & ~a7328;
assign a7566 = ~a7562 & a7328;
assign a7568 = ~a7566 & ~a7564;
assign a7570 = a7568 & ~a2246;
assign a7572 = ~a7570 & ~a7354;
assign a7574 = ~a7572 & ~a7134;
assign a7576 = ~a7340 & ~a4436;
assign a7578 = a7340 & a4436;
assign a7580 = ~a7578 & ~a7576;
assign a7582 = a7580 & a7134;
assign a7584 = ~a7582 & ~a7574;
assign a7586 = ~a7584 & ~l494;
assign a7588 = a5384 & l494;
assign a7592 = a4722 & a2246;
assign a7594 = a7546 & ~a7382;
assign a7596 = a7594 & ~a4706;
assign a7598 = a7594 & a4706;
assign a7600 = ~a7546 & ~a7382;
assign a7602 = a7546 & ~a7420;
assign a7604 = ~a7602 & ~a7600;
assign a7606 = ~a7604 & ~a4706;
assign a7608 = ~a7606 & ~a7598;
assign a7610 = ~a7608 & a4428;
assign a7612 = ~a7610 & ~a7596;
assign a7614 = ~a7612 & a5050;
assign a7616 = ~a4886 & ~a4722;
assign a7618 = ~a4934 & ~a4894;
assign a7620 = ~a7618 & a4722;
assign a7622 = ~a7620 & ~a7616;
assign a7624 = ~a7604 & a4706;
assign a7626 = ~a7546 & ~a7420;
assign a7628 = a7546 & ~a7436;
assign a7630 = ~a7628 & ~a7626;
assign a7632 = ~a7630 & ~a4706;
assign a7634 = ~a7632 & ~a7624;
assign a7636 = ~a7608 & ~a4428;
assign a7638 = ~a7636 & a7634;
assign a7640 = ~a7630 & a4706;
assign a7642 = ~a7546 & ~a7436;
assign a7644 = a7642 & ~a4706;
assign a7646 = ~a7644 & ~a7640;
assign a7648 = ~a7646 & a4428;
assign a7650 = ~a7648 & a7638;
assign a7652 = ~a7650 & a7622;
assign a7654 = ~a7652 & ~a7614;
assign a7656 = ~a7618 & ~a4722;
assign a7658 = ~a4932 & a4722;
assign a7660 = ~a7658 & ~a7656;
assign a7662 = a7642 & a4706;
assign a7664 = ~a7646 & ~a4428;
assign a7666 = ~a7664 & ~a7662;
assign a7668 = ~a7666 & a7660;
assign a7670 = ~a7668 & i490;
assign a7672 = a7670 & a7654;
assign a7674 = ~a5050 & ~a4644;
assign a7676 = a7546 & ~a7464;
assign a7678 = a7676 & ~a4706;
assign a7680 = a7676 & a4706;
assign a7682 = ~a7546 & ~a7464;
assign a7684 = a7546 & ~a7506;
assign a7686 = ~a7684 & ~a7682;
assign a7688 = ~a7686 & ~a4706;
assign a7690 = ~a7688 & ~a7680;
assign a7692 = ~a7690 & a4428;
assign a7694 = ~a7692 & ~a7678;
assign a7696 = ~a7694 & ~a7674;
assign a7698 = ~a7660 & ~a4644;
assign a7700 = ~a7546 & ~a7488;
assign a7702 = a7700 & a4706;
assign a7704 = ~a7546 & ~a7506;
assign a7706 = a7546 & ~a7488;
assign a7708 = ~a7706 & ~a7704;
assign a7710 = ~a7708 & a4706;
assign a7712 = a7700 & ~a4706;
assign a7714 = ~a7712 & ~a7710;
assign a7716 = ~a7714 & ~a4428;
assign a7718 = ~a7716 & ~a7702;
assign a7720 = ~a7718 & ~a7698;
assign a7722 = ~a7720 & ~a7696;
assign a7724 = ~a7686 & a4706;
assign a7726 = ~a7708 & ~a4706;
assign a7728 = ~a7726 & ~a7724;
assign a7730 = ~a7690 & ~a4428;
assign a7732 = ~a7730 & a7728;
assign a7734 = ~a7714 & a4428;
assign a7736 = ~a7734 & a7732;
assign a7738 = ~a7622 & ~a4644;
assign a7740 = ~a7738 & ~a7736;
assign a7742 = ~a7740 & a7722;
assign a7744 = a7742 & a7672;
assign a7746 = ~a7736 & ~a7674;
assign a7748 = ~a7738 & ~a7718;
assign a7750 = ~a7748 & ~a7746;
assign a7752 = a5042 & ~a4644;
assign a7754 = ~a7752 & ~a7694;
assign a7756 = ~a7754 & a7750;
assign a7758 = ~a7666 & a7622;
assign a7760 = ~a7758 & a7756;
assign a7762 = ~a7650 & a5050;
assign a7764 = ~a7762 & a7760;
assign a7766 = ~a7612 & ~a5042;
assign a7768 = ~a7766 & a7764;
assign a7770 = a7768 & ~a7744;
assign a7772 = a7770 & ~a4722;
assign a7774 = ~a7770 & a4722;
assign a7776 = ~a7774 & ~a7772;
assign a7778 = ~a7558 & ~a7550;
assign a7780 = a7778 & ~a7776;
assign a7782 = ~a7778 & a7776;
assign a7784 = ~a7782 & ~a7780;
assign a7786 = a7784 & ~a7566;
assign a7788 = ~a7784 & a7566;
assign a7790 = ~a7788 & ~a7786;
assign a7792 = a7790 & ~a2246;
assign a7794 = ~a7792 & ~a7592;
assign a7796 = ~a7794 & ~a7134;
assign a7798 = ~a7578 & ~a4398;
assign a7800 = a7578 & a4398;
assign a7802 = ~a7800 & ~a7798;
assign a7804 = a7802 & a7134;
assign a7806 = ~a7804 & ~a7796;
assign a7808 = ~a7806 & ~l494;
assign a7810 = a5392 & l494;
assign a7814 = a4738 & a2246;
assign a7816 = ~a7778 & ~a7774;
assign a7818 = ~a7816 & ~a7772;
assign a7820 = ~a7818 & ~a4738;
assign a7822 = a7818 & a4738;
assign a7824 = ~a7822 & ~a7820;
assign a7826 = ~a7824 & ~a7788;
assign a7828 = a7824 & a7788;
assign a7830 = ~a7828 & ~a7826;
assign a7832 = a7830 & ~a2246;
assign a7834 = ~a7832 & ~a7814;
assign a7836 = ~a7834 & ~a7134;
assign a7838 = ~a7800 & ~a2542;
assign a7840 = a7800 & a2542;
assign a7842 = ~a7840 & ~a7838;
assign a7844 = a7842 & a7134;
assign a7846 = ~a7844 & ~a7836;
assign a7848 = ~a7846 & ~l494;
assign a7850 = a5394 & l494;
assign a7854 = ~a6908 & a2268;
assign a7856 = ~a6906 & i196;
assign a7858 = a6906 & a6882;
assign a7860 = ~a7858 & ~a7856;
assign a7862 = ~a7860 & a6908;
assign a7866 = ~a7822 & ~a4752;
assign a7868 = ~a7866 & a7828;
assign a7870 = a7822 & a4752;
assign a7872 = ~a7870 & ~a7868;
assign a7874 = ~a7872 & ~a2246;
assign a7876 = ~a7874 & a4760;
assign a7878 = a7874 & ~a4760;
assign a7880 = ~a7878 & ~a7876;
assign a7882 = ~a7880 & ~a7134;
assign a7884 = a7840 & a2526;
assign a7886 = a7884 & ~a2266;
assign a7888 = ~a7884 & a2266;
assign a7890 = ~a7888 & ~a7886;
assign a7892 = ~a7890 & a7134;
assign a7894 = ~a7892 & ~a7882;
assign a7896 = ~a7894 & ~l494;
assign a7898 = a5398 & l494;
assign a7902 = a4752 & a2246;
assign a7904 = ~a7870 & ~a7866;
assign a7906 = ~a7904 & a7828;
assign a7908 = a7904 & ~a7828;
assign a7910 = ~a7908 & ~a7906;
assign a7912 = ~a7910 & ~a2246;
assign a7914 = ~a7912 & ~a7902;
assign a7916 = ~a7914 & ~a7134;
assign a7918 = ~a7840 & ~a2526;
assign a7920 = ~a7918 & ~a7884;
assign a7922 = a7920 & a7134;
assign a7924 = ~a7922 & ~a7916;
assign a7926 = ~a7924 & ~l494;
assign a7928 = a5396 & l494;
assign a7932 = ~a6908 & a2548;
assign a7934 = ~a6906 & i182;
assign a7936 = a6906 & a6714;
assign a7938 = ~a7936 & ~a7934;
assign a7940 = ~a7938 & a6908;
assign a7944 = ~a6908 & a4404;
assign a7946 = ~a6906 & i184;
assign a7948 = a6906 & a6720;
assign a7950 = ~a7948 & ~a7946;
assign a7952 = ~a7950 & a6908;
assign a7956 = ~a6908 & a2566;
assign a7958 = ~a6906 & i186;
assign a7960 = a6906 & a6726;
assign a7962 = ~a7960 & ~a7958;
assign a7964 = ~a7962 & a6908;
assign a7968 = ~a6908 & a4428;
assign a7970 = ~a6906 & i188;
assign a7972 = a6906 & a6744;
assign a7974 = ~a7972 & ~a7970;
assign a7976 = ~a7974 & a6908;
assign a7980 = ~a6908 & a4464;
assign a7982 = ~a6906 & i190;
assign a7984 = a6906 & a6806;
assign a7986 = ~a7984 & ~a7982;
assign a7988 = ~a7986 & a6908;
assign a7992 = ~a6908 & a4536;
assign a7994 = ~a6906 & i194;
assign a7996 = a6906 & a6852;
assign a7998 = ~a7996 & ~a7994;
assign a8000 = ~a7998 & a6908;
assign a8004 = a4656 & a2246;
assign a8006 = ~a7122 & ~a2246;
assign a8008 = ~a8006 & ~a8004;
assign a8010 = ~a8008 & ~a7134;
assign a8012 = a7134 & ~a4544;
assign a8014 = ~a8012 & ~a8010;
assign a8016 = ~a8014 & ~l494;
assign a8018 = a5514 & l494;
assign a8022 = ~l494 & i206;
assign a8024 = ~a1698 & i208;
assign a8026 = ~a8024 & ~i14;
assign a8028 = ~a8026 & ~l1686;
assign a8030 = l1686 & l944;
assign a8032 = ~a8030 & ~a8028;
assign a8034 = l1686 & ~l878;
assign a8036 = a8034 & ~l494;
assign a8038 = ~a8036 & ~a7898;
assign a8040 = ~a8038 & ~a6908;
assign a8044 = a8042 & i350;
assign a8046 = ~a6592 & l972;
assign a8048 = ~l998 & ~l988;
assign a8050 = l1686 & ~l1006;
assign a8052 = l1686 & ~l1002;
assign a8054 = l1686 & ~l1004;
assign a8056 = a8054 & a8052;
assign a8058 = ~a1704 & ~l1686;
assign a8060 = l1686 & l1064;
assign a8062 = ~a8060 & ~a8058;
assign a8064 = ~a6732 & ~l1686;
assign a8066 = l1686 & l1066;
assign a8068 = ~a8066 & ~a8064;
assign a8070 = ~a8068 & ~a8032;
assign a8072 = a8070 & a8062;
assign a8074 = i132 & ~i90;
assign a8076 = ~a8074 & ~a4212;
assign a8078 = ~i132 & i90;
assign a8080 = ~a8078 & ~a8076;
assign a8082 = a8080 & a3838;
assign a8084 = ~a1716 & a1704;
assign a8086 = ~a3828 & a1716;
assign a8088 = ~a8086 & ~a8084;
assign a8090 = ~a8088 & ~a1698;
assign a8092 = ~a8090 & ~a1802;
assign a8094 = a8084 & ~a3776;
assign a8096 = a8094 & a3828;
assign a8098 = ~a3828 & ~a3782;
assign a8100 = ~a8098 & ~a8096;
assign a8102 = a8100 & ~a8092;
assign a8104 = ~a8102 & a3852;
assign a8106 = ~a8090 & ~a1886;
assign a8108 = a8084 & ~a3878;
assign a8110 = a8108 & a3828;
assign a8112 = ~a3884 & ~a3828;
assign a8114 = ~a8112 & ~a8110;
assign a8116 = a8114 & ~a8106;
assign a8118 = ~a8116 & a3922;
assign a8120 = ~a8118 & ~a8104;
assign a8122 = a8116 & ~a3922;
assign a8124 = ~a8122 & ~a8120;
assign a8126 = ~a8090 & ~a1970;
assign a8128 = a8084 & ~a3952;
assign a8130 = a8128 & a3828;
assign a8132 = ~a3958 & ~a3828;
assign a8134 = ~a8132 & ~a8130;
assign a8136 = a8134 & ~a8126;
assign a8138 = ~a8136 & a4000;
assign a8140 = ~a8138 & ~a8124;
assign a8142 = a8136 & ~a4000;
assign a8144 = ~a8142 & ~a8140;
assign a8146 = ~a4036 & ~a3828;
assign a8148 = ~a8090 & ~a2052;
assign a8150 = a8084 & ~a4030;
assign a8152 = a8150 & a3828;
assign a8154 = ~a8152 & ~a8148;
assign a8156 = a8154 & ~a8146;
assign a8158 = ~a8156 & a4078;
assign a8160 = ~a8158 & ~a8144;
assign a8162 = a8156 & ~a4078;
assign a8164 = ~a8162 & ~a8160;
assign a8166 = ~a4114 & ~a3828;
assign a8168 = ~a8090 & ~a2134;
assign a8170 = a8084 & ~a4108;
assign a8172 = a8170 & a3828;
assign a8174 = ~a8172 & ~a8168;
assign a8176 = a8174 & ~a8166;
assign a8178 = ~a8176 & a4156;
assign a8180 = ~a8178 & ~a8164;
assign a8182 = a8176 & ~a4156;
assign a8184 = ~a8182 & ~a8180;
assign a8186 = ~a4188 & ~a3828;
assign a8188 = ~a8090 & a2192;
assign a8190 = a8084 & ~a4182;
assign a8192 = a8190 & a3828;
assign a8194 = ~a8192 & ~a8188;
assign a8196 = a8194 & ~a8186;
assign a8198 = ~a8196 & a4226;
assign a8200 = ~a8198 & ~a8184;
assign a8202 = a8196 & ~a4226;
assign a8204 = ~a8202 & ~a8200;
assign a8206 = ~a8090 & a2184;
assign a8208 = a3828 & i8;
assign a8210 = a8208 & a2182;
assign a8212 = ~a8210 & ~a8206;
assign a8214 = a8212 & ~a8204;
assign a8216 = ~a8214 & ~a8082;
assign a8218 = a8090 & i242;
assign a8220 = a8218 & ~a8216;
assign a8222 = a8220 & a3828;
assign a8224 = a8220 & ~a3828;
assign a8226 = ~a8220 & a3828;
assign a8228 = ~a8226 & ~a8224;
assign a8230 = ~a6732 & ~a1730;
assign a8232 = ~a8230 & ~a6750;
assign a8234 = ~a8232 & a8228;
assign a8236 = ~a8222 & a5550;
assign a8238 = ~a8236 & ~a8234;
assign a8240 = ~a8238 & ~a6732;
assign a8242 = ~a8240 & ~a1814;
assign a8244 = a8228 & ~a8222;
assign a8246 = ~a6764 & a1720;
assign a8248 = a8246 & a8228;
assign a8250 = a1704 & i62;
assign a8252 = a8250 & a1716;
assign a8254 = a8252 & ~a6764;
assign a8256 = ~a8254 & ~a8094;
assign a8258 = ~a8256 & ~a8228;
assign a8260 = ~a8258 & ~a8248;
assign a8262 = ~a8260 & ~a8244;
assign a8264 = a1718 & ~a1704;
assign a8266 = a8264 & ~a6764;
assign a8268 = ~a8266 & a3782;
assign a8270 = ~a8268 & a8244;
assign a8272 = ~a8270 & ~a8262;
assign a8274 = a8272 & ~a8242;
assign a8276 = i248 & ~i246;
assign a8278 = i254 & i252;
assign a8280 = a8278 & i250;
assign a8282 = a8280 & a8276;
assign a8284 = ~a8282 & i244;
assign a8286 = ~a8256 & a8222;
assign a8288 = ~a8268 & ~a8228;
assign a8290 = ~a8288 & ~a8286;
assign a8292 = a8290 & a8284;
assign a8294 = ~a8292 & a6732;
assign a8296 = a3838 & ~i256;
assign a8298 = ~i260 & i258;
assign a8300 = a8298 & a8216;
assign a8302 = a8300 & ~a8296;
assign a8304 = ~a8274 & a3852;
assign a8306 = ~a8240 & ~a1912;
assign a8308 = ~a6756 & a1720;
assign a8310 = a8308 & a8228;
assign a8312 = a8252 & ~a6756;
assign a8314 = ~a8312 & ~a8108;
assign a8316 = ~a8314 & ~a8228;
assign a8318 = ~a8316 & ~a8310;
assign a8320 = ~a8318 & ~a8244;
assign a8322 = a8264 & ~a6756;
assign a8324 = ~a8322 & a3884;
assign a8326 = ~a8324 & a8244;
assign a8328 = ~a8326 & ~a8320;
assign a8330 = a8328 & ~a8306;
assign a8332 = ~a8330 & a3922;
assign a8334 = ~a8332 & ~a8304;
assign a8336 = a8330 & ~a3922;
assign a8338 = ~a8336 & ~a8334;
assign a8340 = ~a8240 & ~a1994;
assign a8342 = ~a6778 & a1720;
assign a8344 = a8342 & a8228;
assign a8346 = a8252 & ~a6778;
assign a8348 = ~a8346 & ~a8128;
assign a8350 = ~a8348 & ~a8228;
assign a8352 = ~a8350 & ~a8344;
assign a8354 = ~a8352 & ~a8244;
assign a8356 = a8264 & ~a6778;
assign a8358 = ~a8356 & a3958;
assign a8360 = ~a8358 & a8244;
assign a8362 = ~a8360 & ~a8354;
assign a8364 = a8362 & ~a8340;
assign a8366 = ~a8364 & a4000;
assign a8368 = ~a8366 & ~a8338;
assign a8370 = a8364 & ~a4000;
assign a8372 = ~a8370 & ~a8368;
assign a8374 = ~a8240 & ~a2076;
assign a8376 = ~a2076 & i62;
assign a8378 = i262 & ~i62;
assign a8380 = ~a8378 & ~a8376;
assign a8382 = ~a8380 & a1720;
assign a8384 = a8382 & a8228;
assign a8386 = ~a8380 & a8252;
assign a8388 = ~a8386 & ~a8150;
assign a8390 = ~a8388 & ~a8228;
assign a8392 = ~a8390 & ~a8384;
assign a8394 = ~a8392 & ~a8244;
assign a8396 = ~a8380 & a8264;
assign a8398 = ~a8396 & a4036;
assign a8400 = ~a8398 & a8244;
assign a8402 = ~a8400 & ~a8394;
assign a8404 = a8402 & ~a8374;
assign a8406 = ~a8404 & a4078;
assign a8408 = ~a8406 & ~a8372;
assign a8410 = a8404 & ~a4078;
assign a8412 = ~a8410 & ~a8408;
assign a8414 = ~a8240 & ~a2158;
assign a8416 = ~a2158 & i62;
assign a8418 = i264 & ~i62;
assign a8420 = ~a8418 & ~a8416;
assign a8422 = ~a8420 & a1720;
assign a8424 = a8422 & a8228;
assign a8426 = ~a8420 & a8252;
assign a8428 = ~a8426 & ~a8170;
assign a8430 = ~a8428 & ~a8228;
assign a8432 = ~a8430 & ~a8424;
assign a8434 = ~a8432 & ~a8244;
assign a8436 = ~a8420 & a8264;
assign a8438 = ~a8436 & a4114;
assign a8440 = ~a8438 & a8244;
assign a8442 = ~a8440 & ~a8434;
assign a8444 = a8442 & ~a8414;
assign a8446 = ~a8444 & a4156;
assign a8448 = ~a8446 & ~a8412;
assign a8450 = a8444 & ~a4156;
assign a8452 = ~a8450 & ~a8448;
assign a8454 = ~a8240 & ~a2214;
assign a8456 = ~a2214 & i62;
assign a8458 = i266 & ~i62;
assign a8460 = ~a8458 & ~a8456;
assign a8462 = ~a8460 & a1720;
assign a8464 = a8462 & a8228;
assign a8466 = ~a8460 & a8252;
assign a8468 = ~a8466 & ~a8190;
assign a8470 = ~a8468 & ~a8228;
assign a8472 = ~a8470 & ~a8464;
assign a8474 = ~a8472 & ~a8244;
assign a8476 = ~a8460 & a8264;
assign a8478 = ~a8476 & a4188;
assign a8480 = ~a8478 & a8244;
assign a8482 = ~a8480 & ~a8474;
assign a8484 = a8482 & ~a8454;
assign a8486 = ~a8484 & a4226;
assign a8488 = ~a8486 & ~a8452;
assign a8490 = a8484 & ~a4226;
assign a8492 = ~a8490 & ~a8488;
assign a8494 = ~a8240 & ~a2232;
assign a8496 = ~a2232 & i62;
assign a8498 = i268 & ~i62;
assign a8500 = ~a8498 & ~a8496;
assign a8502 = ~a8500 & a1720;
assign a8504 = a8502 & a8228;
assign a8506 = a2184 & i8;
assign a8508 = ~a8500 & a8252;
assign a8510 = ~a8508 & ~a8506;
assign a8512 = ~a8510 & ~a8228;
assign a8514 = ~a8512 & ~a8504;
assign a8516 = ~a8514 & ~a8244;
assign a8518 = ~a8516 & ~a8494;
assign a8520 = ~a8518 & ~a8082;
assign a8522 = ~a8520 & ~a8492;
assign a8524 = a8518 & a8082;
assign a8526 = ~a8524 & a8296;
assign a8528 = a8526 & ~a8522;
assign a8530 = ~a8528 & ~a8302;
assign a8532 = ~a8530 & ~a8284;
assign a8534 = ~a8532 & a3852;
assign a8536 = ~a8284 & ~a3852;
assign a8538 = a8536 & ~a8530;
assign a8540 = ~a8538 & ~a6732;
assign a8542 = a8540 & ~a8534;
assign a8544 = ~a8542 & ~a8294;
assign a8546 = a8544 & ~a8274;
assign a8548 = ~a8314 & a8222;
assign a8550 = ~a8324 & ~a8228;
assign a8552 = ~a8550 & ~a8548;
assign a8554 = a8552 & i250;
assign a8556 = ~a8290 & ~a8284;
assign a8558 = ~a8552 & ~i250;
assign a8560 = ~a8558 & ~a8556;
assign a8562 = a8560 & ~a8554;
assign a8564 = ~a8558 & ~a8554;
assign a8566 = ~a8564 & a8556;
assign a8568 = ~a8566 & ~a8562;
assign a8570 = ~a8568 & a6732;
assign a8572 = a3922 & i250;
assign a8574 = ~a3922 & ~i250;
assign a8576 = ~a8574 & ~a8536;
assign a8578 = a8576 & ~a8572;
assign a8580 = ~a8574 & ~a8572;
assign a8582 = ~a8580 & a8536;
assign a8584 = ~a8582 & ~a8578;
assign a8586 = ~a8584 & ~a8530;
assign a8588 = a8530 & ~a3922;
assign a8590 = ~a8588 & ~a8586;
assign a8592 = ~a8590 & ~a6732;
assign a8594 = ~a8592 & ~a8570;
assign a8596 = a8594 & ~a8330;
assign a8598 = ~a8596 & ~a8546;
assign a8600 = ~a8594 & a8330;
assign a8602 = ~a8600 & ~a8598;
assign a8604 = ~a8560 & ~a8554;
assign a8606 = ~a8348 & a8222;
assign a8608 = ~a8358 & ~a8228;
assign a8610 = ~a8608 & ~a8606;
assign a8612 = a8610 & i248;
assign a8614 = ~a8610 & ~i248;
assign a8616 = ~a8614 & ~a8612;
assign a8618 = a8616 & ~a8604;
assign a8620 = ~a8616 & a8604;
assign a8622 = ~a8620 & ~a8618;
assign a8624 = ~a8622 & a6732;
assign a8626 = ~a8576 & ~a8572;
assign a8628 = a4000 & i248;
assign a8630 = ~a4000 & ~i248;
assign a8632 = ~a8630 & ~a8628;
assign a8634 = a8632 & ~a8626;
assign a8636 = ~a8632 & a8626;
assign a8638 = ~a8636 & ~a8634;
assign a8640 = ~a8638 & ~a8530;
assign a8642 = a8530 & ~a4000;
assign a8644 = ~a8642 & ~a8640;
assign a8646 = ~a8644 & ~a6732;
assign a8648 = ~a8646 & ~a8624;
assign a8650 = a8648 & ~a8364;
assign a8652 = ~a8650 & ~a8602;
assign a8654 = ~a8648 & a8364;
assign a8656 = ~a8654 & ~a8652;
assign a8658 = ~a8614 & ~a8604;
assign a8660 = ~a8658 & ~a8612;
assign a8662 = ~a8388 & a8222;
assign a8664 = ~a8398 & ~a8228;
assign a8666 = ~a8664 & ~a8662;
assign a8668 = a8666 & i252;
assign a8670 = ~a8666 & ~i252;
assign a8672 = ~a8670 & ~a8668;
assign a8674 = a8672 & ~a8660;
assign a8676 = ~a8672 & a8660;
assign a8678 = ~a8676 & ~a8674;
assign a8680 = ~a8678 & a6732;
assign a8682 = ~a8630 & ~a8626;
assign a8684 = ~a8682 & ~a8628;
assign a8686 = a4078 & i252;
assign a8688 = ~a4078 & ~i252;
assign a8690 = ~a8688 & ~a8686;
assign a8692 = a8690 & ~a8684;
assign a8694 = ~a8690 & a8684;
assign a8696 = ~a8694 & ~a8692;
assign a8698 = ~a8696 & ~a8530;
assign a8700 = a8530 & ~a4078;
assign a8702 = ~a8700 & ~a8698;
assign a8704 = ~a8702 & ~a6732;
assign a8706 = ~a8704 & ~a8680;
assign a8708 = a8706 & ~a8404;
assign a8710 = ~a8708 & ~a8656;
assign a8712 = ~a8706 & a8404;
assign a8714 = ~a8712 & ~a8710;
assign a8716 = ~a8670 & ~a8660;
assign a8718 = ~a8716 & ~a8668;
assign a8720 = ~a8428 & a8222;
assign a8722 = ~a8438 & ~a8228;
assign a8724 = ~a8722 & ~a8720;
assign a8726 = a8724 & i254;
assign a8728 = ~a8724 & ~i254;
assign a8730 = ~a8728 & ~a8726;
assign a8732 = a8730 & ~a8718;
assign a8734 = ~a8730 & a8718;
assign a8736 = ~a8734 & ~a8732;
assign a8738 = ~a8736 & a6732;
assign a8740 = ~a8688 & ~a8684;
assign a8742 = ~a8740 & ~a8686;
assign a8744 = a4156 & i254;
assign a8746 = ~a4156 & ~i254;
assign a8748 = ~a8746 & ~a8744;
assign a8750 = a8748 & ~a8742;
assign a8752 = ~a8748 & a8742;
assign a8754 = ~a8752 & ~a8750;
assign a8756 = ~a8754 & ~a8530;
assign a8758 = a8530 & ~a4156;
assign a8760 = ~a8758 & ~a8756;
assign a8762 = ~a8760 & ~a6732;
assign a8764 = ~a8762 & ~a8738;
assign a8766 = a8764 & ~a8444;
assign a8768 = ~a8766 & ~a8714;
assign a8770 = ~a8764 & a8444;
assign a8772 = ~a8770 & ~a8768;
assign a8774 = ~a8728 & ~a8718;
assign a8776 = ~a8774 & ~a8726;
assign a8778 = ~a8468 & a8222;
assign a8780 = ~a8478 & ~a8228;
assign a8782 = ~a8780 & ~a8778;
assign a8784 = ~a8782 & ~i246;
assign a8786 = a8782 & i246;
assign a8788 = ~a8786 & ~a8784;
assign a8790 = ~a8788 & ~a8776;
assign a8792 = a8788 & a8776;
assign a8794 = ~a8792 & ~a8790;
assign a8796 = ~a8794 & a6732;
assign a8798 = ~a8746 & ~a8742;
assign a8800 = ~a8798 & ~a8744;
assign a8802 = a4226 & ~i246;
assign a8804 = ~a4226 & i246;
assign a8806 = ~a8804 & ~a8802;
assign a8808 = a8806 & ~a8800;
assign a8810 = ~a8806 & a8800;
assign a8812 = ~a8810 & ~a8808;
assign a8814 = ~a8812 & ~a8530;
assign a8816 = a8530 & ~a4226;
assign a8818 = ~a8816 & ~a8814;
assign a8820 = ~a8818 & ~a6732;
assign a8822 = ~a8820 & ~a8796;
assign a8824 = a8822 & ~a8484;
assign a8826 = ~a8824 & ~a8772;
assign a8828 = ~a8822 & a8484;
assign a8830 = ~a8828 & ~a8826;
assign a8832 = ~a8804 & ~a8800;
assign a8834 = ~a8832 & ~a8802;
assign a8836 = a8834 & ~a8530;
assign a8838 = ~a8836 & a8520;
assign a8840 = ~a8838 & ~a8830;
assign a8842 = ~a8836 & ~a8082;
assign a8844 = ~a8842 & a8518;
assign a8846 = ~a8844 & ~a8840;
assign a8848 = a8240 & i270;
assign a8850 = a8848 & ~a8846;
assign a8852 = a8850 & ~a8228;
assign a8854 = ~a8852 & ~a8222;
assign a8856 = a8854 & ~l1686;
assign a8858 = l1686 & l1060;
assign a8860 = ~a8858 & ~a8856;
assign a8862 = l1686 & ~l1058;
assign a8864 = l1686 & ~l1008;
assign a8866 = l1686 & ~l1010;
assign a8868 = l1686 & ~l992;
assign a8870 = l1686 & ~l1012;
assign a8872 = l1686 & ~l1014;
assign a8874 = l1686 & ~l1020;
assign a8876 = a1712 & i14;
assign a8878 = a4384 & a3760;
assign a8880 = a8878 & a3864;
assign a8882 = ~a8878 & ~a3864;
assign a8884 = ~a8882 & ~a8880;
assign a8886 = a4384 & a4260;
assign a8888 = ~a8886 & ~a3930;
assign a8890 = a8886 & a3930;
assign a8892 = ~a8890 & ~a8888;
assign a8894 = ~a8892 & ~a8880;
assign a8896 = a8892 & a8880;
assign a8898 = ~a8896 & ~a8894;
assign a8900 = ~a8890 & ~a8880;
assign a8902 = ~a8900 & ~a8888;
assign a8904 = a4384 & a4286;
assign a8906 = ~a8904 & ~a4008;
assign a8908 = a8904 & a4008;
assign a8910 = ~a8908 & ~a8906;
assign a8912 = ~a8910 & ~a8902;
assign a8914 = a8910 & a8902;
assign a8916 = ~a8914 & ~a8912;
assign a8918 = ~a8908 & ~a8902;
assign a8920 = ~a8918 & ~a8906;
assign a8922 = a4384 & a4312;
assign a8924 = ~a8922 & ~a4086;
assign a8926 = a8922 & a4086;
assign a8928 = ~a8926 & ~a8924;
assign a8930 = ~a8928 & ~a8920;
assign a8932 = a8928 & a8920;
assign a8934 = ~a8932 & ~a8930;
assign a8936 = a4384 & a3758;
assign a8938 = ~a8936 & ~a4164;
assign a8940 = ~a8926 & ~a8920;
assign a8942 = ~a8940 & ~a8924;
assign a8944 = a8936 & a4164;
assign a8946 = ~a8944 & ~a8942;
assign a8948 = ~a8946 & ~a8938;
assign a8950 = ~a8948 & ~a4230;
assign a8952 = ~a8944 & ~a8938;
assign a8954 = ~a8952 & ~a8942;
assign a8956 = a8952 & a8942;
assign a8958 = ~a8956 & ~a8954;
assign a8960 = a8958 & ~a8950;
assign a8962 = a8960 & a8934;
assign a8964 = a8962 & a8916;
assign a8966 = a8964 & a8898;
assign a8968 = a8966 & a8884;
assign a8970 = ~i222 & ~i220;
assign a8972 = ~a8970 & i224;
assign a8974 = i228 & i226;
assign a8976 = i232 & i230;
assign a8978 = a8976 & a8974;
assign a8980 = a8978 & a8972;
assign a8982 = ~a8980 & ~i234;
assign a8984 = ~a8982 & ~a8884;
assign a8986 = i236 & i234;
assign a8988 = a8986 & i238;
assign a8990 = a8988 & i240;
assign a8992 = a8990 & i222;
assign a8994 = a8992 & i220;
assign a8996 = ~a8992 & ~i220;
assign a8998 = ~a8996 & ~a8980;
assign a9000 = a8998 & ~a8994;
assign a9002 = ~a9000 & ~a8884;
assign a9004 = a8994 & i232;
assign a9006 = ~a8994 & ~i232;
assign a9008 = ~a9006 & ~a9004;
assign a9010 = ~a9008 & ~a8980;
assign a9012 = a9010 & ~a8884;
assign a9014 = a9004 & i224;
assign a9016 = ~a9004 & ~i224;
assign a9018 = ~a9016 & ~a9014;
assign a9020 = ~a9018 & ~a8980;
assign a9022 = a9020 & ~a8884;
assign a9024 = a9014 & i230;
assign a9026 = ~a9014 & ~i230;
assign a9028 = ~a9026 & ~a9024;
assign a9030 = ~a9028 & ~a8980;
assign a9032 = a9030 & ~a8884;
assign a9034 = a9024 & i228;
assign a9036 = ~a9024 & ~i228;
assign a9038 = ~a9036 & ~a9034;
assign a9040 = ~a9038 & ~a8980;
assign a9042 = a9040 & ~a8884;
assign a9044 = ~a9034 & ~i226;
assign a9046 = a8966 & ~a8884;
assign a9048 = ~a9046 & ~a9044;
assign a9050 = ~a9048 & ~a8898;
assign a9052 = ~a9050 & ~a9042;
assign a9054 = a9048 & a8898;
assign a9056 = ~a9054 & ~a9052;
assign a9058 = ~a9056 & a8964;
assign a9060 = a9058 & ~a8884;
assign a9062 = ~a9060 & ~a9040;
assign a9064 = ~a9062 & ~a8898;
assign a9066 = ~a9064 & ~a9032;
assign a9068 = a9062 & a8898;
assign a9070 = ~a9068 & ~a9066;
assign a9072 = a9058 & ~a8898;
assign a9074 = ~a9072 & a9048;
assign a9076 = ~a9074 & ~a8916;
assign a9078 = ~a9076 & ~a9070;
assign a9080 = a9074 & a8916;
assign a9082 = ~a9080 & ~a9078;
assign a9084 = ~a9082 & a8962;
assign a9086 = a9084 & ~a8884;
assign a9088 = a9086 & a9030;
assign a9090 = ~a9086 & ~a9030;
assign a9092 = ~a9090 & ~a9088;
assign a9094 = a9092 & ~a8898;
assign a9096 = ~a9094 & ~a9022;
assign a9098 = ~a9092 & a8898;
assign a9100 = ~a9098 & ~a9096;
assign a9102 = ~a9100 & a8916;
assign a9104 = a9084 & ~a8898;
assign a9106 = a9104 & ~a9062;
assign a9108 = ~a9104 & a9062;
assign a9110 = ~a9108 & ~a9106;
assign a9112 = ~a9110 & ~a9088;
assign a9114 = a9100 & ~a8916;
assign a9116 = ~a9114 & a9112;
assign a9118 = ~a9116 & ~a9102;
assign a9120 = ~a9118 & a8934;
assign a9122 = a9084 & ~a8916;
assign a9124 = ~a9122 & a9074;
assign a9126 = a9124 & ~a9106;
assign a9128 = a9118 & ~a8934;
assign a9130 = ~a9128 & a9126;
assign a9132 = ~a9130 & ~a9120;
assign a9134 = ~a9132 & a8960;
assign a9136 = a9134 & ~a8884;
assign a9138 = ~a9136 & ~a9020;
assign a9140 = a9134 & a9022;
assign a9142 = ~a9140 & ~a9138;
assign a9144 = a9142 & ~a8898;
assign a9146 = ~a9144 & ~a9012;
assign a9148 = ~a9142 & a8898;
assign a9150 = ~a9148 & ~a9146;
assign a9152 = a9150 & ~a8916;
assign a9154 = a9134 & ~a8898;
assign a9156 = a9154 & a9092;
assign a9158 = ~a9154 & ~a9092;
assign a9160 = ~a9158 & ~a9156;
assign a9162 = ~a9160 & ~a9140;
assign a9164 = a9160 & a9140;
assign a9166 = ~a9164 & ~a9162;
assign a9168 = ~a9150 & a8916;
assign a9170 = ~a9168 & a9166;
assign a9172 = ~a9170 & ~a9152;
assign a9174 = a9172 & a8934;
assign a9176 = ~a9114 & ~a9102;
assign a9178 = a9176 & a9134;
assign a9180 = a9178 & a9112;
assign a9182 = ~a9178 & ~a9112;
assign a9184 = ~a9182 & ~a9180;
assign a9186 = ~a9172 & ~a8934;
assign a9188 = ~a9186 & a9184;
assign a9190 = ~a9188 & ~a9174;
assign a9192 = ~a9190 & a8958;
assign a9194 = a9134 & ~a9120;
assign a9196 = ~a9194 & a9126;
assign a9198 = a9190 & ~a8958;
assign a9200 = ~a9198 & a9196;
assign a9202 = ~a9200 & ~a9192;
assign a9204 = ~a9202 & ~a8950;
assign a9206 = a9204 & ~a8884;
assign a9208 = ~a9206 & ~a9010;
assign a9210 = a9204 & a9012;
assign a9212 = ~a9210 & ~a9208;
assign a9214 = a9212 & ~a8898;
assign a9216 = ~a9214 & ~a9002;
assign a9218 = ~a9212 & a8898;
assign a9220 = ~a9218 & ~a9216;
assign a9222 = a9220 & ~a8916;
assign a9224 = a9204 & ~a8898;
assign a9226 = a9224 & a9142;
assign a9228 = ~a9224 & ~a9142;
assign a9230 = ~a9228 & ~a9226;
assign a9232 = ~a9230 & ~a9210;
assign a9234 = a9230 & a9210;
assign a9236 = ~a9234 & ~a9232;
assign a9238 = ~a9220 & a8916;
assign a9240 = ~a9238 & a9236;
assign a9242 = ~a9240 & ~a9222;
assign a9244 = ~a9242 & ~a8934;
assign a9246 = a9242 & a8934;
assign a9248 = ~a9168 & ~a9152;
assign a9250 = a9248 & a9204;
assign a9252 = a9250 & a9166;
assign a9254 = ~a9250 & ~a9166;
assign a9256 = ~a9254 & ~a9252;
assign a9258 = a9256 & ~a9246;
assign a9260 = ~a9258 & ~a9244;
assign a9262 = ~a9260 & ~a8958;
assign a9264 = ~a9186 & ~a9174;
assign a9266 = a9264 & a9204;
assign a9268 = a9266 & a9184;
assign a9270 = ~a9266 & ~a9184;
assign a9272 = ~a9270 & ~a9268;
assign a9274 = a9260 & a8958;
assign a9276 = ~a9274 & ~a9272;
assign a9278 = ~a9276 & ~a9262;
assign a9280 = a9278 & ~a8950;
assign a9282 = ~a9278 & a8950;
assign a9284 = a9204 & ~a9192;
assign a9286 = ~a9284 & a9196;
assign a9288 = a9286 & ~a9282;
assign a9290 = ~a9288 & ~a9280;
assign a9292 = ~a9290 & a9002;
assign a9294 = ~a9290 & ~a8898;
assign a9296 = a9294 & a9212;
assign a9298 = ~a9294 & ~a9212;
assign a9300 = ~a9298 & ~a9296;
assign a9302 = ~a9300 & ~a9292;
assign a9304 = a9300 & a9292;
assign a9306 = ~a9304 & ~a9302;
assign a9308 = ~a8990 & ~i222;
assign a9310 = ~a9308 & ~a8992;
assign a9312 = ~a9310 & ~a8980;
assign a9314 = a9312 & ~a8884;
assign a9316 = ~a9290 & ~a8884;
assign a9318 = ~a9316 & a9000;
assign a9320 = ~a9318 & ~a9292;
assign a9322 = a9320 & ~a8898;
assign a9324 = ~a9322 & ~a9314;
assign a9326 = ~a9320 & a8898;
assign a9328 = ~a9326 & ~a9324;
assign a9330 = a9306 & ~a8916;
assign a9332 = ~a9330 & ~a9328;
assign a9334 = ~a9306 & a8916;
assign a9336 = ~a9334 & ~a9332;
assign a9338 = ~a9238 & ~a9222;
assign a9340 = a9338 & ~a9290;
assign a9342 = a9340 & a9236;
assign a9344 = ~a9340 & ~a9236;
assign a9346 = ~a9344 & ~a9342;
assign a9348 = a9346 & ~a8934;
assign a9350 = ~a9348 & ~a9336;
assign a9352 = ~a9346 & a8934;
assign a9354 = ~a9352 & ~a9350;
assign a9356 = ~a9246 & ~a9244;
assign a9358 = a9356 & ~a9290;
assign a9360 = a9358 & a9256;
assign a9362 = ~a9358 & ~a9256;
assign a9364 = ~a9362 & ~a9360;
assign a9366 = a9364 & ~a8958;
assign a9368 = ~a9366 & ~a9354;
assign a9370 = ~a9364 & a8958;
assign a9372 = ~a9370 & ~a9368;
assign a9374 = ~a9274 & ~a9262;
assign a9376 = a9374 & ~a9290;
assign a9378 = a9376 & ~a9272;
assign a9380 = ~a9376 & a9272;
assign a9382 = ~a9380 & ~a9378;
assign a9384 = a9382 & a8950;
assign a9386 = ~a9384 & ~a9372;
assign a9388 = ~a9382 & ~a8950;
assign a9390 = a9288 & ~a9280;
assign a9392 = ~a9390 & a9286;
assign a9394 = ~a9392 & ~a9388;
assign a9396 = a9394 & ~a9386;
assign a9398 = ~a9396 & ~a8916;
assign a9400 = a9398 & a9306;
assign a9402 = ~a9398 & ~a9306;
assign a9404 = ~a9402 & ~a9400;
assign a9406 = ~a9396 & ~a8898;
assign a9408 = ~a9406 & ~a9320;
assign a9410 = ~a9396 & ~a8884;
assign a9412 = a9410 & a9312;
assign a9414 = a9406 & a9320;
assign a9416 = ~a9414 & ~a9412;
assign a9418 = ~a9416 & ~a9408;
assign a9420 = ~a9418 & ~a9404;
assign a9422 = a9418 & a9404;
assign a9424 = ~a9422 & ~a9420;
assign a9426 = ~a8988 & ~i240;
assign a9428 = ~a8990 & ~a8980;
assign a9430 = a9428 & ~a9426;
assign a9432 = ~a9430 & ~a8884;
assign a9434 = ~a9410 & ~a9312;
assign a9436 = ~a9434 & ~a9412;
assign a9438 = a9436 & ~a8898;
assign a9440 = ~a9438 & ~a9432;
assign a9442 = ~a9436 & a8898;
assign a9444 = ~a9442 & ~a9440;
assign a9446 = a9444 & ~a8916;
assign a9448 = ~a9414 & ~a9408;
assign a9450 = ~a9448 & ~a9412;
assign a9452 = a9448 & a9412;
assign a9454 = ~a9452 & ~a9450;
assign a9456 = ~a9444 & a8916;
assign a9458 = ~a9456 & a9454;
assign a9460 = ~a9458 & ~a9446;
assign a9462 = a9460 & a8934;
assign a9464 = ~a9460 & ~a8934;
assign a9466 = ~a9464 & ~a9424;
assign a9468 = ~a9466 & ~a9462;
assign a9470 = a9468 & ~a8958;
assign a9472 = ~a9396 & ~a8934;
assign a9474 = a9472 & a9346;
assign a9476 = ~a9472 & ~a9346;
assign a9478 = ~a9476 & ~a9474;
assign a9480 = ~a9418 & ~a9400;
assign a9482 = ~a9480 & ~a9402;
assign a9484 = ~a9482 & ~a9478;
assign a9486 = a9482 & a9478;
assign a9488 = ~a9486 & ~a9484;
assign a9490 = ~a9468 & a8958;
assign a9492 = ~a9490 & a9488;
assign a9494 = ~a9492 & ~a9470;
assign a9496 = ~a9396 & ~a8958;
assign a9498 = a9496 & a9364;
assign a9500 = ~a9496 & ~a9364;
assign a9502 = ~a9500 & ~a9498;
assign a9504 = ~a9482 & ~a9474;
assign a9506 = ~a9504 & ~a9476;
assign a9508 = ~a9506 & ~a9502;
assign a9510 = a9506 & a9502;
assign a9512 = ~a9510 & ~a9508;
assign a9514 = a9512 & a8950;
assign a9516 = ~a9514 & a9494;
assign a9518 = ~a9396 & a8950;
assign a9520 = a9518 & a9382;
assign a9522 = ~a9518 & ~a9382;
assign a9524 = ~a9522 & ~a9520;
assign a9526 = ~a9506 & ~a9498;
assign a9528 = ~a9526 & ~a9500;
assign a9530 = ~a9528 & ~a9524;
assign a9532 = a9528 & a9524;
assign a9534 = ~a9512 & ~a8950;
assign a9536 = ~a9534 & ~a9532;
assign a9538 = a9536 & ~a9530;
assign a9540 = a9538 & ~a9516;
assign a9542 = ~a9464 & ~a9462;
assign a9544 = a9542 & ~a9540;
assign a9546 = a9544 & a9424;
assign a9548 = ~a9544 & ~a9424;
assign a9550 = ~a9548 & ~a9546;
assign a9552 = ~a8986 & ~i238;
assign a9554 = ~a9552 & ~a8988;
assign a9556 = a9554 & ~a8980;
assign a9558 = ~a9556 & ~a8884;
assign a9560 = ~a9540 & a9432;
assign a9562 = ~a9540 & ~a8884;
assign a9564 = ~a9562 & a9430;
assign a9566 = ~a9564 & ~a9560;
assign a9568 = a9566 & ~a8898;
assign a9570 = ~a9568 & ~a9558;
assign a9572 = ~a9566 & a8898;
assign a9574 = ~a9572 & ~a9570;
assign a9576 = a9574 & ~a8916;
assign a9578 = ~a9540 & ~a8898;
assign a9580 = ~a9578 & ~a9436;
assign a9582 = a9578 & a9436;
assign a9584 = ~a9582 & ~a9580;
assign a9586 = ~a9584 & ~a9560;
assign a9588 = a9584 & a9560;
assign a9590 = ~a9588 & ~a9586;
assign a9592 = ~a9574 & a8916;
assign a9594 = ~a9592 & a9590;
assign a9596 = ~a9594 & ~a9576;
assign a9598 = ~a9596 & ~a8934;
assign a9600 = ~a9456 & ~a9446;
assign a9602 = a9600 & ~a9540;
assign a9604 = a9602 & a9454;
assign a9606 = ~a9602 & ~a9454;
assign a9608 = ~a9606 & ~a9604;
assign a9610 = a9596 & a8934;
assign a9612 = ~a9610 & a9608;
assign a9614 = ~a9612 & ~a9598;
assign a9616 = ~a9614 & ~a8958;
assign a9618 = a9614 & a8958;
assign a9620 = ~a9618 & a9550;
assign a9622 = ~a9620 & ~a9616;
assign a9624 = ~a9490 & ~a9470;
assign a9626 = a9624 & ~a9540;
assign a9628 = a9626 & a9488;
assign a9630 = ~a9626 & ~a9488;
assign a9632 = ~a9630 & ~a9628;
assign a9634 = a9632 & a8950;
assign a9636 = ~a9634 & a9622;
assign a9638 = ~a9540 & a8950;
assign a9640 = a9638 & a9512;
assign a9642 = ~a9638 & ~a9512;
assign a9644 = ~a9642 & ~a9640;
assign a9646 = ~a9540 & ~a9494;
assign a9648 = ~a9646 & ~a9644;
assign a9650 = a9646 & a9644;
assign a9652 = ~a9632 & ~a8950;
assign a9654 = ~a9652 & ~a9650;
assign a9656 = a9654 & ~a9648;
assign a9658 = a9656 & ~a9636;
assign a9660 = ~a9618 & ~a9616;
assign a9662 = a9660 & ~a9658;
assign a9664 = a9662 & a9550;
assign a9666 = ~a9662 & ~a9550;
assign a9668 = ~a9666 & ~a9664;
assign a9670 = ~i236 & ~i234;
assign a9672 = ~a9670 & ~a8986;
assign a9674 = a9672 & ~a8980;
assign a9676 = ~a9674 & ~a8884;
assign a9678 = ~a9658 & a9558;
assign a9680 = ~a9658 & ~a8884;
assign a9682 = ~a9680 & a9556;
assign a9684 = ~a9682 & ~a9678;
assign a9686 = a9684 & ~a8898;
assign a9688 = ~a9686 & ~a9676;
assign a9690 = ~a9684 & a8898;
assign a9692 = ~a9690 & ~a9688;
assign a9694 = a9692 & ~a8916;
assign a9696 = ~a9658 & ~a8898;
assign a9698 = ~a9696 & ~a9566;
assign a9700 = a9696 & a9566;
assign a9702 = ~a9700 & ~a9698;
assign a9704 = ~a9702 & ~a9678;
assign a9706 = a9702 & a9678;
assign a9708 = ~a9706 & ~a9704;
assign a9710 = ~a9692 & a8916;
assign a9712 = ~a9710 & a9708;
assign a9714 = ~a9712 & ~a9694;
assign a9716 = ~a9714 & ~a8934;
assign a9718 = ~a9592 & ~a9576;
assign a9720 = a9718 & ~a9658;
assign a9722 = a9720 & a9590;
assign a9724 = ~a9720 & ~a9590;
assign a9726 = ~a9724 & ~a9722;
assign a9728 = a9714 & a8934;
assign a9730 = ~a9728 & a9726;
assign a9732 = ~a9730 & ~a9716;
assign a9734 = ~a9732 & ~a8958;
assign a9736 = ~a9610 & ~a9598;
assign a9738 = a9736 & ~a9658;
assign a9740 = a9738 & a9608;
assign a9742 = ~a9738 & ~a9608;
assign a9744 = ~a9742 & ~a9740;
assign a9746 = a9732 & a8958;
assign a9748 = ~a9746 & a9744;
assign a9750 = ~a9748 & ~a9734;
assign a9752 = a9668 & a8950;
assign a9754 = ~a9752 & a9750;
assign a9756 = ~a9658 & a8950;
assign a9758 = a9756 & a9632;
assign a9760 = ~a9756 & ~a9632;
assign a9762 = ~a9760 & ~a9758;
assign a9764 = ~a9658 & ~a9622;
assign a9766 = ~a9764 & ~a9762;
assign a9768 = a9764 & a9762;
assign a9770 = ~a9668 & ~a8950;
assign a9772 = ~a9770 & ~a9768;
assign a9774 = a9772 & ~a9766;
assign a9776 = a9774 & ~a9754;
assign a9778 = ~a9750 & a8950;
assign a9780 = a9750 & ~a8950;
assign a9782 = ~a9780 & ~a9778;
assign a9784 = a9782 & ~a9776;
assign a9786 = a9784 & a9668;
assign a9788 = ~a9784 & ~a9668;
assign a9790 = ~a9788 & ~a9786;
assign a9792 = ~a9776 & a9676;
assign a9794 = ~a9776 & ~a8884;
assign a9796 = ~a9794 & a9674;
assign a9798 = ~a9796 & ~a9792;
assign a9800 = a9798 & ~a8898;
assign a9802 = ~a9800 & ~a8984;
assign a9804 = ~a9798 & a8898;
assign a9806 = ~a9804 & ~a9802;
assign a9808 = a9806 & ~a8916;
assign a9810 = ~a9776 & ~a8898;
assign a9812 = ~a9810 & ~a9684;
assign a9814 = a9810 & a9684;
assign a9816 = ~a9814 & ~a9812;
assign a9818 = ~a9816 & ~a9792;
assign a9820 = a9816 & a9792;
assign a9822 = ~a9820 & ~a9818;
assign a9824 = ~a9806 & a8916;
assign a9826 = ~a9824 & a9822;
assign a9828 = ~a9826 & ~a9808;
assign a9830 = ~a9828 & ~a8934;
assign a9832 = ~a9710 & ~a9694;
assign a9834 = a9832 & ~a9776;
assign a9836 = a9834 & a9708;
assign a9838 = ~a9834 & ~a9708;
assign a9840 = ~a9838 & ~a9836;
assign a9842 = a9828 & a8934;
assign a9844 = ~a9842 & a9840;
assign a9846 = ~a9844 & ~a9830;
assign a9848 = ~a9846 & ~a8958;
assign a9850 = ~a9728 & ~a9716;
assign a9852 = a9850 & ~a9776;
assign a9854 = a9852 & a9726;
assign a9856 = ~a9852 & ~a9726;
assign a9858 = ~a9856 & ~a9854;
assign a9860 = a9846 & a8958;
assign a9862 = ~a9860 & a9858;
assign a9864 = ~a9862 & ~a9848;
assign a9866 = ~a9864 & a8950;
assign a9868 = a9864 & ~a8950;
assign a9870 = ~a9746 & ~a9734;
assign a9872 = a9870 & ~a9776;
assign a9874 = a9872 & a9744;
assign a9876 = ~a9872 & ~a9744;
assign a9878 = ~a9876 & ~a9874;
assign a9880 = a9878 & ~a9868;
assign a9882 = ~a9880 & ~a9866;
assign a9884 = ~a9882 & a9790;
assign a9886 = ~a9884 & a8984;
assign a9888 = ~a9884 & ~a8884;
assign a9890 = ~a9888 & a8982;
assign a9892 = ~a9890 & ~a9886;
assign a9894 = ~a9884 & ~a8898;
assign a9896 = ~a9894 & ~a9798;
assign a9898 = a9894 & a9798;
assign a9900 = ~a9898 & ~a9896;
assign a9902 = ~a9900 & ~a9886;
assign a9904 = a9900 & a9886;
assign a9906 = ~a9904 & ~a9902;
assign a9908 = ~a9906 & ~a9892;
assign a9910 = ~a9824 & ~a9808;
assign a9912 = a9910 & ~a9884;
assign a9914 = a9912 & a9822;
assign a9916 = ~a9912 & ~a9822;
assign a9918 = ~a9916 & ~a9914;
assign a9920 = ~a9918 & a9908;
assign a9922 = ~a9842 & ~a9830;
assign a9924 = a9922 & ~a9884;
assign a9926 = a9924 & a9840;
assign a9928 = ~a9924 & ~a9840;
assign a9930 = ~a9928 & ~a9926;
assign a9932 = ~a9930 & a9920;
assign a9934 = ~a9860 & ~a9848;
assign a9936 = a9934 & ~a9884;
assign a9938 = a9936 & a9858;
assign a9940 = ~a9936 & ~a9858;
assign a9942 = ~a9940 & ~a9938;
assign a9944 = ~a9942 & a9932;
assign a9946 = ~a9868 & ~a9866;
assign a9948 = a9946 & ~a9884;
assign a9950 = a9948 & a9878;
assign a9952 = ~a9948 & ~a9878;
assign a9954 = ~a9952 & ~a9950;
assign a9956 = ~a9954 & ~a9944;
assign a9958 = a9954 & a9944;
assign a9960 = ~a9958 & ~a9956;
assign a9962 = ~a9960 & ~a8968;
assign a9964 = a9962 & ~a8876;
assign a9966 = a9892 & ~a8968;
assign a9968 = a9966 & a3760;
assign a9970 = a9906 & a9892;
assign a9972 = ~a9970 & ~a9908;
assign a9974 = a9972 & ~a8968;
assign a9976 = a9974 & a4260;
assign a9978 = ~a9976 & ~a9968;
assign a9980 = ~a9974 & ~a4260;
assign a9982 = ~a9980 & ~a9978;
assign a9984 = a9918 & ~a9908;
assign a9986 = ~a9984 & ~a9920;
assign a9988 = a9986 & ~a8968;
assign a9990 = a9988 & a4286;
assign a9992 = ~a9990 & ~a9982;
assign a9994 = ~a9988 & ~a4286;
assign a9996 = ~a9994 & ~a9992;
assign a9998 = a9930 & ~a9920;
assign a10000 = ~a9998 & ~a9932;
assign a10002 = a10000 & ~a8968;
assign a10004 = a10002 & a4312;
assign a10006 = ~a10004 & ~a9996;
assign a10008 = ~a10002 & ~a4312;
assign a10010 = ~a10008 & ~a10006;
assign a10012 = a9942 & ~a9932;
assign a10014 = ~a10012 & ~a9944;
assign a10016 = a10014 & ~a8968;
assign a10018 = a10016 & a3758;
assign a10020 = ~a10018 & ~a10010;
assign a10022 = ~a10016 & ~a3758;
assign a10024 = ~a10022 & ~a10020;
assign a10026 = a10024 & ~a9962;
assign a10028 = ~a10024 & a9962;
assign a10030 = ~a10028 & ~a10026;
assign a10032 = ~a10030 & a4384;
assign a10034 = ~a10032 & ~a4378;
assign a10036 = ~a10034 & a8876;
assign a10038 = ~a10036 & ~a9964;
assign a10040 = a10038 & ~l1686;
assign a10042 = l1686 & l1026;
assign a10044 = ~a10042 & ~a10040;
assign a10046 = ~a8968 & ~a8876;
assign a10048 = a10046 & a10014;
assign a10050 = ~a10022 & a10020;
assign a10052 = ~a10022 & ~a10018;
assign a10054 = ~a10052 & a10010;
assign a10056 = ~a10054 & ~a10050;
assign a10058 = ~a10056 & a4384;
assign a10060 = ~a4384 & a1712;
assign a10062 = a10060 & a3756;
assign a10064 = ~a10062 & ~a10058;
assign a10066 = ~a10064 & a8876;
assign a10068 = ~a10066 & ~a10048;
assign a10070 = a10068 & ~l1686;
assign a10072 = l1686 & l1032;
assign a10074 = ~a10072 & ~a10070;
assign a10076 = a10046 & a10000;
assign a10078 = ~a10008 & a10006;
assign a10080 = ~a10008 & ~a10004;
assign a10082 = ~a10080 & a9996;
assign a10084 = ~a10082 & ~a10078;
assign a10086 = ~a10084 & a4384;
assign a10088 = a10060 & a4310;
assign a10090 = ~a10088 & ~a10086;
assign a10092 = ~a10090 & a8876;
assign a10094 = ~a10092 & ~a10076;
assign a10096 = a10094 & ~l1686;
assign a10098 = l1686 & l1038;
assign a10100 = ~a10098 & ~a10096;
assign a10102 = a10046 & a9986;
assign a10104 = ~a9994 & a9992;
assign a10106 = ~a9994 & ~a9990;
assign a10108 = ~a10106 & a9982;
assign a10110 = ~a10108 & ~a10104;
assign a10112 = ~a10110 & a4384;
assign a10114 = a10060 & a4284;
assign a10116 = ~a10114 & ~a10112;
assign a10118 = ~a10116 & a8876;
assign a10120 = ~a10118 & ~a10102;
assign a10122 = a10120 & ~l1686;
assign a10124 = l1686 & l1044;
assign a10126 = ~a10124 & ~a10122;
assign a10128 = a10046 & a9972;
assign a10130 = ~a9980 & a9978;
assign a10132 = ~a9980 & ~a9976;
assign a10134 = ~a10132 & a9968;
assign a10136 = ~a10134 & ~a10130;
assign a10138 = ~a10136 & a4384;
assign a10140 = a10060 & a4258;
assign a10142 = ~a10140 & ~a10138;
assign a10144 = ~a10142 & a8876;
assign a10146 = ~a10144 & ~a10128;
assign a10148 = a10146 & ~l1686;
assign a10150 = l1686 & l1050;
assign a10152 = ~a10150 & ~a10148;
assign a10154 = a3782 & ~l1686;
assign a10156 = l1686 & l1054;
assign a10158 = ~a10156 & ~a10154;
assign a10160 = a10046 & a9892;
assign a10162 = a9966 & a4384;
assign a10164 = a10162 & a3760;
assign a10166 = ~a10162 & ~a3760;
assign a10168 = ~a10166 & a8876;
assign a10170 = a10168 & ~a10164;
assign a10172 = ~a10170 & ~a10160;
assign a10174 = a10172 & ~l1686;
assign a10176 = l1686 & l1052;
assign a10178 = ~a10176 & ~a10174;
assign a10180 = l1686 & ~l1056;
assign a10182 = a10180 & ~a10178;
assign a10184 = a10182 & a10158;
assign a10186 = a10184 & ~a10152;
assign a10188 = l1686 & ~l1048;
assign a10190 = ~a10180 & ~a10178;
assign a10192 = a10190 & a10158;
assign a10194 = a10192 & ~a10152;
assign a10196 = a10194 & a10188;
assign a10198 = ~a10196 & ~a10186;
assign a10200 = a3884 & ~l1686;
assign a10202 = l1686 & l1046;
assign a10204 = ~a10202 & ~a10200;
assign a10206 = a10182 & ~a10158;
assign a10208 = a10206 & ~a10152;
assign a10210 = a10184 & a10152;
assign a10212 = a10190 & ~a10158;
assign a10214 = ~a10212 & ~a10178;
assign a10216 = ~a10214 & ~a10152;
assign a10218 = ~a10216 & ~a10210;
assign a10220 = ~a10218 & a10188;
assign a10222 = ~a10220 & ~a10208;
assign a10224 = ~a10222 & a10204;
assign a10226 = ~a10224 & a10198;
assign a10228 = ~a10226 & ~a10126;
assign a10230 = l1686 & ~l1042;
assign a10232 = a10194 & ~a10188;
assign a10234 = a10192 & a10152;
assign a10236 = ~a10218 & ~a10188;
assign a10238 = ~a10236 & ~a10234;
assign a10240 = ~a10238 & a10204;
assign a10242 = ~a10240 & ~a10232;
assign a10244 = ~a10242 & ~a10126;
assign a10246 = a10244 & a10230;
assign a10248 = ~a10246 & ~a10228;
assign a10250 = a3958 & ~l1686;
assign a10252 = l1686 & l1040;
assign a10254 = ~a10252 & ~a10250;
assign a10256 = a10206 & a10152;
assign a10258 = a10256 & a10188;
assign a10260 = ~a10222 & ~a10204;
assign a10262 = ~a10260 & ~a10258;
assign a10264 = ~a10262 & ~a10126;
assign a10266 = ~a10226 & a10126;
assign a10268 = a10256 & ~a10188;
assign a10270 = ~a10214 & a10152;
assign a10272 = ~a10270 & ~a10268;
assign a10274 = ~a10238 & ~a10204;
assign a10276 = ~a10274 & a10272;
assign a10278 = ~a10276 & ~a10126;
assign a10280 = ~a10278 & ~a10266;
assign a10282 = ~a10280 & a10230;
assign a10284 = ~a10282 & ~a10264;
assign a10286 = ~a10284 & a10254;
assign a10288 = ~a10286 & a10248;
assign a10290 = ~a10288 & ~a10100;
assign a10292 = l1686 & ~l1036;
assign a10294 = a10244 & ~a10230;
assign a10296 = ~a10242 & a10126;
assign a10298 = ~a10280 & ~a10230;
assign a10300 = ~a10298 & ~a10296;
assign a10302 = ~a10300 & a10254;
assign a10304 = ~a10302 & ~a10294;
assign a10306 = ~a10304 & ~a10100;
assign a10308 = a10306 & a10292;
assign a10310 = ~a10308 & ~a10290;
assign a10312 = a4036 & ~l1686;
assign a10314 = l1686 & l1034;
assign a10316 = ~a10314 & ~a10312;
assign a10318 = ~a10262 & a10126;
assign a10320 = a10318 & a10230;
assign a10322 = ~a10284 & ~a10254;
assign a10324 = ~a10322 & ~a10320;
assign a10326 = ~a10324 & ~a10100;
assign a10328 = ~a10288 & a10100;
assign a10330 = a10318 & ~a10230;
assign a10332 = ~a10276 & a10126;
assign a10334 = ~a10332 & ~a10330;
assign a10336 = ~a10300 & ~a10254;
assign a10338 = ~a10336 & a10334;
assign a10340 = ~a10338 & ~a10100;
assign a10342 = ~a10340 & ~a10328;
assign a10344 = ~a10342 & a10292;
assign a10346 = ~a10344 & ~a10326;
assign a10348 = ~a10346 & a10316;
assign a10350 = ~a10348 & a10310;
assign a10352 = ~a10350 & ~a10074;
assign a10354 = l1686 & ~l1030;
assign a10356 = a10306 & ~a10292;
assign a10358 = ~a10304 & a10100;
assign a10360 = ~a10342 & ~a10292;
assign a10362 = ~a10360 & ~a10358;
assign a10364 = ~a10362 & a10316;
assign a10366 = ~a10364 & ~a10356;
assign a10368 = ~a10366 & ~a10074;
assign a10370 = a10368 & a10354;
assign a10372 = ~a10370 & ~a10352;
assign a10374 = a4114 & ~l1686;
assign a10376 = l1686 & l1028;
assign a10378 = ~a10376 & ~a10374;
assign a10380 = ~a10324 & a10100;
assign a10382 = a10380 & a10292;
assign a10384 = ~a10346 & ~a10316;
assign a10386 = ~a10384 & ~a10382;
assign a10388 = ~a10386 & ~a10074;
assign a10390 = ~a10350 & a10074;
assign a10392 = a10380 & ~a10292;
assign a10394 = ~a10338 & a10100;
assign a10396 = ~a10394 & ~a10392;
assign a10398 = ~a10362 & ~a10316;
assign a10400 = ~a10398 & a10396;
assign a10402 = ~a10400 & ~a10074;
assign a10404 = ~a10402 & ~a10390;
assign a10406 = ~a10404 & a10354;
assign a10408 = ~a10406 & ~a10388;
assign a10410 = ~a10408 & a10378;
assign a10412 = ~a10410 & a10372;
assign a10414 = ~a10412 & ~a10044;
assign a10416 = l1686 & ~l1024;
assign a10418 = a10368 & ~a10354;
assign a10420 = ~a10366 & a10074;
assign a10422 = ~a10404 & ~a10354;
assign a10424 = ~a10422 & ~a10420;
assign a10426 = ~a10424 & a10378;
assign a10428 = ~a10426 & ~a10418;
assign a10430 = ~a10428 & ~a10044;
assign a10432 = a10430 & a10416;
assign a10434 = ~a10432 & ~a10414;
assign a10436 = a4188 & ~l1686;
assign a10438 = l1686 & l1022;
assign a10440 = ~a10438 & ~a10436;
assign a10442 = ~a10386 & a10074;
assign a10444 = a10442 & a10354;
assign a10446 = ~a10408 & ~a10378;
assign a10448 = ~a10446 & ~a10444;
assign a10450 = ~a10448 & ~a10044;
assign a10452 = ~a10412 & a10044;
assign a10454 = a10442 & ~a10354;
assign a10456 = ~a10400 & a10074;
assign a10458 = ~a10456 & ~a10454;
assign a10460 = ~a10424 & ~a10378;
assign a10462 = ~a10460 & a10458;
assign a10464 = ~a10462 & ~a10044;
assign a10466 = ~a10464 & ~a10452;
assign a10468 = ~a10466 & a10416;
assign a10470 = ~a10468 & ~a10450;
assign a10472 = ~a10470 & a10440;
assign a10474 = ~a10472 & a10434;
assign a10476 = ~a10474 & ~a8874;
assign a10478 = l1686 & ~l1018;
assign a10480 = a10430 & ~a10416;
assign a10482 = ~a10428 & a10044;
assign a10484 = ~a10466 & ~a10416;
assign a10486 = ~a10484 & ~a10482;
assign a10488 = ~a10486 & a10440;
assign a10490 = ~a10488 & ~a10480;
assign a10492 = ~a10490 & ~a8874;
assign a10494 = a10492 & a10478;
assign a10496 = ~a10494 & ~a10476;
assign a10498 = l1686 & ~l1016;
assign a10500 = ~a10448 & a10044;
assign a10502 = a10500 & a10416;
assign a10504 = ~a10470 & ~a10440;
assign a10506 = ~a10504 & ~a10502;
assign a10508 = ~a10506 & ~a8874;
assign a10510 = ~a10474 & a8874;
assign a10512 = a10500 & ~a10416;
assign a10514 = ~a10462 & a10044;
assign a10516 = ~a10514 & ~a10512;
assign a10518 = ~a10486 & ~a10440;
assign a10520 = ~a10518 & a10516;
assign a10522 = ~a10520 & ~a8874;
assign a10524 = ~a10522 & ~a10510;
assign a10526 = ~a10524 & a10478;
assign a10528 = ~a10526 & ~a10508;
assign a10530 = ~a10528 & a10498;
assign a10532 = ~a10530 & a10496;
assign a10534 = ~a10532 & ~a8872;
assign a10536 = a10492 & ~a10478;
assign a10538 = ~a10490 & a8874;
assign a10540 = ~a10524 & ~a10478;
assign a10542 = ~a10540 & ~a10538;
assign a10544 = ~a10542 & a10498;
assign a10546 = ~a10544 & ~a10536;
assign a10548 = ~a10546 & a8872;
assign a10550 = ~a10548 & ~a10534;
assign a10552 = ~a10550 & a8870;
assign a10554 = ~a10506 & a8874;
assign a10556 = a10554 & a10478;
assign a10558 = ~a10528 & ~a10498;
assign a10560 = ~a10558 & ~a10556;
assign a10562 = ~a10560 & ~a8872;
assign a10564 = a10554 & ~a10478;
assign a10566 = ~a10520 & a8874;
assign a10568 = ~a10566 & ~a10564;
assign a10570 = ~a10542 & ~a10498;
assign a10572 = ~a10570 & a10568;
assign a10574 = ~a10572 & a8872;
assign a10576 = ~a10574 & ~a10562;
assign a10578 = ~a10576 & ~a8870;
assign a10580 = ~a10578 & ~a10552;
assign a10582 = ~a10580 & ~a8868;
assign a10584 = ~a10532 & a8872;
assign a10586 = ~a10546 & ~a8872;
assign a10588 = ~a10586 & ~a10584;
assign a10590 = ~a10588 & ~a8870;
assign a10592 = ~a10560 & a8872;
assign a10594 = ~a10572 & ~a8872;
assign a10596 = ~a10594 & ~a10592;
assign a10598 = ~a10596 & a8870;
assign a10600 = ~a10598 & ~a10590;
assign a10602 = ~a10600 & a8868;
assign a10604 = ~a10602 & ~a10582;
assign a10606 = a10588 & a10576;
assign a10608 = a10606 & ~a8870;
assign a10610 = ~a10606 & a8870;
assign a10612 = ~a10610 & ~a10608;
assign a10614 = a10612 & a10604;
assign a10616 = ~a10614 & a8866;
assign a10618 = a10616 & a8864;
assign a10620 = a10618 & ~a8050;
assign a10622 = a10620 & ~a8862;
assign a10624 = a10622 & ~a8054;
assign a10626 = a10624 & a8860;
assign a10628 = a10620 & a8862;
assign a10630 = ~a10614 & ~a8866;
assign a10632 = a10630 & a8864;
assign a10634 = a10632 & ~a8050;
assign a10636 = ~a10634 & ~a10628;
assign a10638 = ~a10636 & ~a8054;
assign a10640 = ~a10638 & ~a10626;
assign a10642 = ~a10640 & ~a8052;
assign a10644 = a10630 & ~a8864;
assign a10646 = ~a10644 & ~a10618;
assign a10648 = ~a10646 & a8050;
assign a10650 = a10648 & a8862;
assign a10652 = a10644 & ~a8050;
assign a10654 = a10652 & ~a8862;
assign a10656 = ~a10654 & ~a10650;
assign a10658 = a10656 & ~a10622;
assign a10660 = ~a10658 & a8054;
assign a10662 = a10660 & ~a8860;
assign a10664 = ~a10662 & ~a10642;
assign a10666 = a10616 & ~a8864;
assign a10668 = a10632 & a8050;
assign a10670 = ~a10668 & ~a10666;
assign a10672 = a10652 & a8862;
assign a10674 = ~a10672 & a10670;
assign a10676 = a10648 & ~a8862;
assign a10678 = ~a10676 & a10674;
assign a10680 = ~a10636 & a8054;
assign a10682 = ~a10680 & a10678;
assign a10684 = ~a10656 & ~a8054;
assign a10686 = a10684 & a8860;
assign a10688 = ~a10686 & a10682;
assign a10690 = a10688 & a10664;
assign a10692 = a10660 & a8860;
assign a10694 = a10684 & ~a8860;
assign a10696 = ~a10694 & ~a10692;
assign a10698 = ~a8850 & a8228;
assign a10700 = ~a10698 & ~a8852;
assign a10702 = ~a10700 & ~l1686;
assign a10704 = l1686 & l1062;
assign a10706 = ~a10704 & ~a10702;
assign a10708 = ~a10706 & a8052;
assign a10710 = a10708 & ~a10696;
assign a10712 = ~a10710 & a10690;
assign a10714 = a10706 & ~a8052;
assign a10716 = a10624 & ~a8860;
assign a10718 = ~a10716 & a10696;
assign a10720 = ~a10718 & a10714;
assign a10722 = ~a10720 & a10712;
assign a10724 = ~a10722 & ~a8072;
assign a10726 = ~a10580 & a8868;
assign a10728 = ~a10600 & ~a8868;
assign a10730 = ~a10718 & ~a10714;
assign a10732 = a10730 & ~a10708;
assign a10734 = ~a10732 & ~a10728;
assign a10736 = a10734 & ~a10726;
assign a10738 = a10736 & ~a10724;
assign a10740 = a10716 & ~a10706;
assign a10742 = ~a10740 & a10640;
assign a10744 = ~a10742 & a8052;
assign a10746 = ~a10744 & a10738;
assign a10748 = a10746 & i218;
assign a10750 = a10748 & a8056;
assign a10752 = ~a10750 & a8050;
assign a10754 = a10750 & ~a8050;
assign a10756 = ~a10754 & ~a10752;
assign a10758 = ~a10756 & a8048;
assign a10760 = l1686 & ~l1070;
assign a10762 = a10760 & ~a8048;
assign a10764 = ~a10762 & ~a10758;
assign a10766 = ~a4388 & a4384;
assign a10768 = a10766 & i212;
assign a10770 = a10768 & ~l1686;
assign a10772 = l1686 & l986;
assign a10774 = ~a10772 & ~a10770;
assign a10776 = l1686 & l980;
assign a10778 = ~a10776 & ~a10770;
assign a10780 = l1686 & l982;
assign a10782 = ~a10780 & ~a10770;
assign a10784 = ~a10782 & ~a10778;
assign a10786 = a10784 & ~a10774;
assign a10788 = ~a10786 & ~a10764;
assign a10790 = l1686 & ~l1068;
assign a10792 = a10790 & a10786;
assign a10794 = ~a10792 & ~a10788;
assign a10796 = ~a10794 & ~l972;
assign a10798 = ~a10796 & ~a8046;
assign a10800 = a10782 & a10778;
assign a10802 = a10800 & l984;
assign a10804 = ~a10802 & ~a10798;
assign a10806 = a10802 & a10790;
assign a10808 = ~a10806 & ~a10804;
assign a10810 = ~a10808 & ~l972;
assign a10812 = ~a10810 & ~a8046;
assign a10814 = ~a10812 & ~l494;
assign a10818 = ~a6476 & l972;
assign a10820 = a10744 & ~a8072;
assign a10822 = ~a10820 & a10722;
assign a10824 = a10822 & a10736;
assign a10826 = a10824 & i272;
assign a10828 = ~a10826 & ~a10748;
assign a10830 = a10828 & a8864;
assign a10832 = a8056 & a8050;
assign a10834 = a10832 & ~a8864;
assign a10836 = ~a10832 & a8864;
assign a10838 = ~a10836 & ~a10834;
assign a10840 = ~a10838 & a10748;
assign a10842 = ~a10840 & ~a10830;
assign a10844 = ~a10842 & a8048;
assign a10846 = l1686 & ~l1000;
assign a10848 = a10846 & ~a8048;
assign a10850 = ~a10848 & ~a10844;
assign a10852 = ~a10850 & ~a10786;
assign a10854 = l1686 & ~l996;
assign a10856 = a10854 & a10786;
assign a10858 = ~a10856 & ~a10852;
assign a10860 = ~a10858 & ~l972;
assign a10862 = ~a10860 & ~a10818;
assign a10864 = ~a10862 & ~a10802;
assign a10866 = a10854 & a10802;
assign a10868 = ~a10866 & ~a10864;
assign a10870 = ~a10868 & ~l972;
assign a10872 = ~a10870 & ~a10818;
assign a10874 = ~a10872 & ~l494;
assign a10878 = ~a10876 & a10816;
assign a10880 = ~a6512 & l972;
assign a10882 = a10828 & a8052;
assign a10884 = a10748 & ~a8052;
assign a10886 = ~a10884 & ~a10882;
assign a10888 = ~a10886 & a8048;
assign a10890 = l1686 & ~l1078;
assign a10892 = a10890 & ~a8048;
assign a10894 = ~a10892 & ~a10888;
assign a10896 = ~a10894 & ~a10786;
assign a10898 = l1686 & ~l1076;
assign a10900 = a10898 & a10786;
assign a10902 = ~a10900 & ~a10896;
assign a10904 = ~a10902 & ~l972;
assign a10906 = ~a10904 & ~a10880;
assign a10908 = ~a10906 & ~a10802;
assign a10910 = a10898 & a10802;
assign a10912 = ~a10910 & ~a10908;
assign a10914 = ~a10912 & ~l972;
assign a10916 = ~a10914 & ~a10880;
assign a10918 = ~a10916 & ~l494;
assign a10922 = ~a6548 & l972;
assign a10924 = a10748 & a8052;
assign a10926 = ~a10924 & ~a8054;
assign a10928 = ~a10926 & ~a10750;
assign a10930 = a10928 & a8048;
assign a10932 = l1686 & ~l1074;
assign a10934 = a10932 & ~a8048;
assign a10936 = ~a10934 & ~a10930;
assign a10938 = ~a10936 & ~a10786;
assign a10940 = l1686 & ~l1072;
assign a10942 = a10940 & a10786;
assign a10944 = ~a10942 & ~a10938;
assign a10946 = ~a10944 & ~l972;
assign a10948 = ~a10946 & ~a10922;
assign a10950 = ~a10948 & ~a10802;
assign a10952 = a10940 & a10802;
assign a10954 = ~a10952 & ~a10950;
assign a10956 = ~a10954 & ~l972;
assign a10958 = ~a10956 & ~a10922;
assign a10960 = ~a10958 & ~l494;
assign a10964 = a10962 & ~a10920;
assign a10966 = a10964 & a10878;
assign a10968 = a10966 & ~a5542;
assign a10970 = ~a10920 & ~a5542;
assign a10972 = a10920 & ~a5548;
assign a10974 = ~a10972 & ~a10970;
assign a10976 = ~a10962 & a10920;
assign a10978 = ~a10976 & ~a10964;
assign a10980 = a10978 & ~a10974;
assign a10982 = a10964 & ~a5556;
assign a10984 = a10976 & ~a5572;
assign a10986 = ~a10984 & ~a10982;
assign a10988 = a10986 & ~a10980;
assign a10990 = ~a10962 & ~a10920;
assign a10992 = ~a10990 & a10816;
assign a10994 = a10990 & ~a10816;
assign a10996 = ~a10994 & ~a10992;
assign a10998 = ~a10996 & ~a10988;
assign a11000 = ~a10920 & l576;
assign a11002 = a10920 & l578;
assign a11004 = ~a11002 & ~a11000;
assign a11006 = ~a11004 & a10978;
assign a11008 = a10964 & l580;
assign a11010 = a10976 & l582;
assign a11012 = ~a11010 & ~a11008;
assign a11014 = a11012 & ~a11006;
assign a11016 = ~a11014 & a10996;
assign a11018 = ~a11016 & ~a10998;
assign a11020 = a10994 & a10876;
assign a11022 = ~a10994 & ~a10876;
assign a11024 = ~a11022 & ~a11020;
assign a11026 = a11024 & ~a11018;
assign a11028 = ~a10920 & l586;
assign a11030 = a10920 & l584;
assign a11032 = ~a11030 & ~a11028;
assign a11034 = ~a11032 & ~a11024;
assign a11036 = ~a11034 & ~a11026;
assign a11038 = ~a11036 & ~a10966;
assign a11042 = a6522 & a5580;
assign a11044 = a6566 & a6522;
assign a11046 = a11044 & a6608;
assign a11048 = a11046 & a6494;
assign a11050 = ~a11048 & ~a5580;
assign a11052 = ~a11050 & ~a11042;
assign a11054 = a11050 & a6522;
assign a11056 = ~a11054 & ~a11052;
assign a11058 = a11056 & ~a10920;
assign a11060 = ~a11056 & a10920;
assign a11062 = ~a11054 & ~a6566;
assign a11064 = a11054 & a6566;
assign a11066 = ~a11064 & ~a11062;
assign a11068 = a11066 & ~a10962;
assign a11070 = ~a11066 & a10962;
assign a11072 = ~a11064 & ~a6608;
assign a11074 = a11064 & a6608;
assign a11076 = ~a11074 & ~a11072;
assign a11078 = a11076 & ~a10816;
assign a11080 = ~a11076 & a10816;
assign a11082 = a11046 & ~a5580;
assign a11084 = ~a11082 & ~a6494;
assign a11086 = a11082 & a6494;
assign a11088 = ~a11086 & ~a11084;
assign a11090 = ~a11088 & a10876;
assign a11092 = a11088 & ~a10876;
assign a11094 = ~a11092 & ~a11090;
assign a11096 = a11094 & ~a11080;
assign a11098 = a11096 & ~a11078;
assign a11100 = a11098 & ~a11070;
assign a11102 = a11100 & ~a11068;
assign a11104 = a11102 & ~a11060;
assign a11106 = a11104 & ~a11058;
assign a11108 = ~a11106 & ~a11040;
assign a11110 = l1686 & ~l1472;
assign a11112 = ~a6710 & ~a1690;
assign a11114 = a11112 & ~a11110;
assign a11116 = a11114 & a11108;
assign a11118 = ~a5098 & ~a4674;
assign a11120 = a4672 & ~a4500;
assign a11122 = ~a11120 & ~a11118;
assign a11124 = ~a4690 & a4464;
assign a11126 = ~a11124 & ~a11122;
assign a11128 = a4690 & ~a4464;
assign a11130 = ~a11128 & ~a11126;
assign a11132 = ~a4706 & a4428;
assign a11134 = ~a11132 & ~a11130;
assign a11136 = a4706 & ~a4428;
assign a11138 = ~a11136 & ~a11134;
assign a11140 = ~a4722 & a2566;
assign a11142 = ~a11140 & ~a11138;
assign a11144 = a4722 & ~a2566;
assign a11146 = ~a11144 & ~a11142;
assign a11148 = ~a4738 & a4404;
assign a11150 = ~a11148 & ~a11146;
assign a11152 = ~a11150 & ~a4926;
assign a11154 = ~a11152 & ~a4770;
assign a11156 = ~a11154 & a4802;
assign a11158 = a4656 & ~a4536;
assign a11160 = ~a11158 & ~a11120;
assign a11162 = ~a11160 & ~a4674;
assign a11164 = ~a11162 & ~a11128;
assign a11166 = ~a11164 & ~a11124;
assign a11168 = ~a11166 & ~a11136;
assign a11170 = ~a11168 & ~a11132;
assign a11172 = ~a11170 & ~a11144;
assign a11174 = ~a11172 & ~a11140;
assign a11176 = ~a11174 & ~a4926;
assign a11178 = ~a11176 & ~a11148;
assign a11180 = ~a11178 & ~a4754;
assign a11182 = ~a11180 & a4778;
assign a11184 = ~a11182 & ~a11156;
assign a11186 = ~a5580 & ~l494;
assign a11188 = a11186 & ~a11184;
assign a11190 = ~a11188 & a4760;
assign a11192 = a11188 & ~a2268;
assign a11194 = ~a11192 & ~a11190;
assign a11196 = ~a11194 & ~a11116;
assign a11198 = ~a10996 & a10978;
assign a11200 = a11198 & ~a11024;
assign a11202 = l1686 & ~l1132;
assign a11204 = a11202 & ~a10920;
assign a11206 = l1686 & ~l1130;
assign a11208 = a11206 & a10920;
assign a11210 = ~a11208 & ~a11204;
assign a11212 = ~a11210 & a11200;
assign a11214 = l1686 & ~l1148;
assign a11216 = a11214 & a10966;
assign a11218 = ~a11216 & ~a11212;
assign a11220 = a11214 & ~a10920;
assign a11222 = l1686 & ~l1146;
assign a11224 = a11222 & a10920;
assign a11226 = ~a11224 & ~a11220;
assign a11228 = ~a11226 & a10978;
assign a11230 = l1686 & ~l1144;
assign a11232 = a11230 & ~a10920;
assign a11234 = l1686 & ~l1142;
assign a11236 = a11234 & a10920;
assign a11238 = ~a11236 & ~a11232;
assign a11240 = ~a11238 & ~a10978;
assign a11242 = ~a11240 & ~a11228;
assign a11244 = ~a11242 & ~a10996;
assign a11246 = l1686 & ~l1140;
assign a11248 = a11246 & ~a10920;
assign a11250 = l1686 & ~l1138;
assign a11252 = a11250 & a10920;
assign a11254 = ~a11252 & ~a11248;
assign a11256 = ~a11254 & a10978;
assign a11258 = l1686 & ~l1136;
assign a11260 = a11258 & ~a10920;
assign a11262 = l1686 & ~l1134;
assign a11264 = a11262 & a10920;
assign a11266 = ~a11264 & ~a11260;
assign a11268 = ~a11266 & ~a10978;
assign a11270 = ~a11268 & ~a11256;
assign a11272 = ~a11270 & a10996;
assign a11274 = ~a11272 & ~a11244;
assign a11276 = ~a11274 & a11024;
assign a11280 = ~a11278 & a11116;
assign a11282 = ~a11280 & ~a11196;
assign a11284 = ~a11188 & a4656;
assign a11286 = a11188 & a4536;
assign a11288 = ~a11286 & ~a11284;
assign a11290 = ~a11288 & ~a11116;
assign a11292 = l1686 & ~l1174;
assign a11294 = a11292 & ~a10920;
assign a11296 = l1686 & ~l1172;
assign a11298 = a11296 & a10920;
assign a11300 = ~a11298 & ~a11294;
assign a11302 = ~a11300 & a11200;
assign a11304 = l1686 & ~l1190;
assign a11306 = a11304 & a10966;
assign a11308 = ~a11306 & ~a11302;
assign a11310 = a11304 & ~a10920;
assign a11312 = a8268 & ~l1686;
assign a11314 = l1686 & l1188;
assign a11316 = ~a11314 & ~a11312;
assign a11318 = a11316 & a10920;
assign a11320 = ~a11318 & ~a11310;
assign a11322 = ~a11320 & a10978;
assign a11324 = a8256 & ~l1686;
assign a11326 = l1686 & l1186;
assign a11328 = ~a11326 & ~a11324;
assign a11330 = a11328 & ~a10920;
assign a11332 = ~a8246 & ~l1686;
assign a11334 = l1686 & l1184;
assign a11336 = ~a11334 & ~a11332;
assign a11338 = a11336 & a10920;
assign a11340 = ~a11338 & ~a11330;
assign a11342 = ~a11340 & ~a10978;
assign a11344 = ~a11342 & ~a11322;
assign a11346 = ~a11344 & ~a10996;
assign a11348 = l1686 & ~l1182;
assign a11350 = a11348 & ~a10920;
assign a11352 = l1686 & ~l1180;
assign a11354 = a11352 & a10920;
assign a11356 = ~a11354 & ~a11350;
assign a11358 = ~a11356 & a10978;
assign a11360 = l1686 & ~l1178;
assign a11362 = a11360 & ~a10920;
assign a11364 = l1686 & ~l1176;
assign a11366 = a11364 & a10920;
assign a11368 = ~a11366 & ~a11362;
assign a11370 = ~a11368 & ~a10978;
assign a11372 = ~a11370 & ~a11358;
assign a11374 = ~a11372 & a10996;
assign a11376 = ~a11374 & ~a11346;
assign a11378 = ~a11376 & a11024;
assign a11382 = ~a11380 & a11116;
assign a11384 = ~a11382 & ~a11290;
assign a11386 = a10774 & ~l984;
assign a11388 = a11386 & a10800;
assign a11390 = ~l964 & ~l962;
assign a11392 = a4390 & ~l1686;
assign a11394 = l1686 & l978;
assign a11396 = ~a11394 & ~a11392;
assign a11398 = a11396 & ~l508;
assign a11400 = a11398 & ~l976;
assign a11402 = a11400 & ~l974;
assign a11404 = a11402 & ~l972;
assign a11406 = a11404 & ~l970;
assign a11408 = a11406 & ~l968;
assign a11410 = a11408 & ~l510;
assign a11412 = a11410 & ~l514;
assign a11414 = a11412 & ~l966;
assign a11416 = a11414 & a11390;
assign a11418 = a11416 & a11388;
assign a11420 = a11418 & i334;
assign a11422 = ~a4384 & ~l1686;
assign a11424 = l1686 & l1460;
assign a11426 = ~a11424 & ~a11422;
assign a11428 = ~a8878 & ~l1686;
assign a11430 = l1686 & l1458;
assign a11432 = ~a11430 & ~a11428;
assign a11434 = ~a11432 & a10178;
assign a11436 = a11432 & ~a10178;
assign a11438 = ~a8886 & ~l1686;
assign a11440 = l1686 & l1456;
assign a11442 = ~a11440 & ~a11438;
assign a11444 = ~a11442 & a10152;
assign a11446 = a11442 & ~a10152;
assign a11448 = ~a8904 & ~l1686;
assign a11450 = l1686 & l1454;
assign a11452 = ~a11450 & ~a11448;
assign a11454 = ~a11452 & a10126;
assign a11456 = a11452 & ~a10126;
assign a11458 = ~a8922 & ~l1686;
assign a11460 = l1686 & l1452;
assign a11462 = ~a11460 & ~a11458;
assign a11464 = ~a11462 & a10100;
assign a11466 = a11462 & ~a10100;
assign a11468 = ~a8936 & ~l1686;
assign a11470 = l1686 & l1450;
assign a11472 = ~a11470 & ~a11468;
assign a11474 = ~a11472 & a10074;
assign a11476 = a11472 & ~a10074;
assign a11478 = l1686 & ~l1448;
assign a11480 = ~a11478 & a10044;
assign a11482 = a11478 & ~a10044;
assign a11484 = a8874 & l1446;
assign a11486 = l1686 & ~l1446;
assign a11488 = a11486 & l1020;
assign a11490 = l1686 & ~l1444;
assign a11492 = a11490 & l992;
assign a11494 = a8868 & l1444;
assign a11496 = ~a11494 & ~a11492;
assign a11498 = a11496 & ~a11488;
assign a11500 = a11498 & ~a11484;
assign a11502 = a11500 & ~a11482;
assign a11504 = a11502 & ~a11480;
assign a11506 = a11504 & ~a11476;
assign a11508 = a11506 & ~a11474;
assign a11510 = a11508 & ~a11466;
assign a11512 = a11510 & ~a11464;
assign a11514 = a11512 & ~a11456;
assign a11516 = a11514 & ~a11454;
assign a11518 = a11516 & ~a11446;
assign a11520 = a11518 & ~a11444;
assign a11522 = a11520 & ~a11436;
assign a11524 = a11522 & ~a11434;
assign a11526 = a11524 & a11426;
assign a11528 = ~a11188 & a4672;
assign a11530 = a11188 & a4500;
assign a11532 = ~a11530 & ~a11528;
assign a11534 = ~a11532 & ~a8062;
assign a11536 = a10204 & a8062;
assign a11538 = ~a11536 & ~a11534;
assign a11540 = ~a11288 & ~a8062;
assign a11542 = a10158 & a8062;
assign a11544 = ~a11542 & ~a11540;
assign a11546 = a11544 & a11538;
assign a11548 = ~a11188 & a4690;
assign a11550 = a11188 & a4464;
assign a11552 = ~a11550 & ~a11548;
assign a11554 = ~a11552 & ~a8062;
assign a11556 = a10254 & a8062;
assign a11558 = ~a11556 & ~a11554;
assign a11560 = a11558 & a11546;
assign a11562 = ~a11188 & a4706;
assign a11564 = a11188 & a4428;
assign a11566 = ~a11564 & ~a11562;
assign a11568 = ~a11566 & ~a8062;
assign a11570 = a10316 & a8062;
assign a11572 = ~a11570 & ~a11568;
assign a11574 = a11572 & a11560;
assign a11576 = ~a11188 & a4722;
assign a11578 = a11188 & a2566;
assign a11580 = ~a11578 & ~a11576;
assign a11582 = ~a11580 & ~a8062;
assign a11584 = a10378 & a8062;
assign a11586 = ~a11584 & ~a11582;
assign a11588 = a11586 & a11574;
assign a11590 = ~a11188 & a4738;
assign a11592 = a11188 & a4404;
assign a11594 = ~a11592 & ~a11590;
assign a11596 = ~a11594 & ~a8062;
assign a11598 = a10440 & a8062;
assign a11600 = ~a11598 & ~a11596;
assign a11602 = a11600 & a11588;
assign a11604 = ~a11188 & a4752;
assign a11606 = a11188 & a2548;
assign a11608 = ~a11606 & ~a11604;
assign a11610 = ~a11608 & ~a8062;
assign a11612 = a10498 & a8062;
assign a11614 = ~a11612 & ~a11610;
assign a11616 = ~a11614 & ~a11602;
assign a11618 = a11614 & a11602;
assign a11620 = ~a11618 & ~a11616;
assign a11622 = l1686 & ~l1082;
assign a11624 = l1686 & ~l1090;
assign a11626 = ~a8222 & ~l1686;
assign a11628 = l1686 & l1092;
assign a11630 = ~a11628 & ~a11626;
assign a11632 = i274 & i24;
assign a11634 = ~a4384 & i276;
assign a11636 = ~a11634 & ~a8904;
assign a11638 = ~a11636 & ~i24;
assign a11640 = ~a11638 & ~a11632;
assign a11642 = ~a11640 & ~a4004;
assign a11644 = i278 & i24;
assign a11646 = ~a4384 & i280;
assign a11648 = ~a11646 & ~a8936;
assign a11650 = ~a11648 & ~i24;
assign a11652 = ~a11650 & ~a11644;
assign a11654 = ~a11652 & ~a4160;
assign a11656 = ~a11654 & ~a11642;
assign a11658 = i282 & i24;
assign a11660 = ~a4384 & i284;
assign a11662 = ~a11660 & ~a8922;
assign a11664 = ~a11662 & ~i24;
assign a11666 = ~a11664 & ~a11658;
assign a11668 = ~a11666 & ~a4082;
assign a11670 = i286 & i24;
assign a11672 = ~a4384 & i288;
assign a11674 = ~a11672 & ~a8886;
assign a11676 = ~a11674 & ~i24;
assign a11678 = ~a11676 & ~a11670;
assign a11680 = a11678 & a3926;
assign a11682 = ~a11680 & ~a11668;
assign a11684 = a11682 & a11656;
assign a11686 = i290 & i24;
assign a11688 = ~a4384 & i292;
assign a11690 = ~a11688 & ~a8878;
assign a11692 = ~a11690 & ~i24;
assign a11694 = ~a11692 & ~a11686;
assign a11696 = a11694 & a3860;
assign a11698 = ~a11678 & ~a3926;
assign a11700 = a4384 & a3838;
assign a11702 = ~i298 & ~i296;
assign a11704 = a11702 & ~i294;
assign a11706 = ~a11704 & i24;
assign a11708 = ~a11706 & a11700;
assign a11710 = a11708 & ~a11698;
assign a11712 = a11710 & ~a11696;
assign a11714 = a11666 & a4082;
assign a11716 = a11640 & a4004;
assign a11718 = ~a11716 & ~a11714;
assign a11720 = ~a11694 & ~a3860;
assign a11722 = a11652 & a4160;
assign a11724 = ~a11722 & ~a11720;
assign a11726 = a11724 & a11718;
assign a11728 = a11726 & a11712;
assign a11730 = a11728 & a11684;
assign a11732 = a8302 & ~a8228;
assign a11734 = a8302 & a8228;
assign a11736 = ~a11734 & ~a3838;
assign a11738 = a11736 & ~a11732;
assign a11740 = ~a11738 & ~a11730;
assign a11742 = ~a11740 & a8224;
assign a11744 = ~a11742 & ~a8226;
assign a11746 = a11744 & ~l1686;
assign a11748 = l1686 & l1084;
assign a11750 = ~a11748 & ~a11746;
assign a11752 = l1686 & ~l1442;
assign a11754 = a11752 & ~a11750;
assign a11756 = l1686 & ~l1440;
assign a11758 = a11756 & a11750;
assign a11760 = ~a11758 & ~a11754;
assign a11762 = ~a11760 & ~a11630;
assign a11764 = a8510 & ~l1686;
assign a11766 = l1686 & l1438;
assign a11768 = ~a11766 & ~a11764;
assign a11770 = a11768 & ~a11750;
assign a11772 = ~a8502 & ~l1686;
assign a11774 = l1686 & l1436;
assign a11776 = ~a11774 & ~a11772;
assign a11778 = a11776 & a11750;
assign a11780 = ~a11778 & ~a11770;
assign a11782 = ~a11780 & a11630;
assign a11784 = ~a11782 & ~a11762;
assign a11786 = ~a11784 & ~a11624;
assign a11788 = l1686 & ~l1434;
assign a11790 = a11788 & ~a11750;
assign a11792 = l1686 & ~l1432;
assign a11794 = a11792 & a11750;
assign a11796 = ~a11794 & ~a11790;
assign a11798 = ~a11796 & ~a11630;
assign a11800 = l1686 & ~l1430;
assign a11802 = a11800 & ~a11750;
assign a11804 = l1686 & ~l1428;
assign a11806 = a11804 & a11750;
assign a11808 = ~a11806 & ~a11802;
assign a11810 = ~a11808 & a11630;
assign a11812 = ~a11810 & ~a11798;
assign a11814 = ~a11812 & a11624;
assign a11816 = ~a11814 & ~a11786;
assign a11818 = ~a11816 & ~a11622;
assign a11820 = l1686 & ~l1426;
assign a11822 = a11820 & ~a11750;
assign a11824 = l1686 & ~l1424;
assign a11826 = a11824 & a11750;
assign a11828 = ~a11826 & ~a11822;
assign a11830 = a11622 & l1090;
assign a11832 = a11830 & ~a11630;
assign a11834 = a11832 & ~a11828;
assign a11836 = ~a11834 & ~a11818;
assign a11838 = ~a11736 & ~l1686;
assign a11840 = l1686 & l1108;
assign a11842 = ~a11840 & ~a11838;
assign a11844 = ~a11842 & ~a11750;
assign a11846 = a11732 & ~l1686;
assign a11848 = l1686 & l1106;
assign a11850 = ~a11848 & ~a11846;
assign a11852 = ~a11850 & a11750;
assign a11854 = ~a11852 & ~a11844;
assign a11856 = ~a11854 & ~a11630;
assign a11858 = ~a11750 & l1104;
assign a11860 = a11750 & l1102;
assign a11862 = ~a11860 & ~a11858;
assign a11864 = ~a11862 & a11630;
assign a11866 = ~a11864 & ~a11856;
assign a11868 = ~a11866 & ~a11624;
assign a11870 = ~a11750 & l1100;
assign a11872 = a11750 & l1098;
assign a11874 = ~a11872 & ~a11870;
assign a11876 = ~a11874 & ~a11630;
assign a11878 = ~a11750 & l1096;
assign a11880 = a11750 & l1094;
assign a11882 = ~a11880 & ~a11878;
assign a11884 = ~a11882 & a11630;
assign a11886 = ~a11884 & ~a11876;
assign a11888 = ~a11886 & a11624;
assign a11890 = ~a11888 & ~a11868;
assign a11892 = ~a11890 & ~a11622;
assign a11894 = ~a11750 & l1088;
assign a11896 = a11750 & l1086;
assign a11898 = ~a11896 & ~a11894;
assign a11900 = ~a11898 & a11622;
assign a11902 = ~a11900 & ~a11892;
assign a11904 = a11902 & ~a11836;
assign a11906 = l1686 & ~l1422;
assign a11908 = a11906 & ~a11750;
assign a11910 = l1686 & ~l1420;
assign a11912 = a11910 & a11750;
assign a11914 = ~a11912 & ~a11908;
assign a11916 = ~a11914 & ~a11630;
assign a11918 = l1686 & ~l1418;
assign a11920 = a11918 & ~a11750;
assign a11922 = l1686 & ~l1416;
assign a11924 = a11922 & a11750;
assign a11926 = ~a11924 & ~a11920;
assign a11928 = ~a11926 & a11630;
assign a11930 = ~a11928 & ~a11916;
assign a11932 = ~a11930 & ~a11624;
assign a11934 = l1686 & ~l1414;
assign a11936 = a11934 & ~a11750;
assign a11938 = l1686 & ~l1412;
assign a11940 = a11938 & a11750;
assign a11942 = ~a11940 & ~a11936;
assign a11944 = ~a11942 & ~a11630;
assign a11946 = l1686 & ~l1410;
assign a11948 = a11946 & ~a11750;
assign a11950 = l1686 & ~l1408;
assign a11952 = a11950 & a11750;
assign a11954 = ~a11952 & ~a11948;
assign a11956 = ~a11954 & a11630;
assign a11958 = ~a11956 & ~a11944;
assign a11960 = ~a11958 & a11624;
assign a11962 = ~a11960 & ~a11932;
assign a11964 = ~a11962 & ~a11622;
assign a11966 = l1686 & ~l1406;
assign a11968 = a11966 & ~a11750;
assign a11970 = l1686 & ~l1404;
assign a11972 = a11970 & a11750;
assign a11974 = ~a11972 & ~a11968;
assign a11976 = ~a11974 & a11832;
assign a11978 = ~a11976 & ~a11964;
assign a11980 = ~a11978 & ~a11902;
assign a11982 = ~a11980 & ~a11904;
assign a11984 = l1686 & l1080;
assign a11986 = ~a11984 & ~a5538;
assign a11988 = ~a11986 & a11902;
assign a11990 = a11988 & a11106;
assign a11992 = ~a11990 & ~a11982;
assign a11994 = a8842 & ~l1686;
assign a11996 = l1686 & l1402;
assign a11998 = ~a11996 & ~a11994;
assign a12000 = a11998 & a11990;
assign a12002 = ~a12000 & ~a11992;
assign a12004 = ~a12002 & a11614;
assign a12006 = a12002 & ~a11614;
assign a12008 = l1686 & ~l1400;
assign a12010 = a12008 & ~a11750;
assign a12012 = a8478 & ~l1686;
assign a12014 = l1686 & l1398;
assign a12016 = ~a12014 & ~a12012;
assign a12018 = a12016 & a11750;
assign a12020 = ~a12018 & ~a12010;
assign a12022 = ~a12020 & ~a11630;
assign a12024 = a8468 & ~l1686;
assign a12026 = l1686 & l1396;
assign a12028 = ~a12026 & ~a12024;
assign a12030 = a12028 & ~a11750;
assign a12032 = ~a8462 & ~l1686;
assign a12034 = l1686 & l1394;
assign a12036 = ~a12034 & ~a12032;
assign a12038 = a12036 & a11750;
assign a12040 = ~a12038 & ~a12030;
assign a12042 = ~a12040 & a11630;
assign a12044 = ~a12042 & ~a12022;
assign a12046 = ~a12044 & ~a11624;
assign a12048 = l1686 & ~l1392;
assign a12050 = a12048 & ~a11750;
assign a12052 = l1686 & ~l1390;
assign a12054 = a12052 & a11750;
assign a12056 = ~a12054 & ~a12050;
assign a12058 = ~a12056 & ~a11630;
assign a12060 = l1686 & ~l1388;
assign a12062 = a12060 & ~a11750;
assign a12064 = l1686 & ~l1386;
assign a12066 = a12064 & a11750;
assign a12068 = ~a12066 & ~a12062;
assign a12070 = ~a12068 & a11630;
assign a12072 = ~a12070 & ~a12058;
assign a12074 = ~a12072 & a11624;
assign a12076 = ~a12074 & ~a12046;
assign a12078 = ~a12076 & ~a11622;
assign a12080 = l1686 & ~l1384;
assign a12082 = a12080 & ~a11750;
assign a12084 = l1686 & ~l1382;
assign a12086 = a12084 & a11750;
assign a12088 = ~a12086 & ~a12082;
assign a12090 = ~a12088 & a11832;
assign a12092 = ~a12090 & ~a12078;
assign a12094 = ~a12092 & a11902;
assign a12096 = l1686 & ~l1380;
assign a12098 = a12096 & ~a11750;
assign a12100 = a11732 & ~a4226;
assign a12102 = ~a12100 & ~l1686;
assign a12104 = l1686 & l1378;
assign a12106 = ~a12104 & ~a12102;
assign a12108 = a12106 & a11750;
assign a12110 = ~a12108 & ~a12098;
assign a12112 = ~a12110 & ~a11630;
assign a12114 = l1686 & ~l1376;
assign a12116 = a12114 & ~a11750;
assign a12118 = l1686 & ~l1374;
assign a12120 = a12118 & a11750;
assign a12122 = ~a12120 & ~a12116;
assign a12124 = ~a12122 & a11630;
assign a12126 = ~a12124 & ~a12112;
assign a12128 = ~a12126 & ~a11624;
assign a12130 = l1686 & ~l1372;
assign a12132 = a12130 & ~a11750;
assign a12134 = l1686 & ~l1370;
assign a12136 = a12134 & a11750;
assign a12138 = ~a12136 & ~a12132;
assign a12140 = ~a12138 & ~a11630;
assign a12142 = l1686 & ~l1368;
assign a12144 = a12142 & ~a11750;
assign a12146 = l1686 & ~l1366;
assign a12148 = a12146 & a11750;
assign a12150 = ~a12148 & ~a12144;
assign a12152 = ~a12150 & a11630;
assign a12154 = ~a12152 & ~a12140;
assign a12156 = ~a12154 & a11624;
assign a12158 = ~a12156 & ~a12128;
assign a12160 = ~a12158 & ~a11622;
assign a12162 = l1686 & ~l1364;
assign a12164 = a12162 & ~a11750;
assign a12166 = l1686 & ~l1362;
assign a12168 = a12166 & a11750;
assign a12170 = ~a12168 & ~a12164;
assign a12172 = ~a12170 & a11832;
assign a12174 = ~a12172 & ~a12160;
assign a12176 = ~a12174 & ~a11902;
assign a12178 = ~a12176 & ~a12094;
assign a12180 = ~a12178 & ~a11990;
assign a12182 = ~a8822 & ~l1686;
assign a12184 = l1686 & l1360;
assign a12186 = ~a12184 & ~a12182;
assign a12188 = ~a12186 & a11990;
assign a12190 = ~a12188 & ~a12180;
assign a12192 = ~a12190 & a11600;
assign a12194 = a12190 & ~a11600;
assign a12196 = l1686 & ~l1358;
assign a12198 = a12196 & ~a11750;
assign a12200 = a8438 & ~l1686;
assign a12202 = l1686 & l1356;
assign a12204 = ~a12202 & ~a12200;
assign a12206 = a12204 & a11750;
assign a12208 = ~a12206 & ~a12198;
assign a12210 = ~a12208 & ~a11630;
assign a12212 = a8428 & ~l1686;
assign a12214 = l1686 & l1354;
assign a12216 = ~a12214 & ~a12212;
assign a12218 = a12216 & ~a11750;
assign a12220 = ~a8422 & ~l1686;
assign a12222 = l1686 & l1352;
assign a12224 = ~a12222 & ~a12220;
assign a12226 = a12224 & a11750;
assign a12228 = ~a12226 & ~a12218;
assign a12230 = ~a12228 & a11630;
assign a12232 = ~a12230 & ~a12210;
assign a12234 = ~a12232 & ~a11624;
assign a12236 = l1686 & ~l1350;
assign a12238 = a12236 & ~a11750;
assign a12240 = l1686 & ~l1348;
assign a12242 = a12240 & a11750;
assign a12244 = ~a12242 & ~a12238;
assign a12246 = ~a12244 & ~a11630;
assign a12248 = l1686 & ~l1346;
assign a12250 = a12248 & ~a11750;
assign a12252 = l1686 & ~l1344;
assign a12254 = a12252 & a11750;
assign a12256 = ~a12254 & ~a12250;
assign a12258 = ~a12256 & a11630;
assign a12260 = ~a12258 & ~a12246;
assign a12262 = ~a12260 & a11624;
assign a12264 = ~a12262 & ~a12234;
assign a12266 = ~a12264 & ~a11622;
assign a12268 = l1686 & ~l1342;
assign a12270 = a12268 & ~a11750;
assign a12272 = l1686 & ~l1340;
assign a12274 = a12272 & a11750;
assign a12276 = ~a12274 & ~a12270;
assign a12278 = ~a12276 & a11832;
assign a12280 = ~a12278 & ~a12266;
assign a12282 = ~a12280 & a11902;
assign a12284 = a8302 & ~a4156;
assign a12286 = a12284 & a8228;
assign a12288 = ~a11734 & a4160;
assign a12290 = ~a12288 & ~a12286;
assign a12292 = a12290 & ~l1686;
assign a12294 = l1686 & l1338;
assign a12296 = ~a12294 & ~a12292;
assign a12298 = a12296 & ~a11750;
assign a12300 = a12284 & ~a8228;
assign a12302 = ~a12300 & ~l1686;
assign a12304 = l1686 & l1336;
assign a12306 = ~a12304 & ~a12302;
assign a12308 = a12306 & a11750;
assign a12310 = ~a12308 & ~a12298;
assign a12312 = ~a12310 & ~a11630;
assign a12314 = l1686 & ~l1334;
assign a12316 = a12314 & ~a11750;
assign a12318 = l1686 & ~l1332;
assign a12320 = a12318 & a11750;
assign a12322 = ~a12320 & ~a12316;
assign a12324 = ~a12322 & a11630;
assign a12326 = ~a12324 & ~a12312;
assign a12328 = ~a12326 & ~a11624;
assign a12330 = l1686 & ~l1330;
assign a12332 = a12330 & ~a11750;
assign a12334 = l1686 & ~l1328;
assign a12336 = a12334 & a11750;
assign a12338 = ~a12336 & ~a12332;
assign a12340 = ~a12338 & ~a11630;
assign a12342 = l1686 & ~l1326;
assign a12344 = a12342 & ~a11750;
assign a12346 = l1686 & ~l1324;
assign a12348 = a12346 & a11750;
assign a12350 = ~a12348 & ~a12344;
assign a12352 = ~a12350 & a11630;
assign a12354 = ~a12352 & ~a12340;
assign a12356 = ~a12354 & a11624;
assign a12358 = ~a12356 & ~a12328;
assign a12360 = ~a12358 & ~a11622;
assign a12362 = l1686 & ~l1322;
assign a12364 = a12362 & ~a11750;
assign a12366 = l1686 & ~l1320;
assign a12368 = a12366 & a11750;
assign a12370 = ~a12368 & ~a12364;
assign a12372 = ~a12370 & a11832;
assign a12374 = ~a12372 & ~a12360;
assign a12376 = ~a12374 & ~a11902;
assign a12378 = ~a12376 & ~a12282;
assign a12380 = ~a12378 & ~a11990;
assign a12382 = ~a8764 & ~l1686;
assign a12384 = l1686 & l1318;
assign a12386 = ~a12384 & ~a12382;
assign a12388 = ~a12386 & a11990;
assign a12390 = ~a12388 & ~a12380;
assign a12392 = ~a12390 & a11586;
assign a12394 = a12390 & ~a11586;
assign a12396 = l1686 & ~l1316;
assign a12398 = a12396 & ~a11750;
assign a12400 = a8398 & ~l1686;
assign a12402 = l1686 & l1314;
assign a12404 = ~a12402 & ~a12400;
assign a12406 = a12404 & a11750;
assign a12408 = ~a12406 & ~a12398;
assign a12410 = ~a12408 & ~a11630;
assign a12412 = a8388 & ~l1686;
assign a12414 = l1686 & l1312;
assign a12416 = ~a12414 & ~a12412;
assign a12418 = a12416 & ~a11750;
assign a12420 = ~a8382 & ~l1686;
assign a12422 = l1686 & l1310;
assign a12424 = ~a12422 & ~a12420;
assign a12426 = a12424 & a11750;
assign a12428 = ~a12426 & ~a12418;
assign a12430 = ~a12428 & a11630;
assign a12432 = ~a12430 & ~a12410;
assign a12434 = ~a12432 & ~a11624;
assign a12436 = l1686 & ~l1308;
assign a12438 = a12436 & ~a11750;
assign a12440 = l1686 & ~l1306;
assign a12442 = a12440 & a11750;
assign a12444 = ~a12442 & ~a12438;
assign a12446 = ~a12444 & ~a11630;
assign a12448 = l1686 & ~l1304;
assign a12450 = a12448 & ~a11750;
assign a12452 = l1686 & ~l1302;
assign a12454 = a12452 & a11750;
assign a12456 = ~a12454 & ~a12450;
assign a12458 = ~a12456 & a11630;
assign a12460 = ~a12458 & ~a12446;
assign a12462 = ~a12460 & a11624;
assign a12464 = ~a12462 & ~a12434;
assign a12466 = ~a12464 & ~a11622;
assign a12468 = l1686 & ~l1300;
assign a12470 = a12468 & ~a11750;
assign a12472 = l1686 & ~l1298;
assign a12474 = a12472 & a11750;
assign a12476 = ~a12474 & ~a12470;
assign a12478 = ~a12476 & a11832;
assign a12480 = ~a12478 & ~a12466;
assign a12482 = ~a12480 & a11902;
assign a12484 = a8302 & ~a4078;
assign a12486 = a12484 & a8228;
assign a12488 = ~a11734 & a4082;
assign a12490 = ~a12488 & ~a12486;
assign a12492 = a12490 & ~l1686;
assign a12494 = l1686 & l1296;
assign a12496 = ~a12494 & ~a12492;
assign a12498 = a12496 & ~a11750;
assign a12500 = a12484 & ~a8228;
assign a12502 = ~a12500 & ~l1686;
assign a12504 = l1686 & l1294;
assign a12506 = ~a12504 & ~a12502;
assign a12508 = a12506 & a11750;
assign a12510 = ~a12508 & ~a12498;
assign a12512 = ~a12510 & ~a11630;
assign a12514 = l1686 & ~l1292;
assign a12516 = a12514 & ~a11750;
assign a12518 = l1686 & ~l1290;
assign a12520 = a12518 & a11750;
assign a12522 = ~a12520 & ~a12516;
assign a12524 = ~a12522 & a11630;
assign a12526 = ~a12524 & ~a12512;
assign a12528 = ~a12526 & ~a11624;
assign a12530 = l1686 & ~l1288;
assign a12532 = a12530 & ~a11750;
assign a12534 = l1686 & ~l1286;
assign a12536 = a12534 & a11750;
assign a12538 = ~a12536 & ~a12532;
assign a12540 = ~a12538 & ~a11630;
assign a12542 = l1686 & ~l1284;
assign a12544 = a12542 & ~a11750;
assign a12546 = l1686 & ~l1282;
assign a12548 = a12546 & a11750;
assign a12550 = ~a12548 & ~a12544;
assign a12552 = ~a12550 & a11630;
assign a12554 = ~a12552 & ~a12540;
assign a12556 = ~a12554 & a11624;
assign a12558 = ~a12556 & ~a12528;
assign a12560 = ~a12558 & ~a11622;
assign a12562 = l1686 & ~l1280;
assign a12564 = a12562 & ~a11750;
assign a12566 = l1686 & ~l1278;
assign a12568 = a12566 & a11750;
assign a12570 = ~a12568 & ~a12564;
assign a12572 = ~a12570 & a11832;
assign a12574 = ~a12572 & ~a12560;
assign a12576 = ~a12574 & ~a11902;
assign a12578 = ~a12576 & ~a12482;
assign a12580 = ~a12578 & ~a11990;
assign a12582 = ~a8706 & ~l1686;
assign a12584 = l1686 & l1276;
assign a12586 = ~a12584 & ~a12582;
assign a12588 = ~a12586 & a11990;
assign a12590 = ~a12588 & ~a12580;
assign a12592 = ~a12590 & a11572;
assign a12594 = a12590 & ~a11572;
assign a12596 = l1686 & ~l1274;
assign a12598 = a12596 & ~a11750;
assign a12600 = a8358 & ~l1686;
assign a12602 = l1686 & l1272;
assign a12604 = ~a12602 & ~a12600;
assign a12606 = a12604 & a11750;
assign a12608 = ~a12606 & ~a12598;
assign a12610 = ~a12608 & ~a11630;
assign a12612 = a8348 & ~l1686;
assign a12614 = l1686 & l1270;
assign a12616 = ~a12614 & ~a12612;
assign a12618 = a12616 & ~a11750;
assign a12620 = ~a8342 & ~l1686;
assign a12622 = l1686 & l1268;
assign a12624 = ~a12622 & ~a12620;
assign a12626 = a12624 & a11750;
assign a12628 = ~a12626 & ~a12618;
assign a12630 = ~a12628 & a11630;
assign a12632 = ~a12630 & ~a12610;
assign a12634 = ~a12632 & ~a11624;
assign a12636 = l1686 & ~l1266;
assign a12638 = a12636 & ~a11750;
assign a12640 = l1686 & ~l1264;
assign a12642 = a12640 & a11750;
assign a12644 = ~a12642 & ~a12638;
assign a12646 = ~a12644 & ~a11630;
assign a12648 = l1686 & ~l1262;
assign a12650 = a12648 & ~a11750;
assign a12652 = l1686 & ~l1260;
assign a12654 = a12652 & a11750;
assign a12656 = ~a12654 & ~a12650;
assign a12658 = ~a12656 & a11630;
assign a12660 = ~a12658 & ~a12646;
assign a12662 = ~a12660 & a11624;
assign a12664 = ~a12662 & ~a12634;
assign a12666 = ~a12664 & ~a11622;
assign a12668 = l1686 & ~l1258;
assign a12670 = a12668 & ~a11750;
assign a12672 = l1686 & ~l1256;
assign a12674 = a12672 & a11750;
assign a12676 = ~a12674 & ~a12670;
assign a12678 = ~a12676 & a11832;
assign a12680 = ~a12678 & ~a12666;
assign a12682 = ~a12680 & a11902;
assign a12684 = a8302 & ~a4000;
assign a12686 = a12684 & a8228;
assign a12688 = ~a11734 & a4004;
assign a12690 = ~a12688 & ~a12686;
assign a12692 = a12690 & ~l1686;
assign a12694 = l1686 & l1254;
assign a12696 = ~a12694 & ~a12692;
assign a12698 = a12696 & ~a11750;
assign a12700 = a12684 & ~a8228;
assign a12702 = ~a12700 & ~l1686;
assign a12704 = l1686 & l1252;
assign a12706 = ~a12704 & ~a12702;
assign a12708 = a12706 & a11750;
assign a12710 = ~a12708 & ~a12698;
assign a12712 = ~a12710 & ~a11630;
assign a12714 = l1686 & ~l1250;
assign a12716 = a12714 & ~a11750;
assign a12718 = l1686 & ~l1248;
assign a12720 = a12718 & a11750;
assign a12722 = ~a12720 & ~a12716;
assign a12724 = ~a12722 & a11630;
assign a12726 = ~a12724 & ~a12712;
assign a12728 = ~a12726 & ~a11624;
assign a12730 = l1686 & ~l1246;
assign a12732 = a12730 & ~a11750;
assign a12734 = l1686 & ~l1244;
assign a12736 = a12734 & a11750;
assign a12738 = ~a12736 & ~a12732;
assign a12740 = ~a12738 & ~a11630;
assign a12742 = l1686 & ~l1242;
assign a12744 = a12742 & ~a11750;
assign a12746 = l1686 & ~l1240;
assign a12748 = a12746 & a11750;
assign a12750 = ~a12748 & ~a12744;
assign a12752 = ~a12750 & a11630;
assign a12754 = ~a12752 & ~a12740;
assign a12756 = ~a12754 & a11624;
assign a12758 = ~a12756 & ~a12728;
assign a12760 = ~a12758 & ~a11622;
assign a12762 = l1686 & ~l1238;
assign a12764 = a12762 & ~a11750;
assign a12766 = l1686 & ~l1236;
assign a12768 = a12766 & a11750;
assign a12770 = ~a12768 & ~a12764;
assign a12772 = ~a12770 & a11832;
assign a12774 = ~a12772 & ~a12760;
assign a12776 = ~a12774 & ~a11902;
assign a12778 = ~a12776 & ~a12682;
assign a12780 = ~a12778 & ~a11990;
assign a12782 = ~a8648 & ~l1686;
assign a12784 = l1686 & l1234;
assign a12786 = ~a12784 & ~a12782;
assign a12788 = ~a12786 & a11990;
assign a12790 = ~a12788 & ~a12780;
assign a12792 = ~a12790 & a11558;
assign a12794 = a12790 & ~a11558;
assign a12796 = l1686 & ~l1232;
assign a12798 = a12796 & ~a11750;
assign a12800 = a8324 & ~l1686;
assign a12802 = l1686 & l1230;
assign a12804 = ~a12802 & ~a12800;
assign a12806 = a12804 & a11750;
assign a12808 = ~a12806 & ~a12798;
assign a12810 = ~a12808 & ~a11630;
assign a12812 = a8314 & ~l1686;
assign a12814 = l1686 & l1228;
assign a12816 = ~a12814 & ~a12812;
assign a12818 = a12816 & ~a11750;
assign a12820 = ~a8308 & ~l1686;
assign a12822 = l1686 & l1226;
assign a12824 = ~a12822 & ~a12820;
assign a12826 = a12824 & a11750;
assign a12828 = ~a12826 & ~a12818;
assign a12830 = ~a12828 & a11630;
assign a12832 = ~a12830 & ~a12810;
assign a12834 = ~a12832 & ~a11624;
assign a12836 = l1686 & ~l1224;
assign a12838 = a12836 & ~a11750;
assign a12840 = l1686 & ~l1222;
assign a12842 = a12840 & a11750;
assign a12844 = ~a12842 & ~a12838;
assign a12846 = ~a12844 & ~a11630;
assign a12848 = l1686 & ~l1220;
assign a12850 = a12848 & ~a11750;
assign a12852 = l1686 & ~l1218;
assign a12854 = a12852 & a11750;
assign a12856 = ~a12854 & ~a12850;
assign a12858 = ~a12856 & a11630;
assign a12860 = ~a12858 & ~a12846;
assign a12862 = ~a12860 & a11624;
assign a12864 = ~a12862 & ~a12834;
assign a12866 = ~a12864 & ~a11622;
assign a12868 = l1686 & ~l1216;
assign a12870 = a12868 & ~a11750;
assign a12872 = l1686 & ~l1214;
assign a12874 = a12872 & a11750;
assign a12876 = ~a12874 & ~a12870;
assign a12878 = ~a12876 & a11832;
assign a12880 = ~a12878 & ~a12866;
assign a12882 = ~a12880 & a11902;
assign a12884 = a8302 & ~a3922;
assign a12886 = a12884 & a8228;
assign a12888 = ~a11734 & a3926;
assign a12890 = ~a12888 & ~a12886;
assign a12892 = a12890 & ~l1686;
assign a12894 = l1686 & l1212;
assign a12896 = ~a12894 & ~a12892;
assign a12898 = a12896 & ~a11750;
assign a12900 = a12884 & ~a8228;
assign a12902 = ~a12900 & ~l1686;
assign a12904 = l1686 & l1210;
assign a12906 = ~a12904 & ~a12902;
assign a12908 = a12906 & a11750;
assign a12910 = ~a12908 & ~a12898;
assign a12912 = ~a12910 & ~a11630;
assign a12914 = l1686 & ~l1208;
assign a12916 = a12914 & ~a11750;
assign a12918 = l1686 & ~l1206;
assign a12920 = a12918 & a11750;
assign a12922 = ~a12920 & ~a12916;
assign a12924 = ~a12922 & a11630;
assign a12926 = ~a12924 & ~a12912;
assign a12928 = ~a12926 & ~a11624;
assign a12930 = l1686 & ~l1204;
assign a12932 = a12930 & ~a11750;
assign a12934 = l1686 & ~l1202;
assign a12936 = a12934 & a11750;
assign a12938 = ~a12936 & ~a12932;
assign a12940 = ~a12938 & ~a11630;
assign a12942 = l1686 & ~l1200;
assign a12944 = a12942 & ~a11750;
assign a12946 = l1686 & ~l1198;
assign a12948 = a12946 & a11750;
assign a12950 = ~a12948 & ~a12944;
assign a12952 = ~a12950 & a11630;
assign a12954 = ~a12952 & ~a12940;
assign a12956 = ~a12954 & a11624;
assign a12958 = ~a12956 & ~a12928;
assign a12960 = ~a12958 & ~a11622;
assign a12962 = l1686 & ~l1196;
assign a12964 = a12962 & ~a11750;
assign a12966 = l1686 & ~l1194;
assign a12968 = a12966 & a11750;
assign a12970 = ~a12968 & ~a12964;
assign a12972 = ~a12970 & a11832;
assign a12974 = ~a12972 & ~a12960;
assign a12976 = ~a12974 & ~a11902;
assign a12978 = ~a12976 & ~a12882;
assign a12980 = ~a12978 & ~a11990;
assign a12982 = ~a8594 & ~l1686;
assign a12984 = l1686 & l1192;
assign a12986 = ~a12984 & ~a12982;
assign a12988 = ~a12986 & a11990;
assign a12990 = ~a12988 & ~a12980;
assign a12992 = ~a12990 & a11538;
assign a12994 = a12990 & ~a11538;
assign a12996 = ~a11750 & a11304;
assign a12998 = a11750 & a11316;
assign a13000 = ~a12998 & ~a12996;
assign a13002 = ~a13000 & ~a11630;
assign a13004 = ~a11750 & a11328;
assign a13006 = a11750 & a11336;
assign a13008 = ~a13006 & ~a13004;
assign a13010 = ~a13008 & a11630;
assign a13012 = ~a13010 & ~a13002;
assign a13014 = ~a13012 & ~a11624;
assign a13016 = ~a11750 & a11348;
assign a13018 = a11750 & a11352;
assign a13020 = ~a13018 & ~a13016;
assign a13022 = ~a13020 & ~a11630;
assign a13024 = ~a11750 & a11360;
assign a13026 = a11750 & a11364;
assign a13028 = ~a13026 & ~a13024;
assign a13030 = ~a13028 & a11630;
assign a13032 = ~a13030 & ~a13022;
assign a13034 = ~a13032 & a11624;
assign a13036 = ~a13034 & ~a13014;
assign a13038 = ~a13036 & ~a11622;
assign a13040 = ~a11750 & a11292;
assign a13042 = a11750 & a11296;
assign a13044 = ~a13042 & ~a13040;
assign a13046 = ~a13044 & a11832;
assign a13048 = ~a13046 & ~a13038;
assign a13050 = ~a13048 & a11902;
assign a13052 = a8302 & a3852;
assign a13054 = ~a8302 & i300;
assign a13056 = ~a13054 & ~a13052;
assign a13058 = a13056 & a11734;
assign a13060 = ~a11734 & a3860;
assign a13062 = ~a13060 & ~a13058;
assign a13064 = a13062 & ~l1686;
assign a13066 = l1686 & l1170;
assign a13068 = ~a13066 & ~a13064;
assign a13070 = a13068 & ~a11750;
assign a13072 = a13056 & a11732;
assign a13074 = ~a13072 & ~l1686;
assign a13076 = l1686 & l1168;
assign a13078 = ~a13076 & ~a13074;
assign a13080 = a13078 & a11750;
assign a13082 = ~a13080 & ~a13070;
assign a13084 = ~a13082 & ~a11630;
assign a13086 = l1686 & ~l1166;
assign a13088 = a13086 & ~a11750;
assign a13090 = l1686 & ~l1164;
assign a13092 = a13090 & a11750;
assign a13094 = ~a13092 & ~a13088;
assign a13096 = ~a13094 & a11630;
assign a13098 = ~a13096 & ~a13084;
assign a13100 = ~a13098 & ~a11624;
assign a13102 = l1686 & ~l1162;
assign a13104 = a13102 & ~a11750;
assign a13106 = l1686 & ~l1160;
assign a13108 = a13106 & a11750;
assign a13110 = ~a13108 & ~a13104;
assign a13112 = ~a13110 & ~a11630;
assign a13114 = l1686 & ~l1158;
assign a13116 = a13114 & ~a11750;
assign a13118 = l1686 & ~l1156;
assign a13120 = a13118 & a11750;
assign a13122 = ~a13120 & ~a13116;
assign a13124 = ~a13122 & a11630;
assign a13126 = ~a13124 & ~a13112;
assign a13128 = ~a13126 & a11624;
assign a13130 = ~a13128 & ~a13100;
assign a13132 = ~a13130 & ~a11622;
assign a13134 = l1686 & ~l1154;
assign a13136 = a13134 & ~a11750;
assign a13138 = l1686 & ~l1152;
assign a13140 = a13138 & a11750;
assign a13142 = ~a13140 & ~a13136;
assign a13144 = ~a13142 & a11832;
assign a13146 = ~a13144 & ~a13132;
assign a13148 = ~a13146 & ~a11902;
assign a13150 = ~a13148 & ~a13050;
assign a13152 = ~a13150 & ~a11990;
assign a13154 = ~a8544 & ~l1686;
assign a13156 = l1686 & l1150;
assign a13158 = ~a13156 & ~a13154;
assign a13160 = ~a13158 & a11990;
assign a13162 = ~a13160 & ~a13152;
assign a13164 = a13162 & ~a11544;
assign a13166 = ~a13164 & ~a12994;
assign a13168 = ~a13166 & ~a12992;
assign a13170 = ~a13168 & ~a12794;
assign a13172 = ~a13170 & ~a12792;
assign a13174 = ~a13172 & ~a12594;
assign a13176 = ~a13174 & ~a12592;
assign a13178 = ~a13176 & ~a12394;
assign a13180 = ~a13178 & ~a12392;
assign a13182 = ~a13180 & ~a12194;
assign a13184 = ~a13182 & ~a12192;
assign a13186 = ~a13184 & ~a12006;
assign a13188 = ~a13186 & ~a12004;
assign a13190 = ~a11194 & ~a8062;
assign a13192 = a8870 & a8062;
assign a13194 = ~a13192 & ~a13190;
assign a13196 = ~a11750 & a11214;
assign a13198 = a11750 & a11222;
assign a13200 = ~a13198 & ~a13196;
assign a13202 = ~a13200 & ~a11630;
assign a13204 = ~a11750 & a11230;
assign a13206 = a11750 & a11234;
assign a13208 = ~a13206 & ~a13204;
assign a13210 = ~a13208 & a11630;
assign a13212 = ~a13210 & ~a13202;
assign a13214 = ~a13212 & ~a11624;
assign a13216 = ~a11750 & a11246;
assign a13218 = a11750 & a11250;
assign a13220 = ~a13218 & ~a13216;
assign a13222 = ~a13220 & ~a11630;
assign a13224 = ~a11750 & a11258;
assign a13226 = a11750 & a11262;
assign a13228 = ~a13226 & ~a13224;
assign a13230 = ~a13228 & a11630;
assign a13232 = ~a13230 & ~a13222;
assign a13234 = ~a13232 & a11624;
assign a13236 = ~a13234 & ~a13214;
assign a13238 = ~a13236 & ~a11622;
assign a13240 = ~a11750 & a11202;
assign a13242 = a11750 & a11206;
assign a13244 = ~a13242 & ~a13240;
assign a13246 = ~a13244 & a11832;
assign a13248 = ~a13246 & ~a13238;
assign a13250 = ~a13248 & a11902;
assign a13252 = l1686 & ~l1128;
assign a13254 = a13252 & ~a11750;
assign a13256 = l1686 & ~l1126;
assign a13258 = a13256 & a11750;
assign a13260 = ~a13258 & ~a13254;
assign a13262 = ~a13260 & ~a11630;
assign a13264 = l1686 & ~l1124;
assign a13266 = a13264 & ~a11750;
assign a13268 = l1686 & ~l1122;
assign a13270 = a13268 & a11750;
assign a13272 = ~a13270 & ~a13266;
assign a13274 = ~a13272 & a11630;
assign a13276 = ~a13274 & ~a13262;
assign a13278 = ~a13276 & ~a11624;
assign a13280 = l1686 & ~l1120;
assign a13282 = a13280 & ~a11750;
assign a13284 = l1686 & ~l1118;
assign a13286 = a13284 & a11750;
assign a13288 = ~a13286 & ~a13282;
assign a13290 = ~a13288 & ~a11630;
assign a13292 = l1686 & ~l1116;
assign a13294 = a13292 & ~a11750;
assign a13296 = l1686 & ~l1114;
assign a13298 = a13296 & a11750;
assign a13300 = ~a13298 & ~a13294;
assign a13302 = ~a13300 & a11630;
assign a13304 = ~a13302 & ~a13290;
assign a13306 = ~a13304 & a11624;
assign a13308 = ~a13306 & ~a13278;
assign a13310 = ~a13308 & ~a11622;
assign a13312 = l1686 & ~l1112;
assign a13314 = a13312 & ~a11750;
assign a13316 = l1686 & ~l1110;
assign a13318 = a13316 & a11750;
assign a13320 = ~a13318 & ~a13314;
assign a13322 = ~a13320 & a11832;
assign a13324 = ~a13322 & ~a13310;
assign a13326 = ~a13324 & ~a11902;
assign a13328 = ~a13326 & ~a13250;
assign a13330 = ~a13328 & ~a11990;
assign a13332 = l1686 & ~l994;
assign a13334 = a13332 & a11990;
assign a13336 = ~a13334 & ~a13330;
assign a13338 = a13336 & ~a13194;
assign a13340 = ~a13336 & a13194;
assign a13342 = ~a13340 & ~a13338;
assign a13344 = ~a13342 & ~a13188;
assign a13346 = a13342 & a13188;
assign a13348 = ~a13346 & ~a13344;
assign a13350 = a13348 & ~a11620;
assign a13352 = ~a13348 & ~a12002;
assign a13354 = ~a13352 & ~a13350;
assign a13356 = ~a13354 & ~a8874;
assign a13358 = a13354 & a8874;
assign a13360 = ~a11600 & ~a11588;
assign a13362 = ~a13360 & ~a11602;
assign a13364 = ~a13362 & a13348;
assign a13366 = ~a13348 & ~a12190;
assign a13368 = ~a13366 & ~a13364;
assign a13370 = ~a13368 & ~a10044;
assign a13372 = a13368 & a10044;
assign a13374 = ~a11586 & ~a11574;
assign a13376 = ~a13374 & ~a11588;
assign a13378 = ~a13376 & a13348;
assign a13380 = ~a13348 & ~a12390;
assign a13382 = ~a13380 & ~a13378;
assign a13384 = ~a13382 & ~a10074;
assign a13386 = a13382 & a10074;
assign a13388 = ~a11572 & ~a11560;
assign a13390 = ~a13388 & ~a11574;
assign a13392 = ~a13390 & a13348;
assign a13394 = ~a13348 & ~a12590;
assign a13396 = ~a13394 & ~a13392;
assign a13398 = ~a13396 & ~a10100;
assign a13400 = a13396 & a10100;
assign a13402 = ~a11558 & ~a11546;
assign a13404 = ~a13402 & ~a11560;
assign a13406 = ~a13404 & a13348;
assign a13408 = ~a13348 & ~a12790;
assign a13410 = ~a13408 & ~a13406;
assign a13412 = ~a13410 & ~a10126;
assign a13414 = a13410 & a10126;
assign a13416 = ~a11544 & ~a11538;
assign a13418 = ~a13416 & ~a11546;
assign a13420 = ~a13418 & a13348;
assign a13422 = ~a13348 & ~a12990;
assign a13424 = ~a13422 & ~a13420;
assign a13426 = ~a13424 & ~a10152;
assign a13428 = a13424 & a10152;
assign a13430 = ~a13348 & ~a13162;
assign a13432 = a13348 & a11544;
assign a13434 = ~a13432 & a10178;
assign a13436 = a13434 & ~a13430;
assign a13438 = ~a13436 & ~a13428;
assign a13440 = ~a13438 & ~a13426;
assign a13442 = ~a13440 & ~a13414;
assign a13444 = ~a13442 & ~a13412;
assign a13446 = ~a13444 & ~a13400;
assign a13448 = ~a13446 & ~a13398;
assign a13450 = ~a13448 & ~a13386;
assign a13452 = ~a13450 & ~a13384;
assign a13454 = ~a13452 & ~a13372;
assign a13456 = ~a13454 & ~a13370;
assign a13458 = ~a13456 & ~a13358;
assign a13460 = ~a13458 & ~a13356;
assign a13462 = a13194 & a11618;
assign a13464 = ~a13194 & ~a11618;
assign a13466 = ~a13464 & ~a13462;
assign a13468 = ~a13466 & a13348;
assign a13470 = ~a13348 & ~a13336;
assign a13472 = ~a13470 & ~a13468;
assign a13474 = ~a13472 & ~a8868;
assign a13476 = a13472 & a8868;
assign a13478 = ~a13476 & ~a13474;
assign a13480 = ~a13478 & a13460;
assign a13482 = a13478 & ~a13460;
assign a13484 = ~a13482 & ~a13480;
assign a13486 = ~a13484 & ~l988;
assign a13488 = a13486 & ~a11526;
assign a13490 = a13488 & ~a8032;
assign a13492 = ~a6682 & ~l494;
assign a13494 = a13492 & ~l664;
assign a13496 = a13494 & a13490;
assign a13498 = ~l1686 & i214;
assign a13500 = l1686 & l990;
assign a13502 = ~a13500 & ~a13498;
assign a13504 = ~a13502 & ~l988;
assign a13506 = a13504 & ~i216;
assign a13508 = a13506 & a13496;
assign a13510 = a13508 & l582;
assign a13512 = i312 & i216;
assign a13514 = ~a13508 & i310;
assign a13516 = a13508 & a10178;
assign a13518 = ~a13516 & ~a13514;
assign a13520 = ~a13518 & ~i216;
assign a13522 = ~a13520 & ~a13512;
assign a13524 = ~a13522 & ~a11364;
assign a13526 = i316 & i216;
assign a13528 = ~a13508 & i314;
assign a13530 = a13508 & a10152;
assign a13532 = ~a13530 & ~a13528;
assign a13534 = ~a13532 & ~i216;
assign a13536 = ~a13534 & ~a13526;
assign a13538 = ~a13536 & ~a12852;
assign a13540 = ~a13538 & ~a13524;
assign a13542 = a13536 & a12852;
assign a13544 = ~a13542 & ~a13540;
assign a13546 = i320 & i216;
assign a13548 = ~a13508 & i318;
assign a13550 = a13508 & a10126;
assign a13552 = ~a13550 & ~a13548;
assign a13554 = ~a13552 & ~i216;
assign a13556 = ~a13554 & ~a13546;
assign a13558 = ~a13556 & ~a12652;
assign a13560 = ~a13558 & ~a13544;
assign a13562 = a13556 & a12652;
assign a13564 = ~a13562 & ~a13560;
assign a13566 = i324 & i216;
assign a13568 = ~a13508 & i322;
assign a13570 = a13508 & a10100;
assign a13572 = ~a13570 & ~a13568;
assign a13574 = ~a13572 & ~i216;
assign a13576 = ~a13574 & ~a13566;
assign a13578 = ~a13576 & ~a12452;
assign a13580 = ~a13578 & ~a13564;
assign a13582 = a13576 & a12452;
assign a13584 = ~a13582 & ~a13580;
assign a13586 = i328 & i216;
assign a13588 = ~a13508 & i326;
assign a13590 = a13508 & a10074;
assign a13592 = ~a13590 & ~a13588;
assign a13594 = ~a13592 & ~i216;
assign a13596 = ~a13594 & ~a13586;
assign a13598 = ~a13596 & ~a12252;
assign a13600 = ~a13598 & ~a13584;
assign a13602 = a13596 & a12252;
assign a13604 = ~a13602 & ~a13600;
assign a13606 = i332 & i216;
assign a13608 = ~a13508 & i330;
assign a13610 = a13508 & a10044;
assign a13612 = ~a13610 & ~a13608;
assign a13614 = ~a13612 & ~i216;
assign a13616 = ~a13614 & ~a13606;
assign a13618 = ~a13616 & ~a12064;
assign a13620 = ~a13618 & ~a13604;
assign a13622 = a13616 & a12064;
assign a13624 = ~a13622 & ~a13620;
assign a13626 = i308 & i216;
assign a13628 = ~a13508 & i306;
assign a13630 = a13508 & a8874;
assign a13632 = ~a13630 & ~a13628;
assign a13634 = ~a13632 & ~i216;
assign a13636 = ~a13634 & ~a13626;
assign a13638 = ~a13636 & ~a11804;
assign a13640 = ~a13638 & ~a13624;
assign a13642 = a13636 & a11804;
assign a13644 = ~a13642 & ~a13640;
assign a13646 = i304 & i216;
assign a13648 = ~a13508 & i302;
assign a13650 = a13508 & a8868;
assign a13652 = ~a13650 & ~a13648;
assign a13654 = ~a13652 & ~i216;
assign a13656 = ~a13654 & ~a13646;
assign a13658 = a13656 & a11262;
assign a13660 = ~a13656 & ~a11262;
assign a13662 = ~a13660 & ~a13658;
assign a13664 = ~a13662 & ~a13644;
assign a13666 = a13522 & a11364;
assign a13668 = ~a13666 & ~a13542;
assign a13670 = ~a13668 & ~a13538;
assign a13672 = ~a13670 & ~a13562;
assign a13674 = ~a13672 & ~a13558;
assign a13676 = ~a13674 & ~a13582;
assign a13678 = ~a13676 & ~a13578;
assign a13680 = ~a13678 & ~a13602;
assign a13682 = ~a13680 & ~a13598;
assign a13684 = ~a13682 & ~a13622;
assign a13686 = ~a13684 & ~a13618;
assign a13688 = ~a13686 & ~a13642;
assign a13690 = ~a13688 & ~a13638;
assign a13692 = ~a13690 & a13662;
assign a13694 = ~a13692 & ~a13664;
assign a13696 = l1686 & ~l1466;
assign a13698 = ~a5550 & ~l1686;
assign a13700 = l1686 & l1468;
assign a13702 = ~a13700 & ~a13698;
assign a13704 = ~a8230 & ~l1686;
assign a13706 = l1686 & l1462;
assign a13708 = ~a13706 & ~a13704;
assign a13710 = l1686 & ~l1464;
assign a13712 = ~a13710 & a13708;
assign a13714 = a13712 & a13702;
assign a13716 = a13714 & a13696;
assign a13718 = a13636 & a11950;
assign a13720 = a13616 & a12146;
assign a13722 = ~a13720 & ~a13718;
assign a13724 = ~a13616 & ~a12146;
assign a13726 = ~a13596 & ~a12346;
assign a13728 = ~a13726 & ~a13724;
assign a13730 = a13596 & a12346;
assign a13732 = a13576 & a12546;
assign a13734 = ~a13732 & ~a13730;
assign a13736 = ~a13576 & ~a12546;
assign a13738 = a13556 & a12746;
assign a13740 = ~a13556 & ~a12746;
assign a13742 = a13536 & a12946;
assign a13744 = ~a13536 & ~a12946;
assign a13746 = ~a13522 & ~a13118;
assign a13748 = ~a13746 & ~a13744;
assign a13750 = ~a13748 & ~a13742;
assign a13752 = ~a13750 & ~a13740;
assign a13754 = ~a13752 & ~a13738;
assign a13756 = ~a13754 & ~a13736;
assign a13758 = ~a13756 & a13734;
assign a13760 = ~a13758 & a13728;
assign a13762 = ~a13760 & a13722;
assign a13764 = ~a13636 & ~a11950;
assign a13766 = ~a13764 & ~a13762;
assign a13768 = a13656 & a13296;
assign a13770 = ~a13656 & ~a13296;
assign a13772 = ~a13770 & ~a13768;
assign a13774 = ~a13772 & ~a13766;
assign a13776 = a13772 & a13766;
assign a13778 = ~a13776 & ~a13774;
assign a13780 = ~a13778 & a13510;
assign a13782 = ~a13780 & ~a13716;
assign a13784 = ~a13782 & ~a13694;
assign a13786 = a13784 & l1094;
assign a13788 = a13786 & a13510;
assign a13790 = a13508 & l578;
assign a13792 = ~a13522 & ~a11352;
assign a13794 = ~a13536 & ~a12840;
assign a13796 = ~a13794 & ~a13792;
assign a13798 = a13536 & a12840;
assign a13800 = ~a13798 & ~a13796;
assign a13802 = ~a13556 & ~a12640;
assign a13804 = ~a13802 & ~a13800;
assign a13806 = a13556 & a12640;
assign a13808 = ~a13806 & ~a13804;
assign a13810 = ~a13576 & ~a12440;
assign a13812 = ~a13810 & ~a13808;
assign a13814 = a13576 & a12440;
assign a13816 = ~a13814 & ~a13812;
assign a13818 = ~a13596 & ~a12240;
assign a13820 = ~a13818 & ~a13816;
assign a13822 = a13596 & a12240;
assign a13824 = ~a13822 & ~a13820;
assign a13826 = ~a13616 & ~a12052;
assign a13828 = ~a13826 & ~a13824;
assign a13830 = a13616 & a12052;
assign a13832 = ~a13830 & ~a13828;
assign a13834 = ~a13636 & ~a11792;
assign a13836 = ~a13834 & ~a13832;
assign a13838 = a13636 & a11792;
assign a13840 = ~a13838 & ~a13836;
assign a13842 = a13656 & a11250;
assign a13844 = ~a13656 & ~a11250;
assign a13846 = ~a13844 & ~a13842;
assign a13848 = ~a13846 & ~a13840;
assign a13850 = a13522 & a11352;
assign a13852 = ~a13850 & ~a13798;
assign a13854 = ~a13852 & ~a13794;
assign a13856 = ~a13854 & ~a13806;
assign a13858 = ~a13856 & ~a13802;
assign a13860 = ~a13858 & ~a13814;
assign a13862 = ~a13860 & ~a13810;
assign a13864 = ~a13862 & ~a13822;
assign a13866 = ~a13864 & ~a13818;
assign a13868 = ~a13866 & ~a13830;
assign a13870 = ~a13868 & ~a13826;
assign a13872 = ~a13870 & ~a13838;
assign a13874 = ~a13872 & ~a13834;
assign a13876 = ~a13874 & a13846;
assign a13878 = ~a13876 & ~a13848;
assign a13880 = ~a13702 & a13696;
assign a13882 = a13880 & a13712;
assign a13884 = a13636 & a11938;
assign a13886 = a13616 & a12134;
assign a13888 = ~a13886 & ~a13884;
assign a13890 = ~a13616 & ~a12134;
assign a13892 = ~a13596 & ~a12334;
assign a13894 = ~a13892 & ~a13890;
assign a13896 = a13596 & a12334;
assign a13898 = a13576 & a12534;
assign a13900 = ~a13898 & ~a13896;
assign a13902 = ~a13576 & ~a12534;
assign a13904 = a13556 & a12734;
assign a13906 = ~a13556 & ~a12734;
assign a13908 = a13536 & a12934;
assign a13910 = ~a13536 & ~a12934;
assign a13912 = ~a13522 & ~a13106;
assign a13914 = ~a13912 & ~a13910;
assign a13916 = ~a13914 & ~a13908;
assign a13918 = ~a13916 & ~a13906;
assign a13920 = ~a13918 & ~a13904;
assign a13922 = ~a13920 & ~a13902;
assign a13924 = ~a13922 & a13900;
assign a13926 = ~a13924 & a13894;
assign a13928 = ~a13926 & a13888;
assign a13930 = ~a13636 & ~a11938;
assign a13932 = ~a13930 & ~a13928;
assign a13934 = a13656 & a13284;
assign a13936 = ~a13656 & ~a13284;
assign a13938 = ~a13936 & ~a13934;
assign a13940 = ~a13938 & ~a13932;
assign a13942 = a13938 & a13932;
assign a13944 = ~a13942 & ~a13940;
assign a13946 = ~a13944 & a13790;
assign a13948 = ~a13946 & ~a13882;
assign a13950 = ~a13948 & ~a13878;
assign a13952 = a13950 & l1098;
assign a13954 = a13952 & a13790;
assign a13956 = ~a13954 & ~a13788;
assign a13958 = a13508 & ~a5542;
assign a13960 = ~a13522 & ~a11304;
assign a13962 = ~a13536 & ~a12796;
assign a13964 = ~a13962 & ~a13960;
assign a13966 = a13536 & a12796;
assign a13968 = ~a13966 & ~a13964;
assign a13970 = ~a13556 & ~a12596;
assign a13972 = ~a13970 & ~a13968;
assign a13974 = a13556 & a12596;
assign a13976 = ~a13974 & ~a13972;
assign a13978 = ~a13576 & ~a12396;
assign a13980 = ~a13978 & ~a13976;
assign a13982 = a13576 & a12396;
assign a13984 = ~a13982 & ~a13980;
assign a13986 = ~a13596 & ~a12196;
assign a13988 = ~a13986 & ~a13984;
assign a13990 = a13596 & a12196;
assign a13992 = ~a13990 & ~a13988;
assign a13994 = ~a13616 & ~a12008;
assign a13996 = ~a13994 & ~a13992;
assign a13998 = a13616 & a12008;
assign a14000 = ~a13998 & ~a13996;
assign a14002 = ~a13636 & ~a11752;
assign a14004 = ~a14002 & ~a14000;
assign a14006 = a13636 & a11752;
assign a14008 = ~a14006 & ~a14004;
assign a14010 = a13656 & a11214;
assign a14012 = ~a13656 & ~a11214;
assign a14014 = ~a14012 & ~a14010;
assign a14016 = ~a14014 & ~a14008;
assign a14018 = a13522 & a11304;
assign a14020 = ~a14018 & ~a13966;
assign a14022 = ~a14020 & ~a13962;
assign a14024 = ~a14022 & ~a13974;
assign a14026 = ~a14024 & ~a13970;
assign a14028 = ~a14026 & ~a13982;
assign a14030 = ~a14028 & ~a13978;
assign a14032 = ~a14030 & ~a13990;
assign a14034 = ~a14032 & ~a13986;
assign a14036 = ~a14034 & ~a13998;
assign a14038 = ~a14036 & ~a13994;
assign a14040 = ~a14038 & ~a14006;
assign a14042 = ~a14040 & ~a14002;
assign a14044 = ~a14042 & a14014;
assign a14046 = ~a14044 & ~a14016;
assign a14048 = ~a13702 & ~a13696;
assign a14050 = ~a13710 & ~a13708;
assign a14052 = a14050 & a14048;
assign a14054 = a13636 & a11906;
assign a14056 = a13616 & a12096;
assign a14058 = ~a14056 & ~a14054;
assign a14060 = ~a13616 & ~a12096;
assign a14062 = ~a13596 & ~a12296;
assign a14064 = ~a14062 & ~a14060;
assign a14066 = a13596 & a12296;
assign a14068 = a13576 & a12496;
assign a14070 = ~a14068 & ~a14066;
assign a14072 = ~a13576 & ~a12496;
assign a14074 = a13556 & a12696;
assign a14076 = ~a13556 & ~a12696;
assign a14078 = a13536 & a12896;
assign a14080 = ~a13536 & ~a12896;
assign a14082 = ~a13522 & ~a13068;
assign a14084 = ~a14082 & ~a14080;
assign a14086 = ~a14084 & ~a14078;
assign a14088 = ~a14086 & ~a14076;
assign a14090 = ~a14088 & ~a14074;
assign a14092 = ~a14090 & ~a14072;
assign a14094 = ~a14092 & a14070;
assign a14096 = ~a14094 & a14064;
assign a14098 = ~a14096 & a14058;
assign a14100 = ~a13636 & ~a11906;
assign a14102 = ~a14100 & ~a14098;
assign a14104 = a13656 & a13252;
assign a14106 = ~a13656 & ~a13252;
assign a14108 = ~a14106 & ~a14104;
assign a14110 = ~a14108 & ~a14102;
assign a14112 = a14108 & a14102;
assign a14114 = ~a14112 & ~a14110;
assign a14116 = ~a14114 & a13958;
assign a14118 = ~a14116 & ~a14052;
assign a14120 = ~a14118 & ~a14046;
assign a14122 = a14120 & ~a11842;
assign a14124 = a14122 & a13958;
assign a14126 = a13508 & l586;
assign a14128 = ~a13522 & ~a11292;
assign a14130 = ~a13536 & ~a12868;
assign a14132 = ~a14130 & ~a14128;
assign a14134 = a13536 & a12868;
assign a14136 = ~a14134 & ~a14132;
assign a14138 = ~a13556 & ~a12668;
assign a14140 = ~a14138 & ~a14136;
assign a14142 = a13556 & a12668;
assign a14144 = ~a14142 & ~a14140;
assign a14146 = ~a13576 & ~a12468;
assign a14148 = ~a14146 & ~a14144;
assign a14150 = a13576 & a12468;
assign a14152 = ~a14150 & ~a14148;
assign a14154 = ~a13596 & ~a12268;
assign a14156 = ~a14154 & ~a14152;
assign a14158 = a13596 & a12268;
assign a14160 = ~a14158 & ~a14156;
assign a14162 = ~a13616 & ~a12080;
assign a14164 = ~a14162 & ~a14160;
assign a14166 = a13616 & a12080;
assign a14168 = ~a14166 & ~a14164;
assign a14170 = ~a13636 & ~a11820;
assign a14172 = ~a14170 & ~a14168;
assign a14174 = a13636 & a11820;
assign a14176 = ~a14174 & ~a14172;
assign a14178 = a13656 & a11202;
assign a14180 = ~a13656 & ~a11202;
assign a14182 = ~a14180 & ~a14178;
assign a14184 = ~a14182 & ~a14176;
assign a14186 = a13522 & a11292;
assign a14188 = ~a14186 & ~a14134;
assign a14190 = ~a14188 & ~a14130;
assign a14192 = ~a14190 & ~a14142;
assign a14194 = ~a14192 & ~a14138;
assign a14196 = ~a14194 & ~a14150;
assign a14198 = ~a14196 & ~a14146;
assign a14200 = ~a14198 & ~a14158;
assign a14202 = ~a14200 & ~a14154;
assign a14204 = ~a14202 & ~a14166;
assign a14206 = ~a14204 & ~a14162;
assign a14208 = ~a14206 & ~a14174;
assign a14210 = ~a14208 & ~a14170;
assign a14212 = ~a14210 & a14182;
assign a14214 = ~a14212 & ~a14184;
assign a14216 = a14048 & a13710;
assign a14218 = a14216 & ~a13708;
assign a14220 = a13636 & a11966;
assign a14222 = a13616 & a12162;
assign a14224 = ~a14222 & ~a14220;
assign a14226 = ~a13616 & ~a12162;
assign a14228 = ~a13596 & ~a12362;
assign a14230 = ~a14228 & ~a14226;
assign a14232 = a13596 & a12362;
assign a14234 = a13576 & a12562;
assign a14236 = ~a14234 & ~a14232;
assign a14238 = ~a13576 & ~a12562;
assign a14240 = a13556 & a12762;
assign a14242 = ~a13556 & ~a12762;
assign a14244 = a13536 & a12962;
assign a14246 = ~a13536 & ~a12962;
assign a14248 = ~a13522 & ~a13134;
assign a14250 = ~a14248 & ~a14246;
assign a14252 = ~a14250 & ~a14244;
assign a14254 = ~a14252 & ~a14242;
assign a14256 = ~a14254 & ~a14240;
assign a14258 = ~a14256 & ~a14238;
assign a14260 = ~a14258 & a14236;
assign a14262 = ~a14260 & a14230;
assign a14264 = ~a14262 & a14224;
assign a14266 = ~a13636 & ~a11966;
assign a14268 = ~a14266 & ~a14264;
assign a14270 = a13656 & a13312;
assign a14272 = ~a13656 & ~a13312;
assign a14274 = ~a14272 & ~a14270;
assign a14276 = ~a14274 & ~a14268;
assign a14278 = a14274 & a14268;
assign a14280 = ~a14278 & ~a14276;
assign a14282 = ~a14280 & a14126;
assign a14284 = ~a14282 & ~a14218;
assign a14286 = ~a14284 & ~a14214;
assign a14288 = a14286 & l1088;
assign a14290 = a14288 & a14126;
assign a14292 = ~a14290 & ~a14124;
assign a14294 = a14292 & a13956;
assign a14296 = ~a13522 & ~a11296;
assign a14298 = ~a13536 & ~a12872;
assign a14300 = ~a14298 & ~a14296;
assign a14302 = a13536 & a12872;
assign a14304 = ~a14302 & ~a14300;
assign a14306 = ~a13556 & ~a12672;
assign a14308 = ~a14306 & ~a14304;
assign a14310 = a13556 & a12672;
assign a14312 = ~a14310 & ~a14308;
assign a14314 = ~a13576 & ~a12472;
assign a14316 = ~a14314 & ~a14312;
assign a14318 = a13576 & a12472;
assign a14320 = ~a14318 & ~a14316;
assign a14322 = ~a13596 & ~a12272;
assign a14324 = ~a14322 & ~a14320;
assign a14326 = a13596 & a12272;
assign a14328 = ~a14326 & ~a14324;
assign a14330 = ~a13616 & ~a12084;
assign a14332 = ~a14330 & ~a14328;
assign a14334 = a13616 & a12084;
assign a14336 = ~a14334 & ~a14332;
assign a14338 = ~a13636 & ~a11824;
assign a14340 = ~a14338 & ~a14336;
assign a14342 = a13636 & a11824;
assign a14344 = ~a14342 & ~a14340;
assign a14346 = a13656 & a11206;
assign a14348 = ~a13656 & ~a11206;
assign a14350 = ~a14348 & ~a14346;
assign a14352 = ~a14350 & ~a14344;
assign a14354 = a13522 & a11296;
assign a14356 = ~a14354 & ~a14302;
assign a14358 = ~a14356 & ~a14298;
assign a14360 = ~a14358 & ~a14310;
assign a14362 = ~a14360 & ~a14306;
assign a14364 = ~a14362 & ~a14318;
assign a14366 = ~a14364 & ~a14314;
assign a14368 = ~a14366 & ~a14326;
assign a14370 = ~a14368 & ~a14322;
assign a14372 = ~a14370 & ~a14334;
assign a14374 = ~a14372 & ~a14330;
assign a14376 = ~a14374 & ~a14342;
assign a14378 = ~a14376 & ~a14338;
assign a14380 = ~a14378 & a14350;
assign a14382 = ~a14380 & ~a14352;
assign a14384 = a14216 & a13708;
assign a14386 = a13636 & a11970;
assign a14388 = ~a13636 & ~a11970;
assign a14390 = a13616 & a12166;
assign a14392 = ~a13616 & ~a12166;
assign a14394 = a13596 & a12366;
assign a14396 = ~a13596 & ~a12366;
assign a14398 = a13576 & a12566;
assign a14400 = ~a13576 & ~a12566;
assign a14402 = a13556 & a12766;
assign a14404 = ~a13556 & ~a12766;
assign a14406 = a13536 & a12966;
assign a14408 = ~a13536 & ~a12966;
assign a14410 = ~a13522 & ~a13138;
assign a14412 = ~a14410 & ~a14408;
assign a14414 = ~a14412 & ~a14406;
assign a14416 = ~a14414 & ~a14404;
assign a14418 = ~a14416 & ~a14402;
assign a14420 = ~a14418 & ~a14400;
assign a14422 = ~a14420 & ~a14398;
assign a14424 = ~a14422 & ~a14396;
assign a14426 = ~a14424 & ~a14394;
assign a14428 = ~a14426 & ~a14392;
assign a14430 = ~a14428 & ~a14390;
assign a14432 = ~a14430 & ~a14388;
assign a14434 = ~a14432 & ~a14386;
assign a14436 = a13656 & a13316;
assign a14438 = ~a13656 & ~a13316;
assign a14440 = ~a14438 & ~a14436;
assign a14442 = ~a14440 & a14434;
assign a14444 = a14440 & ~a14434;
assign a14446 = ~a14444 & ~a14442;
assign a14448 = ~a14446 & l584;
assign a14450 = a14448 & a13508;
assign a14452 = ~a14450 & ~a14384;
assign a14454 = ~a14452 & ~a14382;
assign a14456 = a14454 & l584;
assign a14458 = a13508 & l1086;
assign a14460 = a14458 & a14456;
assign a14462 = ~a14460 & a14294;
assign a14464 = a13508 & ~a5556;
assign a14466 = ~a13522 & ~a11328;
assign a14468 = ~a13536 & ~a12816;
assign a14470 = ~a14468 & ~a14466;
assign a14472 = a13536 & a12816;
assign a14474 = ~a14472 & ~a14470;
assign a14476 = ~a13556 & ~a12616;
assign a14478 = ~a14476 & ~a14474;
assign a14480 = a13556 & a12616;
assign a14482 = ~a14480 & ~a14478;
assign a14484 = ~a13576 & ~a12416;
assign a14486 = ~a14484 & ~a14482;
assign a14488 = a13576 & a12416;
assign a14490 = ~a14488 & ~a14486;
assign a14492 = ~a13596 & ~a12216;
assign a14494 = ~a14492 & ~a14490;
assign a14496 = a13596 & a12216;
assign a14498 = ~a14496 & ~a14494;
assign a14500 = ~a13616 & ~a12028;
assign a14502 = ~a14500 & ~a14498;
assign a14504 = a13616 & a12028;
assign a14506 = ~a14504 & ~a14502;
assign a14508 = ~a13636 & ~a11768;
assign a14510 = ~a14508 & ~a14506;
assign a14512 = a13636 & a11768;
assign a14514 = ~a14512 & ~a14510;
assign a14516 = a13656 & a11230;
assign a14518 = ~a13656 & ~a11230;
assign a14520 = ~a14518 & ~a14516;
assign a14522 = ~a14520 & ~a14514;
assign a14524 = a13522 & a11328;
assign a14526 = ~a14524 & ~a14472;
assign a14528 = ~a14526 & ~a14468;
assign a14530 = ~a14528 & ~a14480;
assign a14532 = ~a14530 & ~a14476;
assign a14534 = ~a14532 & ~a14488;
assign a14536 = ~a14534 & ~a14484;
assign a14538 = ~a14536 & ~a14496;
assign a14540 = ~a14538 & ~a14492;
assign a14542 = ~a14540 & ~a14504;
assign a14544 = ~a14542 & ~a14500;
assign a14546 = ~a14544 & ~a14512;
assign a14548 = ~a14546 & ~a14508;
assign a14550 = ~a14548 & a14520;
assign a14552 = ~a14550 & ~a14522;
assign a14554 = a14050 & a13702;
assign a14556 = a14554 & ~a13696;
assign a14558 = a13636 & a11918;
assign a14560 = a13616 & a12114;
assign a14562 = ~a14560 & ~a14558;
assign a14564 = ~a13616 & ~a12114;
assign a14566 = ~a13596 & ~a12314;
assign a14568 = ~a14566 & ~a14564;
assign a14570 = a13596 & a12314;
assign a14572 = a13576 & a12514;
assign a14574 = ~a14572 & ~a14570;
assign a14576 = ~a13576 & ~a12514;
assign a14578 = a13556 & a12714;
assign a14580 = ~a13556 & ~a12714;
assign a14582 = a13536 & a12914;
assign a14584 = ~a13536 & ~a12914;
assign a14586 = ~a13522 & ~a13086;
assign a14588 = ~a14586 & ~a14584;
assign a14590 = ~a14588 & ~a14582;
assign a14592 = ~a14590 & ~a14580;
assign a14594 = ~a14592 & ~a14578;
assign a14596 = ~a14594 & ~a14576;
assign a14598 = ~a14596 & a14574;
assign a14600 = ~a14598 & a14568;
assign a14602 = ~a14600 & a14562;
assign a14604 = ~a13636 & ~a11918;
assign a14606 = ~a14604 & ~a14602;
assign a14608 = a13656 & a13264;
assign a14610 = ~a13656 & ~a13264;
assign a14612 = ~a14610 & ~a14608;
assign a14614 = ~a14612 & ~a14606;
assign a14616 = a14612 & a14606;
assign a14618 = ~a14616 & ~a14614;
assign a14620 = ~a14618 & a14464;
assign a14622 = ~a14620 & ~a14556;
assign a14624 = ~a14622 & ~a14552;
assign a14626 = a14624 & l1104;
assign a14628 = a14626 & a14464;
assign a14630 = a13508 & ~a5548;
assign a14632 = ~a13522 & ~a11316;
assign a14634 = ~a13536 & ~a12804;
assign a14636 = ~a14634 & ~a14632;
assign a14638 = a13536 & a12804;
assign a14640 = ~a14638 & ~a14636;
assign a14642 = ~a13556 & ~a12604;
assign a14644 = ~a14642 & ~a14640;
assign a14646 = a13556 & a12604;
assign a14648 = ~a14646 & ~a14644;
assign a14650 = ~a13576 & ~a12404;
assign a14652 = ~a14650 & ~a14648;
assign a14654 = a13576 & a12404;
assign a14656 = ~a14654 & ~a14652;
assign a14658 = ~a13596 & ~a12204;
assign a14660 = ~a14658 & ~a14656;
assign a14662 = a13596 & a12204;
assign a14664 = ~a14662 & ~a14660;
assign a14666 = ~a13616 & ~a12016;
assign a14668 = ~a14666 & ~a14664;
assign a14670 = a13616 & a12016;
assign a14672 = ~a14670 & ~a14668;
assign a14674 = ~a13636 & ~a11756;
assign a14676 = ~a14674 & ~a14672;
assign a14678 = a13636 & a11756;
assign a14680 = ~a14678 & ~a14676;
assign a14682 = a13656 & a11222;
assign a14684 = ~a13656 & ~a11222;
assign a14686 = ~a14684 & ~a14682;
assign a14688 = ~a14686 & ~a14680;
assign a14690 = a13522 & a11316;
assign a14692 = ~a14690 & ~a14638;
assign a14694 = ~a14692 & ~a14634;
assign a14696 = ~a14694 & ~a14646;
assign a14698 = ~a14696 & ~a14642;
assign a14700 = ~a14698 & ~a14654;
assign a14702 = ~a14700 & ~a14650;
assign a14704 = ~a14702 & ~a14662;
assign a14706 = ~a14704 & ~a14658;
assign a14708 = ~a14706 & ~a14670;
assign a14710 = ~a14708 & ~a14666;
assign a14712 = ~a14710 & ~a14678;
assign a14714 = ~a14712 & ~a14674;
assign a14716 = ~a14714 & a14686;
assign a14718 = ~a14716 & ~a14688;
assign a14720 = a14048 & a13712;
assign a14722 = a13636 & a11910;
assign a14724 = a13616 & a12106;
assign a14726 = ~a14724 & ~a14722;
assign a14728 = ~a13616 & ~a12106;
assign a14730 = ~a13596 & ~a12306;
assign a14732 = ~a14730 & ~a14728;
assign a14734 = a13596 & a12306;
assign a14736 = a13576 & a12506;
assign a14738 = ~a14736 & ~a14734;
assign a14740 = ~a13576 & ~a12506;
assign a14742 = a13556 & a12706;
assign a14744 = ~a13556 & ~a12706;
assign a14746 = a13536 & a12906;
assign a14748 = ~a13536 & ~a12906;
assign a14750 = ~a13522 & ~a13078;
assign a14752 = ~a14750 & ~a14748;
assign a14754 = ~a14752 & ~a14746;
assign a14756 = ~a14754 & ~a14744;
assign a14758 = ~a14756 & ~a14742;
assign a14760 = ~a14758 & ~a14740;
assign a14762 = ~a14760 & a14738;
assign a14764 = ~a14762 & a14732;
assign a14766 = ~a14764 & a14726;
assign a14768 = ~a13636 & ~a11910;
assign a14770 = ~a14768 & ~a14766;
assign a14772 = a13656 & a13256;
assign a14774 = ~a13656 & ~a13256;
assign a14776 = ~a14774 & ~a14772;
assign a14778 = ~a14776 & ~a14770;
assign a14780 = a14776 & a14770;
assign a14782 = ~a14780 & ~a14778;
assign a14784 = ~a14782 & a14630;
assign a14786 = ~a14784 & ~a14720;
assign a14788 = ~a14786 & ~a14718;
assign a14790 = a14788 & ~a11850;
assign a14792 = a14790 & a14630;
assign a14794 = ~a14792 & ~a14628;
assign a14796 = a13508 & ~a5572;
assign a14798 = ~a13522 & ~a11336;
assign a14800 = ~a13536 & ~a12824;
assign a14802 = ~a14800 & ~a14798;
assign a14804 = a13536 & a12824;
assign a14806 = ~a14804 & ~a14802;
assign a14808 = ~a13556 & ~a12624;
assign a14810 = ~a14808 & ~a14806;
assign a14812 = a13556 & a12624;
assign a14814 = ~a14812 & ~a14810;
assign a14816 = ~a13576 & ~a12424;
assign a14818 = ~a14816 & ~a14814;
assign a14820 = a13576 & a12424;
assign a14822 = ~a14820 & ~a14818;
assign a14824 = ~a13596 & ~a12224;
assign a14826 = ~a14824 & ~a14822;
assign a14828 = a13596 & a12224;
assign a14830 = ~a14828 & ~a14826;
assign a14832 = ~a13616 & ~a12036;
assign a14834 = ~a14832 & ~a14830;
assign a14836 = a13616 & a12036;
assign a14838 = ~a14836 & ~a14834;
assign a14840 = ~a13636 & ~a11776;
assign a14842 = ~a14840 & ~a14838;
assign a14844 = a13636 & a11776;
assign a14846 = ~a14844 & ~a14842;
assign a14848 = a13656 & a11234;
assign a14850 = ~a13656 & ~a11234;
assign a14852 = ~a14850 & ~a14848;
assign a14854 = ~a14852 & ~a14846;
assign a14856 = a13522 & a11336;
assign a14858 = ~a14856 & ~a14804;
assign a14860 = ~a14858 & ~a14800;
assign a14862 = ~a14860 & ~a14812;
assign a14864 = ~a14862 & ~a14808;
assign a14866 = ~a14864 & ~a14820;
assign a14868 = ~a14866 & ~a14816;
assign a14870 = ~a14868 & ~a14828;
assign a14872 = ~a14870 & ~a14824;
assign a14874 = ~a14872 & ~a14836;
assign a14876 = ~a14874 & ~a14832;
assign a14878 = ~a14876 & ~a14844;
assign a14880 = ~a14878 & ~a14840;
assign a14882 = ~a14880 & a14852;
assign a14884 = ~a14882 & ~a14854;
assign a14886 = a13714 & ~a13696;
assign a14888 = a13636 & a11922;
assign a14890 = a13616 & a12118;
assign a14892 = ~a14890 & ~a14888;
assign a14894 = ~a13616 & ~a12118;
assign a14896 = ~a13596 & ~a12318;
assign a14898 = ~a14896 & ~a14894;
assign a14900 = a13596 & a12318;
assign a14902 = a13576 & a12518;
assign a14904 = ~a14902 & ~a14900;
assign a14906 = ~a13576 & ~a12518;
assign a14908 = a13556 & a12718;
assign a14910 = ~a13556 & ~a12718;
assign a14912 = a13536 & a12918;
assign a14914 = ~a13536 & ~a12918;
assign a14916 = ~a13522 & ~a13090;
assign a14918 = ~a14916 & ~a14914;
assign a14920 = ~a14918 & ~a14912;
assign a14922 = ~a14920 & ~a14910;
assign a14924 = ~a14922 & ~a14908;
assign a14926 = ~a14924 & ~a14906;
assign a14928 = ~a14926 & a14904;
assign a14930 = ~a14928 & a14898;
assign a14932 = ~a14930 & a14892;
assign a14934 = ~a13636 & ~a11922;
assign a14936 = ~a14934 & ~a14932;
assign a14938 = a13656 & a13268;
assign a14940 = ~a13656 & ~a13268;
assign a14942 = ~a14940 & ~a14938;
assign a14944 = ~a14942 & ~a14936;
assign a14946 = a14942 & a14936;
assign a14948 = ~a14946 & ~a14944;
assign a14950 = ~a14948 & a14796;
assign a14952 = ~a14950 & ~a14886;
assign a14954 = ~a14952 & ~a14884;
assign a14956 = a14954 & l1102;
assign a14958 = a14956 & a14796;
assign a14960 = ~a14958 & a14794;
assign a14962 = a13508 & l580;
assign a14964 = ~a13522 & ~a11360;
assign a14966 = ~a13536 & ~a12848;
assign a14968 = ~a14966 & ~a14964;
assign a14970 = a13536 & a12848;
assign a14972 = ~a14970 & ~a14968;
assign a14974 = ~a13556 & ~a12648;
assign a14976 = ~a14974 & ~a14972;
assign a14978 = a13556 & a12648;
assign a14980 = ~a14978 & ~a14976;
assign a14982 = ~a13576 & ~a12448;
assign a14984 = ~a14982 & ~a14980;
assign a14986 = a13576 & a12448;
assign a14988 = ~a14986 & ~a14984;
assign a14990 = ~a13596 & ~a12248;
assign a14992 = ~a14990 & ~a14988;
assign a14994 = a13596 & a12248;
assign a14996 = ~a14994 & ~a14992;
assign a14998 = ~a13616 & ~a12060;
assign a15000 = ~a14998 & ~a14996;
assign a15002 = a13616 & a12060;
assign a15004 = ~a15002 & ~a15000;
assign a15006 = ~a13636 & ~a11800;
assign a15008 = ~a15006 & ~a15004;
assign a15010 = a13636 & a11800;
assign a15012 = ~a15010 & ~a15008;
assign a15014 = a13656 & a11258;
assign a15016 = ~a13656 & ~a11258;
assign a15018 = ~a15016 & ~a15014;
assign a15020 = ~a15018 & ~a15012;
assign a15022 = a13522 & a11360;
assign a15024 = ~a15022 & ~a14970;
assign a15026 = ~a15024 & ~a14966;
assign a15028 = ~a15026 & ~a14978;
assign a15030 = ~a15028 & ~a14974;
assign a15032 = ~a15030 & ~a14986;
assign a15034 = ~a15032 & ~a14982;
assign a15036 = ~a15034 & ~a14994;
assign a15038 = ~a15036 & ~a14990;
assign a15040 = ~a15038 & ~a15002;
assign a15042 = ~a15040 & ~a14998;
assign a15044 = ~a15042 & ~a15010;
assign a15046 = ~a15044 & ~a15006;
assign a15048 = ~a15046 & a15018;
assign a15050 = ~a15048 & ~a15020;
assign a15052 = a14554 & a13696;
assign a15054 = a13636 & a11946;
assign a15056 = a13616 & a12142;
assign a15058 = ~a15056 & ~a15054;
assign a15060 = ~a13616 & ~a12142;
assign a15062 = ~a13596 & ~a12342;
assign a15064 = ~a15062 & ~a15060;
assign a15066 = a13596 & a12342;
assign a15068 = a13576 & a12542;
assign a15070 = ~a15068 & ~a15066;
assign a15072 = ~a13576 & ~a12542;
assign a15074 = a13556 & a12742;
assign a15076 = ~a13556 & ~a12742;
assign a15078 = a13536 & a12942;
assign a15080 = ~a13536 & ~a12942;
assign a15082 = ~a13522 & ~a13114;
assign a15084 = ~a15082 & ~a15080;
assign a15086 = ~a15084 & ~a15078;
assign a15088 = ~a15086 & ~a15076;
assign a15090 = ~a15088 & ~a15074;
assign a15092 = ~a15090 & ~a15072;
assign a15094 = ~a15092 & a15070;
assign a15096 = ~a15094 & a15064;
assign a15098 = ~a15096 & a15058;
assign a15100 = ~a13636 & ~a11946;
assign a15102 = ~a15100 & ~a15098;
assign a15104 = a13656 & a13292;
assign a15106 = ~a13656 & ~a13292;
assign a15108 = ~a15106 & ~a15104;
assign a15110 = ~a15108 & ~a15102;
assign a15112 = a15108 & a15102;
assign a15114 = ~a15112 & ~a15110;
assign a15116 = ~a15114 & a14962;
assign a15118 = ~a15116 & ~a15052;
assign a15120 = ~a15118 & ~a15050;
assign a15122 = a15120 & l1096;
assign a15124 = a15122 & a14962;
assign a15126 = a13508 & l576;
assign a15128 = ~a13522 & ~a11348;
assign a15130 = ~a13536 & ~a12836;
assign a15132 = ~a15130 & ~a15128;
assign a15134 = a13536 & a12836;
assign a15136 = ~a15134 & ~a15132;
assign a15138 = ~a13556 & ~a12636;
assign a15140 = ~a15138 & ~a15136;
assign a15142 = a13556 & a12636;
assign a15144 = ~a15142 & ~a15140;
assign a15146 = ~a13576 & ~a12436;
assign a15148 = ~a15146 & ~a15144;
assign a15150 = a13576 & a12436;
assign a15152 = ~a15150 & ~a15148;
assign a15154 = ~a13596 & ~a12236;
assign a15156 = ~a15154 & ~a15152;
assign a15158 = a13596 & a12236;
assign a15160 = ~a15158 & ~a15156;
assign a15162 = ~a13616 & ~a12048;
assign a15164 = ~a15162 & ~a15160;
assign a15166 = a13616 & a12048;
assign a15168 = ~a15166 & ~a15164;
assign a15170 = ~a13636 & ~a11788;
assign a15172 = ~a15170 & ~a15168;
assign a15174 = a13636 & a11788;
assign a15176 = ~a15174 & ~a15172;
assign a15178 = a13656 & a11246;
assign a15180 = ~a13656 & ~a11246;
assign a15182 = ~a15180 & ~a15178;
assign a15184 = ~a15182 & ~a15176;
assign a15186 = a13522 & a11348;
assign a15188 = ~a15186 & ~a15134;
assign a15190 = ~a15188 & ~a15130;
assign a15192 = ~a15190 & ~a15142;
assign a15194 = ~a15192 & ~a15138;
assign a15196 = ~a15194 & ~a15150;
assign a15198 = ~a15196 & ~a15146;
assign a15200 = ~a15198 & ~a15158;
assign a15202 = ~a15200 & ~a15154;
assign a15204 = ~a15202 & ~a15166;
assign a15206 = ~a15204 & ~a15162;
assign a15208 = ~a15206 & ~a15174;
assign a15210 = ~a15208 & ~a15170;
assign a15212 = ~a15210 & a15182;
assign a15214 = ~a15212 & ~a15184;
assign a15216 = a14050 & a13880;
assign a15218 = a13636 & a11934;
assign a15220 = a13616 & a12130;
assign a15222 = ~a15220 & ~a15218;
assign a15224 = ~a13616 & ~a12130;
assign a15226 = ~a13596 & ~a12330;
assign a15228 = ~a15226 & ~a15224;
assign a15230 = a13596 & a12330;
assign a15232 = a13576 & a12530;
assign a15234 = ~a15232 & ~a15230;
assign a15236 = ~a13576 & ~a12530;
assign a15238 = a13556 & a12730;
assign a15240 = ~a13556 & ~a12730;
assign a15242 = a13536 & a12930;
assign a15244 = ~a13536 & ~a12930;
assign a15246 = ~a13522 & ~a13102;
assign a15248 = ~a15246 & ~a15244;
assign a15250 = ~a15248 & ~a15242;
assign a15252 = ~a15250 & ~a15240;
assign a15254 = ~a15252 & ~a15238;
assign a15256 = ~a15254 & ~a15236;
assign a15258 = ~a15256 & a15234;
assign a15260 = ~a15258 & a15228;
assign a15262 = ~a15260 & a15222;
assign a15264 = ~a13636 & ~a11934;
assign a15266 = ~a15264 & ~a15262;
assign a15268 = a13656 & a13280;
assign a15270 = ~a13656 & ~a13280;
assign a15272 = ~a15270 & ~a15268;
assign a15274 = ~a15272 & ~a15266;
assign a15276 = a15272 & a15266;
assign a15278 = ~a15276 & ~a15274;
assign a15280 = ~a15278 & a15126;
assign a15282 = ~a15280 & ~a15216;
assign a15284 = ~a15282 & ~a15214;
assign a15286 = a15284 & l1100;
assign a15288 = a15286 & a15126;
assign a15290 = ~a15288 & ~a15124;
assign a15292 = a15290 & a14960;
assign a15294 = a15292 & a14462;
assign a15298 = ~a15296 & a11418;
assign a15300 = a15298 & ~l1470;
assign a15302 = a15300 & a10178;
assign a15304 = ~a10786 & a4544;
assign a15306 = a11432 & a10786;
assign a15308 = ~a15306 & ~a15304;
assign a15310 = ~a15308 & ~a15296;
assign a15312 = a15296 & a10178;
assign a15316 = ~a15314 & ~a15300;
assign a15318 = ~a15316 & ~a15302;
assign a15320 = l1686 & ~l950;
assign a15322 = a10766 & i210;
assign a15324 = ~a15322 & ~l1686;
assign a15326 = l1686 & l952;
assign a15328 = ~a15326 & ~a15324;
assign a15330 = l1686 & l956;
assign a15332 = ~a15330 & ~a15324;
assign a15334 = ~a15332 & ~l954;
assign a15336 = a15334 & ~a15328;
assign a15338 = a15336 & ~l958;
assign a15340 = a15338 & ~a15320;
assign a15342 = a15340 & ~a15318;
assign a15344 = a15322 & a3760;
assign a15346 = ~a15344 & ~l1686;
assign a15348 = l1686 & l1474;
assign a15350 = ~a15348 & ~a15346;
assign a15352 = a15350 & ~a15340;
assign a15354 = ~a15352 & ~a15342;
assign a15356 = a15354 & ~a11384;
assign a15358 = a15300 & a10152;
assign a15360 = ~a10786 & a4508;
assign a15362 = a11442 & a10786;
assign a15364 = ~a15362 & ~a15360;
assign a15366 = ~a15364 & ~a15296;
assign a15368 = a15296 & a10152;
assign a15372 = ~a15370 & ~a15300;
assign a15374 = ~a15372 & ~a15358;
assign a15376 = ~a15374 & a15340;
assign a15378 = a15322 & a4260;
assign a15380 = ~a15378 & ~l1686;
assign a15382 = l1686 & l1476;
assign a15384 = ~a15382 & ~a15380;
assign a15386 = a15384 & ~a15340;
assign a15388 = ~a15386 & ~a15376;
assign a15390 = ~a11532 & ~a11116;
assign a15392 = a12868 & ~a10920;
assign a15394 = a12872 & a10920;
assign a15396 = ~a15394 & ~a15392;
assign a15398 = ~a15396 & a11200;
assign a15400 = a12796 & a10966;
assign a15402 = ~a15400 & ~a15398;
assign a15404 = a12796 & ~a10920;
assign a15406 = a12804 & a10920;
assign a15408 = ~a15406 & ~a15404;
assign a15410 = ~a15408 & a10978;
assign a15412 = a12816 & ~a10920;
assign a15414 = a12824 & a10920;
assign a15416 = ~a15414 & ~a15412;
assign a15418 = ~a15416 & ~a10978;
assign a15420 = ~a15418 & ~a15410;
assign a15422 = ~a15420 & ~a10996;
assign a15424 = a12836 & ~a10920;
assign a15426 = a12840 & a10920;
assign a15428 = ~a15426 & ~a15424;
assign a15430 = ~a15428 & a10978;
assign a15432 = a12848 & ~a10920;
assign a15434 = a12852 & a10920;
assign a15436 = ~a15434 & ~a15432;
assign a15438 = ~a15436 & ~a10978;
assign a15440 = ~a15438 & ~a15430;
assign a15442 = ~a15440 & a10996;
assign a15444 = ~a15442 & ~a15422;
assign a15446 = ~a15444 & a11024;
assign a15450 = ~a15448 & a11116;
assign a15452 = ~a15450 & ~a15390;
assign a15454 = ~a15452 & a15388;
assign a15456 = ~a15454 & ~a15356;
assign a15458 = a15452 & ~a15388;
assign a15460 = ~a15458 & ~a15456;
assign a15462 = a15300 & a10126;
assign a15464 = ~a10786 & a4472;
assign a15466 = a11452 & a10786;
assign a15468 = ~a15466 & ~a15464;
assign a15470 = ~a15468 & ~a15296;
assign a15472 = a15296 & a10126;
assign a15476 = ~a15474 & ~a15300;
assign a15478 = ~a15476 & ~a15462;
assign a15480 = ~a15478 & a15340;
assign a15482 = a15322 & a4286;
assign a15484 = ~a15482 & ~l1686;
assign a15486 = l1686 & l1478;
assign a15488 = ~a15486 & ~a15484;
assign a15490 = a15488 & ~a15340;
assign a15492 = ~a15490 & ~a15480;
assign a15494 = ~a11552 & ~a11116;
assign a15496 = a12668 & ~a10920;
assign a15498 = a12672 & a10920;
assign a15500 = ~a15498 & ~a15496;
assign a15502 = ~a15500 & a11200;
assign a15504 = a12596 & a10966;
assign a15506 = ~a15504 & ~a15502;
assign a15508 = a12596 & ~a10920;
assign a15510 = a12604 & a10920;
assign a15512 = ~a15510 & ~a15508;
assign a15514 = ~a15512 & a10978;
assign a15516 = a12616 & ~a10920;
assign a15518 = a12624 & a10920;
assign a15520 = ~a15518 & ~a15516;
assign a15522 = ~a15520 & ~a10978;
assign a15524 = ~a15522 & ~a15514;
assign a15526 = ~a15524 & ~a10996;
assign a15528 = a12636 & ~a10920;
assign a15530 = a12640 & a10920;
assign a15532 = ~a15530 & ~a15528;
assign a15534 = ~a15532 & a10978;
assign a15536 = a12648 & ~a10920;
assign a15538 = a12652 & a10920;
assign a15540 = ~a15538 & ~a15536;
assign a15542 = ~a15540 & ~a10978;
assign a15544 = ~a15542 & ~a15534;
assign a15546 = ~a15544 & a10996;
assign a15548 = ~a15546 & ~a15526;
assign a15550 = ~a15548 & a11024;
assign a15554 = ~a15552 & a11116;
assign a15556 = ~a15554 & ~a15494;
assign a15558 = ~a15556 & a15492;
assign a15560 = ~a15558 & ~a15460;
assign a15562 = a15556 & ~a15492;
assign a15564 = ~a15562 & ~a15560;
assign a15566 = a15300 & a10100;
assign a15568 = ~a10786 & a4436;
assign a15570 = a11462 & a10786;
assign a15572 = ~a15570 & ~a15568;
assign a15574 = ~a15572 & ~a15296;
assign a15576 = a15296 & a10100;
assign a15580 = ~a15578 & ~a15300;
assign a15582 = ~a15580 & ~a15566;
assign a15584 = ~a15582 & a15340;
assign a15586 = a15322 & a4312;
assign a15588 = ~a15586 & ~l1686;
assign a15590 = l1686 & l1480;
assign a15592 = ~a15590 & ~a15588;
assign a15594 = a15592 & ~a15340;
assign a15596 = ~a15594 & ~a15584;
assign a15598 = ~a11566 & ~a11116;
assign a15600 = a12468 & ~a10920;
assign a15602 = a12472 & a10920;
assign a15604 = ~a15602 & ~a15600;
assign a15606 = ~a15604 & a11200;
assign a15608 = a12396 & a10966;
assign a15610 = ~a15608 & ~a15606;
assign a15612 = a12396 & ~a10920;
assign a15614 = a12404 & a10920;
assign a15616 = ~a15614 & ~a15612;
assign a15618 = ~a15616 & a10978;
assign a15620 = a12416 & ~a10920;
assign a15622 = a12424 & a10920;
assign a15624 = ~a15622 & ~a15620;
assign a15626 = ~a15624 & ~a10978;
assign a15628 = ~a15626 & ~a15618;
assign a15630 = ~a15628 & ~a10996;
assign a15632 = a12436 & ~a10920;
assign a15634 = a12440 & a10920;
assign a15636 = ~a15634 & ~a15632;
assign a15638 = ~a15636 & a10978;
assign a15640 = a12448 & ~a10920;
assign a15642 = a12452 & a10920;
assign a15644 = ~a15642 & ~a15640;
assign a15646 = ~a15644 & ~a10978;
assign a15648 = ~a15646 & ~a15638;
assign a15650 = ~a15648 & a10996;
assign a15652 = ~a15650 & ~a15630;
assign a15654 = ~a15652 & a11024;
assign a15658 = ~a15656 & a11116;
assign a15660 = ~a15658 & ~a15598;
assign a15662 = ~a15660 & a15596;
assign a15664 = ~a15662 & ~a15564;
assign a15666 = a15660 & ~a15596;
assign a15668 = ~a15666 & ~a15664;
assign a15670 = a15300 & a10074;
assign a15672 = ~a10786 & a4398;
assign a15674 = a11472 & a10786;
assign a15676 = ~a15674 & ~a15672;
assign a15678 = ~a15676 & ~a15296;
assign a15680 = a15296 & a10074;
assign a15684 = ~a15682 & ~a15300;
assign a15686 = ~a15684 & ~a15670;
assign a15688 = ~a15686 & a15340;
assign a15690 = a15322 & a3758;
assign a15692 = ~a15690 & ~l1686;
assign a15694 = l1686 & l1482;
assign a15696 = ~a15694 & ~a15692;
assign a15698 = a15696 & ~a15340;
assign a15700 = ~a15698 & ~a15688;
assign a15702 = ~a11580 & ~a11116;
assign a15704 = a12268 & ~a10920;
assign a15706 = a12272 & a10920;
assign a15708 = ~a15706 & ~a15704;
assign a15710 = ~a15708 & a11200;
assign a15712 = a12196 & a10966;
assign a15714 = ~a15712 & ~a15710;
assign a15716 = a12196 & ~a10920;
assign a15718 = a12204 & a10920;
assign a15720 = ~a15718 & ~a15716;
assign a15722 = ~a15720 & a10978;
assign a15724 = a12216 & ~a10920;
assign a15726 = a12224 & a10920;
assign a15728 = ~a15726 & ~a15724;
assign a15730 = ~a15728 & ~a10978;
assign a15732 = ~a15730 & ~a15722;
assign a15734 = ~a15732 & ~a10996;
assign a15736 = a12236 & ~a10920;
assign a15738 = a12240 & a10920;
assign a15740 = ~a15738 & ~a15736;
assign a15742 = ~a15740 & a10978;
assign a15744 = a12248 & ~a10920;
assign a15746 = a12252 & a10920;
assign a15748 = ~a15746 & ~a15744;
assign a15750 = ~a15748 & ~a10978;
assign a15752 = ~a15750 & ~a15742;
assign a15754 = ~a15752 & a10996;
assign a15756 = ~a15754 & ~a15734;
assign a15758 = ~a15756 & a11024;
assign a15762 = ~a15760 & a11116;
assign a15764 = ~a15762 & ~a15702;
assign a15766 = ~a15764 & a15700;
assign a15768 = ~a15766 & ~a15668;
assign a15770 = a15764 & ~a15700;
assign a15772 = ~a15770 & ~a15768;
assign a15774 = a15300 & a10044;
assign a15776 = ~a10786 & a2542;
assign a15778 = a11478 & a10786;
assign a15780 = ~a15778 & ~a15776;
assign a15782 = ~a15780 & ~a15296;
assign a15784 = a15296 & a10044;
assign a15788 = ~a15786 & ~a15300;
assign a15790 = ~a15788 & ~a15774;
assign a15792 = ~a15790 & a15340;
assign a15794 = l1686 & ~l1484;
assign a15796 = a15794 & ~a15340;
assign a15798 = ~a15796 & ~a15792;
assign a15800 = ~a11594 & ~a11116;
assign a15802 = a12080 & ~a10920;
assign a15804 = a12084 & a10920;
assign a15806 = ~a15804 & ~a15802;
assign a15808 = ~a15806 & a11200;
assign a15810 = a12008 & a10966;
assign a15812 = ~a15810 & ~a15808;
assign a15814 = a12008 & ~a10920;
assign a15816 = a12016 & a10920;
assign a15818 = ~a15816 & ~a15814;
assign a15820 = ~a15818 & a10978;
assign a15822 = a12028 & ~a10920;
assign a15824 = a12036 & a10920;
assign a15826 = ~a15824 & ~a15822;
assign a15828 = ~a15826 & ~a10978;
assign a15830 = ~a15828 & ~a15820;
assign a15832 = ~a15830 & ~a10996;
assign a15834 = a12048 & ~a10920;
assign a15836 = a12052 & a10920;
assign a15838 = ~a15836 & ~a15834;
assign a15840 = ~a15838 & a10978;
assign a15842 = a12060 & ~a10920;
assign a15844 = a12064 & a10920;
assign a15846 = ~a15844 & ~a15842;
assign a15848 = ~a15846 & ~a10978;
assign a15850 = ~a15848 & ~a15840;
assign a15852 = ~a15850 & a10996;
assign a15854 = ~a15852 & ~a15832;
assign a15856 = ~a15854 & a11024;
assign a15860 = ~a15858 & a11116;
assign a15862 = ~a15860 & ~a15800;
assign a15864 = ~a15862 & a15798;
assign a15866 = ~a15864 & ~a15772;
assign a15868 = a15862 & ~a15798;
assign a15870 = ~a15868 & ~a15866;
assign a15872 = a15300 & a8874;
assign a15874 = ~a10786 & a2526;
assign a15876 = a11486 & a10786;
assign a15878 = ~a15876 & ~a15874;
assign a15880 = ~a15878 & ~a15296;
assign a15882 = a15296 & a8874;
assign a15886 = ~a15884 & ~a15300;
assign a15888 = ~a15886 & ~a15872;
assign a15890 = ~a15888 & a15340;
assign a15892 = l1686 & ~l1486;
assign a15894 = a15892 & ~a15340;
assign a15896 = ~a15894 & ~a15890;
assign a15898 = ~a11608 & ~a11116;
assign a15900 = a11820 & ~a10920;
assign a15902 = a11824 & a10920;
assign a15904 = ~a15902 & ~a15900;
assign a15906 = ~a15904 & a11200;
assign a15908 = a11752 & a10966;
assign a15910 = ~a15908 & ~a15906;
assign a15912 = a11752 & ~a10920;
assign a15914 = a11756 & a10920;
assign a15916 = ~a15914 & ~a15912;
assign a15918 = ~a15916 & a10978;
assign a15920 = a11768 & ~a10920;
assign a15922 = a11776 & a10920;
assign a15924 = ~a15922 & ~a15920;
assign a15926 = ~a15924 & ~a10978;
assign a15928 = ~a15926 & ~a15918;
assign a15930 = ~a15928 & ~a10996;
assign a15932 = a11788 & ~a10920;
assign a15934 = a11792 & a10920;
assign a15936 = ~a15934 & ~a15932;
assign a15938 = ~a15936 & a10978;
assign a15940 = a11800 & ~a10920;
assign a15942 = a11804 & a10920;
assign a15944 = ~a15942 & ~a15940;
assign a15946 = ~a15944 & ~a10978;
assign a15948 = ~a15946 & ~a15938;
assign a15950 = ~a15948 & a10996;
assign a15952 = ~a15950 & ~a15930;
assign a15954 = ~a15952 & a11024;
assign a15958 = ~a15956 & a11116;
assign a15960 = ~a15958 & ~a15898;
assign a15962 = ~a15960 & a15896;
assign a15964 = ~a15962 & ~a15870;
assign a15966 = a15960 & ~a15896;
assign a15968 = ~a15966 & ~a15964;
assign a15970 = a15300 & a8868;
assign a15972 = ~a10786 & a2266;
assign a15974 = a11490 & a10786;
assign a15976 = ~a15974 & ~a15972;
assign a15978 = ~a15976 & ~a15296;
assign a15980 = a15296 & a8868;
assign a15984 = ~a15982 & ~a15300;
assign a15986 = ~a15984 & ~a15970;
assign a15988 = ~a15986 & a15340;
assign a15990 = l1686 & ~l960;
assign a15992 = a15990 & ~a15340;
assign a15994 = ~a15992 & ~a15988;
assign a15996 = ~a15994 & a11282;
assign a15998 = a15994 & ~a11282;
assign a16000 = ~a15998 & ~a15996;
assign a16002 = ~a16000 & ~a15968;
assign a16004 = ~a15354 & a11384;
assign a16006 = ~a16004 & ~a15458;
assign a16008 = ~a16006 & ~a15454;
assign a16010 = ~a16008 & ~a15562;
assign a16012 = ~a16010 & ~a15558;
assign a16014 = ~a16012 & ~a15666;
assign a16016 = ~a16014 & ~a15662;
assign a16018 = ~a16016 & ~a15770;
assign a16020 = ~a16018 & ~a15766;
assign a16022 = ~a16020 & ~a15868;
assign a16024 = ~a16022 & ~a15864;
assign a16026 = ~a16024 & ~a15966;
assign a16028 = ~a16026 & ~a15962;
assign a16030 = ~a16028 & a16000;
assign a16032 = ~a16030 & ~a16002;
assign a16034 = a16032 & ~a11282;
assign a16036 = ~a16032 & ~a15994;
assign a16038 = ~a16036 & ~a16034;
assign a16040 = ~a16038 & ~a8044;
assign a16042 = ~a8042 & ~i350;
assign a16044 = ~a16042 & a16038;
assign a16046 = ~a16044 & ~a16040;
assign a16048 = ~a7928 & ~l724;
assign a16050 = ~a16048 & ~a6908;
assign a16052 = ~a16050 & ~a7940;
assign a16054 = ~a16052 & ~i348;
assign a16056 = ~a16054 & ~a16042;
assign a16058 = a16056 & ~a8044;
assign a16060 = a16052 & i348;
assign a16062 = l1686 & ~l746;
assign a16064 = a16062 & ~l494;
assign a16066 = ~a16064 & ~a7850;
assign a16068 = ~a16066 & ~a6908;
assign a16072 = ~a16070 & ~i346;
assign a16074 = a16070 & i346;
assign a16076 = ~a7810 & ~l768;
assign a16078 = ~a16076 & ~a6908;
assign a16080 = ~a16078 & ~a7964;
assign a16082 = ~a16080 & ~i344;
assign a16084 = a16080 & i344;
assign a16086 = ~a7588 & ~l790;
assign a16088 = ~a16086 & ~a6908;
assign a16090 = ~a16088 & ~a7976;
assign a16092 = ~a16090 & ~i342;
assign a16094 = a16090 & i342;
assign a16096 = ~a7350 & ~l812;
assign a16098 = ~a16096 & ~a6908;
assign a16100 = ~a16098 & ~a7988;
assign a16102 = ~a16100 & ~i340;
assign a16104 = a16100 & i340;
assign a16106 = ~a7150 & ~l834;
assign a16108 = ~a16106 & ~a6908;
assign a16110 = ~a16108 & ~a6918;
assign a16112 = ~a16110 & ~i338;
assign a16114 = a16110 & i338;
assign a16116 = ~a8018 & ~l856;
assign a16118 = ~a16116 & ~a6908;
assign a16120 = ~a16118 & ~a8000;
assign a16122 = a16120 & i336;
assign a16124 = ~a16122 & ~a16114;
assign a16126 = ~a16124 & ~a16112;
assign a16128 = ~a16126 & ~a16104;
assign a16130 = ~a16128 & ~a16102;
assign a16132 = ~a16130 & ~a16094;
assign a16134 = ~a16132 & ~a16092;
assign a16136 = ~a16134 & ~a16084;
assign a16138 = ~a16136 & ~a16082;
assign a16140 = ~a16138 & ~a16074;
assign a16142 = ~a16140 & ~a16072;
assign a16144 = ~a16142 & ~a16060;
assign a16146 = ~a16144 & a16058;
assign a16148 = ~a16146 & ~a16046;
assign a16150 = a16032 & ~a15960;
assign a16152 = ~a16032 & ~a15896;
assign a16154 = ~a16152 & ~a16150;
assign a16156 = a16154 & i348;
assign a16158 = ~a16156 & ~a16148;
assign a16160 = ~a16154 & ~i348;
assign a16162 = a16032 & ~a15862;
assign a16164 = ~a16032 & ~a15798;
assign a16166 = ~a16164 & ~a16162;
assign a16168 = a16166 & i346;
assign a16170 = ~a16166 & ~i346;
assign a16172 = a16032 & ~a15764;
assign a16174 = ~a16032 & ~a15700;
assign a16176 = ~a16174 & ~a16172;
assign a16178 = a16176 & i344;
assign a16180 = ~a16176 & ~i344;
assign a16182 = a16032 & ~a15660;
assign a16184 = ~a16032 & ~a15596;
assign a16186 = ~a16184 & ~a16182;
assign a16188 = a16186 & i342;
assign a16190 = ~a16186 & ~i342;
assign a16192 = a16032 & ~a15556;
assign a16194 = ~a16032 & ~a15492;
assign a16196 = ~a16194 & ~a16192;
assign a16198 = a16196 & i340;
assign a16200 = ~a16196 & ~i340;
assign a16202 = a16032 & ~a15452;
assign a16204 = ~a16032 & ~a15388;
assign a16206 = ~a16204 & ~a16202;
assign a16208 = a16206 & i338;
assign a16210 = ~a16206 & ~i338;
assign a16212 = a16032 & ~a11384;
assign a16214 = ~a16032 & ~a15354;
assign a16216 = ~a16214 & ~a16212;
assign a16218 = ~a16216 & ~i336;
assign a16220 = ~a16218 & ~a16210;
assign a16222 = ~a16220 & ~a16208;
assign a16224 = ~a16222 & ~a16200;
assign a16226 = ~a16224 & ~a16198;
assign a16228 = ~a16226 & ~a16190;
assign a16230 = ~a16228 & ~a16188;
assign a16232 = ~a16230 & ~a16180;
assign a16234 = ~a16232 & ~a16178;
assign a16236 = ~a16234 & ~a16170;
assign a16238 = ~a16236 & ~a16168;
assign a16240 = ~a16238 & ~a16160;
assign a16242 = ~a16240 & a16158;
assign a16244 = ~a16038 & a8042;
assign a16246 = a16038 & ~a8042;
assign a16248 = ~a16246 & ~a16244;
assign a16250 = ~a16248 & a16146;
assign a16252 = ~a16250 & ~a16242;
assign a16254 = ~l948 & ~l946;
assign a16256 = a16254 & a6674;
assign a16258 = a16256 & ~a16252;
assign a16260 = a16258 & ~a8032;
assign a16262 = a16260 & a8022;
assign a16264 = ~a16262 & a5368;
assign a16266 = a16262 & i338;
assign a16270 = ~a16262 & a5376;
assign a16272 = a16262 & i340;
assign a16276 = ~a16262 & a5384;
assign a16278 = a16262 & i342;
assign a16282 = ~a16262 & a5392;
assign a16284 = a16262 & i344;
assign a16288 = ~a16262 & a5394;
assign a16290 = a16262 & i346;
assign a16294 = ~a16262 & a5396;
assign a16296 = a16262 & i348;
assign a16300 = ~a16262 & a5398;
assign a16302 = a16262 & i350;
assign a16306 = ~a16262 & a5514;
assign a16308 = a16262 & i336;
assign a16312 = l1686 & ~l1504;
assign a16314 = l1686 & ~l1530;
assign a16316 = a2246 & i166;
assign a16318 = ~a2246 & a1746;
assign a16320 = ~a16318 & ~a16316;
assign a16322 = a2246 & i164;
assign a16324 = ~a2246 & a1726;
assign a16326 = ~a16324 & ~a16322;
assign a16328 = a16326 & a16320;
assign a16330 = a2246 & i162;
assign a16332 = ~a2246 & a1694;
assign a16334 = ~a16332 & ~a16330;
assign a16336 = a16334 & a16328;
assign a16338 = a2246 & i160;
assign a16340 = ~a16338 & ~a6502;
assign a16342 = ~a16340 & a6934;
assign a16344 = a16342 & a16336;
assign a16346 = ~a16344 & a16314;
assign a16348 = a2246 & i158;
assign a16350 = ~a2246 & a1692;
assign a16352 = ~a16350 & ~a16348;
assign a16354 = ~a16352 & a16344;
assign a16358 = a16356 & a16312;
assign a16360 = ~a16356 & ~a16312;
assign a16362 = ~a16360 & ~a16358;
assign a16364 = ~a11316 & ~a7998;
assign a16366 = ~a12804 & ~a6916;
assign a16368 = ~a16366 & ~a16364;
assign a16370 = a12804 & a6916;
assign a16372 = ~a16370 & ~a16368;
assign a16374 = ~a12604 & ~a7986;
assign a16376 = ~a16374 & ~a16372;
assign a16378 = a12604 & a7986;
assign a16380 = ~a16378 & ~a16376;
assign a16382 = ~a12404 & ~a7974;
assign a16384 = ~a16382 & ~a16380;
assign a16386 = a12404 & a7974;
assign a16388 = ~a16386 & ~a16384;
assign a16390 = ~a12204 & ~a7962;
assign a16392 = ~a16390 & ~a16388;
assign a16394 = a12204 & a7962;
assign a16396 = ~a16394 & ~a16392;
assign a16398 = ~a12016 & ~a7950;
assign a16400 = ~a16398 & ~a16396;
assign a16402 = a12016 & a7950;
assign a16404 = ~a16402 & ~a16400;
assign a16406 = ~a11756 & ~a7938;
assign a16408 = ~a16406 & ~a16404;
assign a16410 = a11756 & a7938;
assign a16412 = ~a16410 & ~a16408;
assign a16414 = a11222 & a7860;
assign a16416 = ~a11222 & ~a7860;
assign a16418 = ~a16416 & ~a16414;
assign a16420 = ~a16418 & ~a16412;
assign a16422 = a11316 & a7998;
assign a16424 = ~a16422 & ~a16370;
assign a16426 = ~a16424 & ~a16366;
assign a16428 = ~a16426 & ~a16378;
assign a16430 = ~a16428 & ~a16374;
assign a16432 = ~a16430 & ~a16386;
assign a16434 = ~a16432 & ~a16382;
assign a16436 = ~a16434 & ~a16394;
assign a16438 = ~a16436 & ~a16390;
assign a16440 = ~a16438 & ~a16402;
assign a16442 = ~a16440 & ~a16398;
assign a16444 = ~a16442 & ~a16410;
assign a16446 = ~a16444 & ~a16406;
assign a16448 = ~a16446 & a16418;
assign a16450 = ~a16448 & ~a16420;
assign a16452 = ~a16450 & a16362;
assign a16454 = a16452 & a6908;
assign a16456 = a16454 & ~a5548;
assign a16458 = ~a16456 & ~a5542;
assign a16460 = a16336 & a6934;
assign a16462 = a16460 & a16340;
assign a16464 = ~a16462 & ~a16458;
assign a16466 = ~a16464 & ~l494;
assign a16468 = a16312 & ~a13708;
assign a16470 = a16314 & a13708;
assign a16472 = ~a16470 & ~a16468;
assign a16474 = ~a16472 & ~a13702;
assign a16476 = l1686 & ~l1528;
assign a16478 = a16476 & ~a13708;
assign a16480 = l1686 & ~l1526;
assign a16482 = a16480 & a13708;
assign a16484 = ~a16482 & ~a16478;
assign a16486 = ~a16484 & a13702;
assign a16488 = ~a16486 & ~a16474;
assign a16490 = ~a16488 & ~a13696;
assign a16492 = l1686 & ~l1524;
assign a16494 = a16492 & ~a13708;
assign a16496 = l1686 & ~l1522;
assign a16498 = a16496 & a13708;
assign a16500 = ~a16498 & ~a16494;
assign a16502 = ~a16500 & ~a13702;
assign a16504 = l1686 & ~l1520;
assign a16506 = a16504 & ~a13708;
assign a16508 = l1686 & ~l1518;
assign a16510 = a16508 & a13708;
assign a16512 = ~a16510 & ~a16506;
assign a16514 = ~a16512 & a13702;
assign a16516 = ~a16514 & ~a16502;
assign a16518 = ~a16516 & a13696;
assign a16520 = ~a16518 & ~a16490;
assign a16522 = ~a16520 & ~a13710;
assign a16524 = l1686 & ~l1516;
assign a16526 = a16524 & ~a13708;
assign a16528 = l1686 & ~l1514;
assign a16530 = a16528 & a13708;
assign a16532 = ~a16530 & ~a16526;
assign a16534 = ~a16532 & a13710;
assign a16536 = ~a16534 & ~a16522;
assign a16538 = ~a16536 & a6424;
assign a16540 = a16536 & ~a6424;
assign a16542 = ~a16540 & ~a16538;
assign a16544 = l1686 & ~l1508;
assign a16546 = a16544 & a6548;
assign a16548 = l1686 & ~l1512;
assign a16550 = ~a16548 & ~a6512;
assign a16552 = ~a16550 & ~a16546;
assign a16554 = l1686 & ~l1510;
assign a16556 = a16554 & a6592;
assign a16558 = a16548 & a6512;
assign a16560 = ~a16558 & ~a16556;
assign a16562 = a16560 & a16552;
assign a16564 = ~a16554 & ~a6592;
assign a16566 = ~a16544 & ~a6548;
assign a16568 = ~a16566 & ~a16564;
assign a16570 = l1686 & ~l1506;
assign a16572 = a16570 & a6476;
assign a16574 = ~a16570 & ~a6476;
assign a16576 = ~a16574 & ~a16572;
assign a16578 = a16576 & a16568;
assign a16580 = a16578 & a16562;
assign a16582 = ~a16580 & ~a16542;
assign a16584 = a6512 & ~a5542;
assign a16586 = ~a6512 & ~a5548;
assign a16588 = ~a16586 & ~a16584;
assign a16590 = ~a16588 & a6548;
assign a16592 = a6512 & ~a5556;
assign a16594 = ~a6512 & ~a5572;
assign a16596 = ~a16594 & ~a16592;
assign a16598 = ~a16596 & ~a6548;
assign a16600 = ~a16598 & ~a16590;
assign a16602 = ~a16600 & a6592;
assign a16604 = a6512 & l576;
assign a16606 = ~a6512 & l578;
assign a16608 = ~a16606 & ~a16604;
assign a16610 = ~a16608 & a6548;
assign a16612 = a6512 & l580;
assign a16614 = ~a6512 & l582;
assign a16616 = ~a16614 & ~a16612;
assign a16618 = ~a16616 & ~a6548;
assign a16620 = ~a16618 & ~a16610;
assign a16622 = ~a16620 & ~a6592;
assign a16624 = ~a16622 & ~a16602;
assign a16626 = ~a16624 & a6476;
assign a16628 = a6512 & l586;
assign a16630 = ~a6512 & l584;
assign a16632 = ~a16630 & ~a16628;
assign a16634 = ~a16632 & ~a6476;
assign a16636 = ~a16634 & ~a16626;
assign a16638 = ~a16636 & a16582;
assign a16640 = a16312 & a6424;
assign a16642 = ~a16312 & ~a6424;
assign a16644 = ~a16642 & ~a16640;
assign a16646 = ~a16644 & a16638;
assign a16648 = a6548 & a6512;
assign a16650 = a16648 & a6592;
assign a16652 = a16650 & a6476;
assign a16654 = a16652 & a16644;
assign a16656 = ~a16654 & ~a16646;
assign a16658 = ~a16656 & a1690;
assign a16662 = a16334 & a16326;
assign a16664 = ~a16320 & a6934;
assign a16666 = a16664 & a16662;
assign a16668 = a16666 & a16340;
assign a16670 = ~a16668 & a16476;
assign a16672 = a16668 & ~a16352;
assign a16676 = a16674 & a16314;
assign a16678 = ~a16674 & ~a16314;
assign a16680 = ~a16678 & ~a16676;
assign a16682 = ~a11328 & ~a7998;
assign a16684 = ~a12816 & ~a6916;
assign a16686 = ~a16684 & ~a16682;
assign a16688 = a12816 & a6916;
assign a16690 = ~a16688 & ~a16686;
assign a16692 = ~a12616 & ~a7986;
assign a16694 = ~a16692 & ~a16690;
assign a16696 = a12616 & a7986;
assign a16698 = ~a16696 & ~a16694;
assign a16700 = ~a12416 & ~a7974;
assign a16702 = ~a16700 & ~a16698;
assign a16704 = a12416 & a7974;
assign a16706 = ~a16704 & ~a16702;
assign a16708 = ~a12216 & ~a7962;
assign a16710 = ~a16708 & ~a16706;
assign a16712 = a12216 & a7962;
assign a16714 = ~a16712 & ~a16710;
assign a16716 = ~a12028 & ~a7950;
assign a16718 = ~a16716 & ~a16714;
assign a16720 = a12028 & a7950;
assign a16722 = ~a16720 & ~a16718;
assign a16724 = ~a11768 & ~a7938;
assign a16726 = ~a16724 & ~a16722;
assign a16728 = a11768 & a7938;
assign a16730 = ~a16728 & ~a16726;
assign a16732 = a11230 & a7860;
assign a16734 = ~a11230 & ~a7860;
assign a16736 = ~a16734 & ~a16732;
assign a16738 = ~a16736 & ~a16730;
assign a16740 = a11328 & a7998;
assign a16742 = ~a16740 & ~a16688;
assign a16744 = ~a16742 & ~a16684;
assign a16746 = ~a16744 & ~a16696;
assign a16748 = ~a16746 & ~a16692;
assign a16750 = ~a16748 & ~a16704;
assign a16752 = ~a16750 & ~a16700;
assign a16754 = ~a16752 & ~a16712;
assign a16756 = ~a16754 & ~a16708;
assign a16758 = ~a16756 & ~a16720;
assign a16760 = ~a16758 & ~a16716;
assign a16762 = ~a16760 & ~a16728;
assign a16764 = ~a16762 & ~a16724;
assign a16766 = ~a16764 & a16736;
assign a16768 = ~a16766 & ~a16738;
assign a16770 = ~a16768 & a16680;
assign a16772 = a16770 & a6908;
assign a16774 = a16772 & ~a5556;
assign a16776 = ~a16774 & ~a5548;
assign a16778 = ~a16776 & ~a16344;
assign a16780 = ~a16778 & ~l494;
assign a16782 = a16314 & a6424;
assign a16784 = ~a16314 & ~a6424;
assign a16786 = ~a16784 & ~a16782;
assign a16788 = ~a16786 & a16638;
assign a16790 = a6592 & a6548;
assign a16792 = a16790 & a6476;
assign a16794 = a16792 & a16786;
assign a16796 = ~a16794 & ~a16788;
assign a16798 = ~a16796 & a1690;
assign a16802 = a16666 & ~a16340;
assign a16804 = ~a16802 & a16480;
assign a16806 = a16802 & ~a16352;
assign a16810 = a16808 & a16476;
assign a16812 = ~a16808 & ~a16476;
assign a16814 = ~a16812 & ~a16810;
assign a16816 = ~a11336 & ~a7998;
assign a16818 = ~a12824 & ~a6916;
assign a16820 = ~a16818 & ~a16816;
assign a16822 = a12824 & a6916;
assign a16824 = ~a16822 & ~a16820;
assign a16826 = ~a12624 & ~a7986;
assign a16828 = ~a16826 & ~a16824;
assign a16830 = a12624 & a7986;
assign a16832 = ~a16830 & ~a16828;
assign a16834 = ~a12424 & ~a7974;
assign a16836 = ~a16834 & ~a16832;
assign a16838 = a12424 & a7974;
assign a16840 = ~a16838 & ~a16836;
assign a16842 = ~a12224 & ~a7962;
assign a16844 = ~a16842 & ~a16840;
assign a16846 = a12224 & a7962;
assign a16848 = ~a16846 & ~a16844;
assign a16850 = ~a12036 & ~a7950;
assign a16852 = ~a16850 & ~a16848;
assign a16854 = a12036 & a7950;
assign a16856 = ~a16854 & ~a16852;
assign a16858 = ~a11776 & ~a7938;
assign a16860 = ~a16858 & ~a16856;
assign a16862 = a11776 & a7938;
assign a16864 = ~a16862 & ~a16860;
assign a16866 = a11234 & a7860;
assign a16868 = ~a11234 & ~a7860;
assign a16870 = ~a16868 & ~a16866;
assign a16872 = ~a16870 & ~a16864;
assign a16874 = a11336 & a7998;
assign a16876 = ~a16874 & ~a16822;
assign a16878 = ~a16876 & ~a16818;
assign a16880 = ~a16878 & ~a16830;
assign a16882 = ~a16880 & ~a16826;
assign a16884 = ~a16882 & ~a16838;
assign a16886 = ~a16884 & ~a16834;
assign a16888 = ~a16886 & ~a16846;
assign a16890 = ~a16888 & ~a16842;
assign a16892 = ~a16890 & ~a16854;
assign a16894 = ~a16892 & ~a16850;
assign a16896 = ~a16894 & ~a16862;
assign a16898 = ~a16896 & ~a16858;
assign a16900 = ~a16898 & a16870;
assign a16902 = ~a16900 & ~a16872;
assign a16904 = ~a16902 & a16814;
assign a16906 = a16904 & a6908;
assign a16908 = a16906 & ~a5572;
assign a16910 = ~a16908 & ~a5556;
assign a16912 = ~a16910 & ~a16668;
assign a16914 = ~a16912 & ~l494;
assign a16916 = a16476 & a6424;
assign a16918 = ~a16476 & ~a6424;
assign a16920 = ~a16918 & ~a16916;
assign a16922 = ~a16920 & a16638;
assign a16924 = a6592 & a6476;
assign a16926 = ~a6548 & ~a6512;
assign a16928 = ~a16926 & a16924;
assign a16930 = a16928 & a16920;
assign a16932 = ~a16930 & ~a16922;
assign a16934 = ~a16932 & a1690;
assign a16938 = ~a16326 & a6934;
assign a16940 = a16938 & a16334;
assign a16942 = a16940 & a16340;
assign a16944 = a16942 & a16320;
assign a16946 = ~a16944 & a16492;
assign a16948 = a16944 & ~a16352;
assign a16952 = a16950 & a16480;
assign a16954 = ~a16950 & ~a16480;
assign a16956 = ~a16954 & ~a16952;
assign a16958 = ~a11348 & ~a7998;
assign a16960 = ~a12836 & ~a6916;
assign a16962 = ~a16960 & ~a16958;
assign a16964 = a12836 & a6916;
assign a16966 = ~a16964 & ~a16962;
assign a16968 = ~a12636 & ~a7986;
assign a16970 = ~a16968 & ~a16966;
assign a16972 = a12636 & a7986;
assign a16974 = ~a16972 & ~a16970;
assign a16976 = ~a12436 & ~a7974;
assign a16978 = ~a16976 & ~a16974;
assign a16980 = a12436 & a7974;
assign a16982 = ~a16980 & ~a16978;
assign a16984 = ~a12236 & ~a7962;
assign a16986 = ~a16984 & ~a16982;
assign a16988 = a12236 & a7962;
assign a16990 = ~a16988 & ~a16986;
assign a16992 = ~a12048 & ~a7950;
assign a16994 = ~a16992 & ~a16990;
assign a16996 = a12048 & a7950;
assign a16998 = ~a16996 & ~a16994;
assign a17000 = ~a11788 & ~a7938;
assign a17002 = ~a17000 & ~a16998;
assign a17004 = a11788 & a7938;
assign a17006 = ~a17004 & ~a17002;
assign a17008 = a11246 & a7860;
assign a17010 = ~a11246 & ~a7860;
assign a17012 = ~a17010 & ~a17008;
assign a17014 = ~a17012 & ~a17006;
assign a17016 = a11348 & a7998;
assign a17018 = ~a17016 & ~a16964;
assign a17020 = ~a17018 & ~a16960;
assign a17022 = ~a17020 & ~a16972;
assign a17024 = ~a17022 & ~a16968;
assign a17026 = ~a17024 & ~a16980;
assign a17028 = ~a17026 & ~a16976;
assign a17030 = ~a17028 & ~a16988;
assign a17032 = ~a17030 & ~a16984;
assign a17034 = ~a17032 & ~a16996;
assign a17036 = ~a17034 & ~a16992;
assign a17038 = ~a17036 & ~a17004;
assign a17040 = ~a17038 & ~a17000;
assign a17042 = ~a17040 & a17012;
assign a17044 = ~a17042 & ~a17014;
assign a17046 = ~a17044 & a16956;
assign a17048 = a17046 & a6908;
assign a17050 = a17048 & l576;
assign a17052 = ~a17050 & ~a5572;
assign a17054 = ~a17052 & ~a16802;
assign a17056 = ~a17054 & ~l494;
assign a17058 = a16480 & a6424;
assign a17060 = ~a16480 & ~a6424;
assign a17062 = ~a17060 & ~a17058;
assign a17064 = ~a17062 & a16638;
assign a17066 = a17062 & a16924;
assign a17068 = ~a17066 & ~a17064;
assign a17070 = ~a17068 & a1690;
assign a17074 = a16940 & ~a16340;
assign a17076 = a17074 & a16320;
assign a17078 = ~a17076 & a16496;
assign a17080 = a17076 & ~a16352;
assign a17084 = a17082 & a16492;
assign a17086 = ~a17082 & ~a16492;
assign a17088 = ~a17086 & ~a17084;
assign a17090 = ~a11352 & ~a7998;
assign a17092 = ~a12840 & ~a6916;
assign a17094 = ~a17092 & ~a17090;
assign a17096 = a12840 & a6916;
assign a17098 = ~a17096 & ~a17094;
assign a17100 = ~a12640 & ~a7986;
assign a17102 = ~a17100 & ~a17098;
assign a17104 = a12640 & a7986;
assign a17106 = ~a17104 & ~a17102;
assign a17108 = ~a12440 & ~a7974;
assign a17110 = ~a17108 & ~a17106;
assign a17112 = a12440 & a7974;
assign a17114 = ~a17112 & ~a17110;
assign a17116 = ~a12240 & ~a7962;
assign a17118 = ~a17116 & ~a17114;
assign a17120 = a12240 & a7962;
assign a17122 = ~a17120 & ~a17118;
assign a17124 = ~a12052 & ~a7950;
assign a17126 = ~a17124 & ~a17122;
assign a17128 = a12052 & a7950;
assign a17130 = ~a17128 & ~a17126;
assign a17132 = ~a11792 & ~a7938;
assign a17134 = ~a17132 & ~a17130;
assign a17136 = a11792 & a7938;
assign a17138 = ~a17136 & ~a17134;
assign a17140 = a11250 & a7860;
assign a17142 = ~a11250 & ~a7860;
assign a17144 = ~a17142 & ~a17140;
assign a17146 = ~a17144 & ~a17138;
assign a17148 = a11352 & a7998;
assign a17150 = ~a17148 & ~a17096;
assign a17152 = ~a17150 & ~a17092;
assign a17154 = ~a17152 & ~a17104;
assign a17156 = ~a17154 & ~a17100;
assign a17158 = ~a17156 & ~a17112;
assign a17160 = ~a17158 & ~a17108;
assign a17162 = ~a17160 & ~a17120;
assign a17164 = ~a17162 & ~a17116;
assign a17166 = ~a17164 & ~a17128;
assign a17168 = ~a17166 & ~a17124;
assign a17170 = ~a17168 & ~a17136;
assign a17172 = ~a17170 & ~a17132;
assign a17174 = ~a17172 & a17144;
assign a17176 = ~a17174 & ~a17146;
assign a17178 = ~a17176 & a17088;
assign a17180 = a17178 & a6908;
assign a17182 = a17180 & l578;
assign a17184 = ~a17182 & l576;
assign a17186 = ~a17184 & ~a16944;
assign a17188 = ~a17186 & ~l494;
assign a17190 = a16492 & a6424;
assign a17192 = ~a16492 & ~a6424;
assign a17194 = ~a17192 & ~a17190;
assign a17196 = ~a17194 & a16638;
assign a17198 = ~a16648 & ~a6592;
assign a17200 = ~a17198 & a6476;
assign a17202 = a17200 & a17194;
assign a17204 = ~a17202 & ~a17196;
assign a17206 = ~a17204 & a1690;
assign a17210 = a16942 & ~a16320;
assign a17212 = ~a17210 & a16504;
assign a17214 = a17210 & ~a16352;
assign a17218 = a17216 & a16496;
assign a17220 = ~a17216 & ~a16496;
assign a17222 = ~a17220 & ~a17218;
assign a17224 = ~a11360 & ~a7998;
assign a17226 = ~a12848 & ~a6916;
assign a17228 = ~a17226 & ~a17224;
assign a17230 = a12848 & a6916;
assign a17232 = ~a17230 & ~a17228;
assign a17234 = ~a12648 & ~a7986;
assign a17236 = ~a17234 & ~a17232;
assign a17238 = a12648 & a7986;
assign a17240 = ~a17238 & ~a17236;
assign a17242 = ~a12448 & ~a7974;
assign a17244 = ~a17242 & ~a17240;
assign a17246 = a12448 & a7974;
assign a17248 = ~a17246 & ~a17244;
assign a17250 = ~a12248 & ~a7962;
assign a17252 = ~a17250 & ~a17248;
assign a17254 = a12248 & a7962;
assign a17256 = ~a17254 & ~a17252;
assign a17258 = ~a12060 & ~a7950;
assign a17260 = ~a17258 & ~a17256;
assign a17262 = a12060 & a7950;
assign a17264 = ~a17262 & ~a17260;
assign a17266 = ~a11800 & ~a7938;
assign a17268 = ~a17266 & ~a17264;
assign a17270 = a11800 & a7938;
assign a17272 = ~a17270 & ~a17268;
assign a17274 = a11258 & a7860;
assign a17276 = ~a11258 & ~a7860;
assign a17278 = ~a17276 & ~a17274;
assign a17280 = ~a17278 & ~a17272;
assign a17282 = a11360 & a7998;
assign a17284 = ~a17282 & ~a17230;
assign a17286 = ~a17284 & ~a17226;
assign a17288 = ~a17286 & ~a17238;
assign a17290 = ~a17288 & ~a17234;
assign a17292 = ~a17290 & ~a17246;
assign a17294 = ~a17292 & ~a17242;
assign a17296 = ~a17294 & ~a17254;
assign a17298 = ~a17296 & ~a17250;
assign a17300 = ~a17298 & ~a17262;
assign a17302 = ~a17300 & ~a17258;
assign a17304 = ~a17302 & ~a17270;
assign a17306 = ~a17304 & ~a17266;
assign a17308 = ~a17306 & a17278;
assign a17310 = ~a17308 & ~a17280;
assign a17312 = ~a17310 & a17222;
assign a17314 = a17312 & a6908;
assign a17316 = a17314 & l580;
assign a17318 = ~a17316 & l578;
assign a17320 = ~a17318 & ~a17076;
assign a17322 = ~a17320 & ~l494;
assign a17324 = a16496 & a6424;
assign a17326 = ~a16496 & ~a6424;
assign a17328 = ~a17326 & ~a17324;
assign a17330 = ~a17328 & a16638;
assign a17332 = ~a6592 & ~a6548;
assign a17334 = ~a17332 & a6476;
assign a17336 = a17334 & a17328;
assign a17338 = ~a17336 & ~a17330;
assign a17340 = ~a17338 & a1690;
assign a17344 = a17074 & ~a16320;
assign a17346 = ~a17344 & a16508;
assign a17348 = a17344 & ~a16352;
assign a17352 = a17350 & a16504;
assign a17354 = ~a17350 & ~a16504;
assign a17356 = ~a17354 & ~a17352;
assign a17358 = ~a11364 & ~a7998;
assign a17360 = ~a12852 & ~a6916;
assign a17362 = ~a17360 & ~a17358;
assign a17364 = a12852 & a6916;
assign a17366 = ~a17364 & ~a17362;
assign a17368 = ~a12652 & ~a7986;
assign a17370 = ~a17368 & ~a17366;
assign a17372 = a12652 & a7986;
assign a17374 = ~a17372 & ~a17370;
assign a17376 = ~a12452 & ~a7974;
assign a17378 = ~a17376 & ~a17374;
assign a17380 = a12452 & a7974;
assign a17382 = ~a17380 & ~a17378;
assign a17384 = ~a12252 & ~a7962;
assign a17386 = ~a17384 & ~a17382;
assign a17388 = a12252 & a7962;
assign a17390 = ~a17388 & ~a17386;
assign a17392 = ~a12064 & ~a7950;
assign a17394 = ~a17392 & ~a17390;
assign a17396 = a12064 & a7950;
assign a17398 = ~a17396 & ~a17394;
assign a17400 = ~a11804 & ~a7938;
assign a17402 = ~a17400 & ~a17398;
assign a17404 = a11804 & a7938;
assign a17406 = ~a17404 & ~a17402;
assign a17408 = a11262 & a7860;
assign a17410 = ~a11262 & ~a7860;
assign a17412 = ~a17410 & ~a17408;
assign a17414 = ~a17412 & ~a17406;
assign a17416 = a11364 & a7998;
assign a17418 = ~a17416 & ~a17364;
assign a17420 = ~a17418 & ~a17360;
assign a17422 = ~a17420 & ~a17372;
assign a17424 = ~a17422 & ~a17368;
assign a17426 = ~a17424 & ~a17380;
assign a17428 = ~a17426 & ~a17376;
assign a17430 = ~a17428 & ~a17388;
assign a17432 = ~a17430 & ~a17384;
assign a17434 = ~a17432 & ~a17396;
assign a17436 = ~a17434 & ~a17392;
assign a17438 = ~a17436 & ~a17404;
assign a17440 = ~a17438 & ~a17400;
assign a17442 = ~a17440 & a17412;
assign a17444 = ~a17442 & ~a17414;
assign a17446 = ~a17444 & a17356;
assign a17448 = a17446 & a6908;
assign a17450 = a17448 & l582;
assign a17452 = ~a17450 & l580;
assign a17454 = ~a17452 & ~a17210;
assign a17456 = ~a17454 & ~l494;
assign a17458 = a16504 & a6424;
assign a17460 = ~a16504 & ~a6424;
assign a17462 = ~a17460 & ~a17458;
assign a17464 = ~a17462 & a16638;
assign a17466 = a17332 & ~a6512;
assign a17468 = ~a17466 & a6476;
assign a17470 = a17468 & a17462;
assign a17472 = ~a17470 & ~a17464;
assign a17474 = ~a17472 & a1690;
assign a17478 = ~a16334 & a6934;
assign a17480 = a17478 & a16328;
assign a17482 = a17480 & a16340;
assign a17484 = ~a17482 & a16524;
assign a17486 = a17482 & ~a16352;
assign a17490 = a17488 & a16508;
assign a17492 = ~a17488 & ~a16508;
assign a17494 = ~a17492 & ~a17490;
assign a17496 = ~a11292 & ~a7998;
assign a17498 = ~a12868 & ~a6916;
assign a17500 = ~a17498 & ~a17496;
assign a17502 = a12868 & a6916;
assign a17504 = ~a17502 & ~a17500;
assign a17506 = ~a12668 & ~a7986;
assign a17508 = ~a17506 & ~a17504;
assign a17510 = a12668 & a7986;
assign a17512 = ~a17510 & ~a17508;
assign a17514 = ~a12468 & ~a7974;
assign a17516 = ~a17514 & ~a17512;
assign a17518 = a12468 & a7974;
assign a17520 = ~a17518 & ~a17516;
assign a17522 = ~a12268 & ~a7962;
assign a17524 = ~a17522 & ~a17520;
assign a17526 = a12268 & a7962;
assign a17528 = ~a17526 & ~a17524;
assign a17530 = ~a12080 & ~a7950;
assign a17532 = ~a17530 & ~a17528;
assign a17534 = a12080 & a7950;
assign a17536 = ~a17534 & ~a17532;
assign a17538 = ~a11820 & ~a7938;
assign a17540 = ~a17538 & ~a17536;
assign a17542 = a11820 & a7938;
assign a17544 = ~a17542 & ~a17540;
assign a17546 = a11202 & a7860;
assign a17548 = ~a11202 & ~a7860;
assign a17550 = ~a17548 & ~a17546;
assign a17552 = ~a17550 & ~a17544;
assign a17554 = a11292 & a7998;
assign a17556 = ~a17554 & ~a17502;
assign a17558 = ~a17556 & ~a17498;
assign a17560 = ~a17558 & ~a17510;
assign a17562 = ~a17560 & ~a17506;
assign a17564 = ~a17562 & ~a17518;
assign a17566 = ~a17564 & ~a17514;
assign a17568 = ~a17566 & ~a17526;
assign a17570 = ~a17568 & ~a17522;
assign a17572 = ~a17570 & ~a17534;
assign a17574 = ~a17572 & ~a17530;
assign a17576 = ~a17574 & ~a17542;
assign a17578 = ~a17576 & ~a17538;
assign a17580 = ~a17578 & a17550;
assign a17582 = ~a17580 & ~a17552;
assign a17584 = ~a17582 & a17494;
assign a17586 = a17584 & a6908;
assign a17588 = a17586 & l586;
assign a17590 = ~a17588 & l582;
assign a17592 = ~a17590 & ~a17344;
assign a17594 = ~a17592 & ~l494;
assign a17596 = a16508 & a6424;
assign a17598 = ~a16508 & ~a6424;
assign a17600 = ~a17598 & ~a17596;
assign a17602 = ~a17600 & a16638;
assign a17604 = a17600 & a6476;
assign a17606 = ~a17604 & ~a17602;
assign a17608 = ~a17606 & a1690;
assign a17612 = ~a16462 & a16312;
assign a17614 = a16462 & ~a16352;
assign a17618 = a17616 & a16528;
assign a17620 = ~a17616 & ~a16528;
assign a17622 = ~a17620 & ~a17618;
assign a17624 = ~a11304 & ~a7998;
assign a17626 = ~a12796 & ~a6916;
assign a17628 = ~a17626 & ~a17624;
assign a17630 = a12796 & a6916;
assign a17632 = ~a17630 & ~a17628;
assign a17634 = ~a12596 & ~a7986;
assign a17636 = ~a17634 & ~a17632;
assign a17638 = a12596 & a7986;
assign a17640 = ~a17638 & ~a17636;
assign a17642 = ~a12396 & ~a7974;
assign a17644 = ~a17642 & ~a17640;
assign a17646 = a12396 & a7974;
assign a17648 = ~a17646 & ~a17644;
assign a17650 = ~a12196 & ~a7962;
assign a17652 = ~a17650 & ~a17648;
assign a17654 = a12196 & a7962;
assign a17656 = ~a17654 & ~a17652;
assign a17658 = ~a12008 & ~a7950;
assign a17660 = ~a17658 & ~a17656;
assign a17662 = a12008 & a7950;
assign a17664 = ~a17662 & ~a17660;
assign a17666 = ~a11752 & ~a7938;
assign a17668 = ~a17666 & ~a17664;
assign a17670 = a11752 & a7938;
assign a17672 = ~a17670 & ~a17668;
assign a17674 = a11214 & a7860;
assign a17676 = ~a11214 & ~a7860;
assign a17678 = ~a17676 & ~a17674;
assign a17680 = ~a17678 & ~a17672;
assign a17682 = a11304 & a7998;
assign a17684 = ~a17682 & ~a17630;
assign a17686 = ~a17684 & ~a17626;
assign a17688 = ~a17686 & ~a17638;
assign a17690 = ~a17688 & ~a17634;
assign a17692 = ~a17690 & ~a17646;
assign a17694 = ~a17692 & ~a17642;
assign a17696 = ~a17694 & ~a17654;
assign a17698 = ~a17696 & ~a17650;
assign a17700 = ~a17698 & ~a17662;
assign a17702 = ~a17700 & ~a17658;
assign a17704 = ~a17702 & ~a17670;
assign a17706 = ~a17704 & ~a17666;
assign a17708 = ~a17706 & a17678;
assign a17710 = ~a17708 & ~a17680;
assign a17712 = ~a17710 & ~a17622;
assign a17714 = a17712 & a6908;
assign a17716 = a17714 & ~a5542;
assign a17718 = ~a17716 & l584;
assign a17720 = a17480 & ~a16340;
assign a17722 = ~a17720 & ~a17718;
assign a17724 = ~a17722 & ~l494;
assign a17726 = a16528 & a6424;
assign a17728 = ~a16528 & ~a6424;
assign a17730 = ~a17728 & ~a17726;
assign a17732 = ~a17730 & a16638;
assign a17734 = ~a16790 & ~a6476;
assign a17736 = ~a17734 & a17730;
assign a17738 = ~a17736 & ~a17732;
assign a17740 = ~a17738 & a1690;
assign a17744 = ~a17720 & a16528;
assign a17746 = a17720 & ~a16352;
assign a17750 = a17748 & a16524;
assign a17752 = ~a17748 & ~a16524;
assign a17754 = ~a17752 & ~a17750;
assign a17756 = ~a11296 & ~a7998;
assign a17758 = ~a12872 & ~a6916;
assign a17760 = ~a17758 & ~a17756;
assign a17762 = a12872 & a6916;
assign a17764 = ~a17762 & ~a17760;
assign a17766 = ~a12672 & ~a7986;
assign a17768 = ~a17766 & ~a17764;
assign a17770 = a12672 & a7986;
assign a17772 = ~a17770 & ~a17768;
assign a17774 = ~a12472 & ~a7974;
assign a17776 = ~a17774 & ~a17772;
assign a17778 = a12472 & a7974;
assign a17780 = ~a17778 & ~a17776;
assign a17782 = ~a12272 & ~a7962;
assign a17784 = ~a17782 & ~a17780;
assign a17786 = a12272 & a7962;
assign a17788 = ~a17786 & ~a17784;
assign a17790 = ~a12084 & ~a7950;
assign a17792 = ~a17790 & ~a17788;
assign a17794 = a12084 & a7950;
assign a17796 = ~a17794 & ~a17792;
assign a17798 = ~a11824 & ~a7938;
assign a17800 = ~a17798 & ~a17796;
assign a17802 = a11824 & a7938;
assign a17804 = ~a17802 & ~a17800;
assign a17806 = a11206 & a7860;
assign a17808 = ~a11206 & ~a7860;
assign a17810 = ~a17808 & ~a17806;
assign a17812 = ~a17810 & ~a17804;
assign a17814 = a11296 & a7998;
assign a17816 = ~a17814 & ~a17762;
assign a17818 = ~a17816 & ~a17758;
assign a17820 = ~a17818 & ~a17770;
assign a17822 = ~a17820 & ~a17766;
assign a17824 = ~a17822 & ~a17778;
assign a17826 = ~a17824 & ~a17774;
assign a17828 = ~a17826 & ~a17786;
assign a17830 = ~a17828 & ~a17782;
assign a17832 = ~a17830 & ~a17794;
assign a17834 = ~a17832 & ~a17790;
assign a17836 = ~a17834 & ~a17802;
assign a17838 = ~a17836 & ~a17798;
assign a17840 = ~a17838 & a17810;
assign a17842 = ~a17840 & ~a17812;
assign a17844 = ~a17842 & a17754;
assign a17846 = a17844 & l584;
assign a17848 = a17846 & a6908;
assign a17850 = ~a17848 & l586;
assign a17852 = ~a17850 & ~a17482;
assign a17854 = ~a17852 & ~l494;
assign a17856 = a16524 & a6424;
assign a17858 = ~a16524 & ~a6424;
assign a17860 = ~a17858 & ~a17856;
assign a17862 = ~a17860 & a16638;
assign a17864 = ~a16650 & ~a6476;
assign a17866 = ~a17864 & a17860;
assign a17868 = ~a17866 & ~a17862;
assign a17870 = ~a17868 & a1690;
assign a17874 = ~a5124 & l664;
assign a17876 = a6646 & ~a2270;
assign a17878 = ~a17876 & ~a17874;
assign a17880 = a6642 & a2270;
assign a17884 = a6642 & a2280;
assign a17886 = a2280 & l604;
assign a17888 = ~a2296 & ~a2280;
assign a17890 = a17888 & a2270;
assign a17892 = ~a17890 & ~a17886;
assign a17894 = ~a17892 & a6646;
assign a17896 = ~a17894 & ~a17884;
assign a17898 = ~a6562 & l664;
assign a17902 = a6642 & a2302;
assign a17904 = ~a6650 & a2302;
assign a17906 = a6650 & ~a2302;
assign a17908 = ~a17906 & ~a17904;
assign a17910 = ~a17908 & a6646;
assign a17912 = ~a17910 & ~a17902;
assign a17914 = ~a6604 & l664;
assign a17918 = l1686 & ~l1674;
assign a17920 = l1686 & ~l1670;
assign a17922 = l1686 & ~l1666;
assign a17924 = l1686 & ~l1662;
assign a17926 = l1686 & ~l680;
assign a17928 = a6696 & ~a6690;
assign a17930 = a17928 & a6702;
assign a17932 = a17930 & a17926;
assign a17934 = l1686 & ~l668;
assign a17936 = ~a6708 & a6702;
assign a17938 = a17936 & a6690;
assign a17940 = a17938 & a17934;
assign a17942 = ~a17940 & ~a17932;
assign a17944 = l1686 & ~l670;
assign a17946 = ~a6696 & ~a6690;
assign a17948 = a17946 & a6708;
assign a17950 = a17948 & ~a6702;
assign a17952 = a17950 & a17944;
assign a17954 = ~a17952 & a17942;
assign a17956 = l1686 & ~l684;
assign a17958 = a17956 & a6702;
assign a17960 = a17958 & a17948;
assign a17962 = l1686 & ~l672;
assign a17964 = a6708 & a6696;
assign a17966 = a17964 & a6690;
assign a17968 = a17966 & a6702;
assign a17970 = a17968 & a17962;
assign a17972 = ~a17970 & ~a17960;
assign a17974 = a17972 & a17954;
assign a17976 = l1686 & ~l686;
assign a17978 = ~a6702 & ~a6696;
assign a17980 = a17978 & a6690;
assign a17982 = a17980 & a17976;
assign a17984 = a17982 & a6708;
assign a17986 = l1686 & ~l678;
assign a17988 = a17986 & ~a6702;
assign a17990 = a17988 & a17928;
assign a17992 = l1686 & ~l674;
assign a17994 = ~a6708 & ~a6702;
assign a17996 = a17994 & a6690;
assign a17998 = a17996 & a17992;
assign a18000 = ~a17998 & ~a17990;
assign a18002 = a18000 & ~a17984;
assign a18004 = l1686 & ~l682;
assign a18006 = ~a6702 & a6696;
assign a18008 = a18006 & a6708;
assign a18010 = a18008 & a18004;
assign a18012 = l1686 & ~l676;
assign a18014 = a6702 & ~a6696;
assign a18016 = a18014 & a6708;
assign a18018 = a18016 & a18012;
assign a18020 = ~a18018 & ~a18010;
assign a18022 = ~a18020 & a6690;
assign a18024 = ~a18022 & a18002;
assign a18028 = l1686 & ~l1600;
assign a18030 = a6642 & a1688;
assign a18032 = ~a6444 & l664;
assign a18034 = ~a18032 & ~a18030;
assign a18036 = a17886 & ~a2302;
assign a18038 = a18036 & a17976;
assign a18040 = a2302 & l610;
assign a18042 = a18040 & a2270;
assign a18044 = a18042 & a17956;
assign a18046 = ~a18044 & ~a18038;
assign a18048 = a17888 & ~a2270;
assign a18050 = a18048 & ~a2302;
assign a18052 = a18050 & a18004;
assign a18054 = ~a18052 & a18046;
assign a18056 = a17926 & a17906;
assign a18058 = a18040 & ~a2270;
assign a18060 = a18058 & a17986;
assign a18062 = ~a18060 & ~a18056;
assign a18064 = a17890 & ~a2302;
assign a18066 = a18064 & a18012;
assign a18068 = ~a18066 & a18062;
assign a18070 = a18068 & a18054;
assign a18072 = a17992 & a6648;
assign a18074 = a2296 & a2270;
assign a18076 = a18074 & ~a2302;
assign a18078 = a18076 & a17962;
assign a18080 = ~a18078 & ~a18072;
assign a18082 = a2370 & ~a2270;
assign a18084 = a18082 & a17944;
assign a18086 = ~a18084 & a18080;
assign a18088 = a6652 & ~a2296;
assign a18090 = a18088 & a17934;
assign a18092 = ~a18090 & a18086;
assign a18094 = a18092 & a18070;
assign a18096 = ~a18094 & a6646;
assign a18100 = a1704 & ~l1686;
assign a18102 = l1686 & l908;
assign a18104 = ~a18102 & ~a18100;
assign a18106 = ~a18104 & a18076;
assign a18108 = a17906 & l910;
assign a18110 = ~a18108 & ~a18106;
assign a18112 = a18088 & l906;
assign a18114 = ~a18112 & a18110;
assign a18116 = a18042 & l902;
assign a18118 = a18058 & l912;
assign a18120 = ~a18118 & ~a18116;
assign a18122 = a8084 & ~l1686;
assign a18124 = l1686 & l900;
assign a18126 = ~a18124 & ~a18122;
assign a18128 = ~a18126 & a18050;
assign a18130 = ~a18128 & a18120;
assign a18132 = a18130 & a18114;
assign a18134 = l1686 & l918;
assign a18136 = ~a18134 & ~a8064;
assign a18138 = ~a18136 & a6648;
assign a18140 = a18036 & l916;
assign a18142 = ~a18140 & ~a18138;
assign a18144 = l914 & ~l664;
assign a18146 = a18144 & a18082;
assign a18148 = ~a18146 & a18142;
assign a18150 = a18064 & l904;
assign a18152 = ~a18150 & a18148;
assign a18154 = a18152 & a18132;
assign a18156 = ~a18154 & l666;
assign a18158 = ~a18136 & a18076;
assign a18160 = a17906 & l916;
assign a18162 = ~a18160 & ~a18158;
assign a18164 = a18144 & a18088;
assign a18166 = ~a18164 & a18162;
assign a18168 = a18042 & l912;
assign a18170 = a18058 & l910;
assign a18172 = ~a18170 & ~a18168;
assign a18174 = ~a18104 & a18050;
assign a18176 = ~a18174 & a18172;
assign a18178 = a18176 & a18166;
assign a18180 = a6648 & l906;
assign a18182 = a18036 & l904;
assign a18184 = ~a18182 & ~a18180;
assign a18186 = a18082 & l902;
assign a18188 = ~a18186 & a18184;
assign a18190 = ~a18126 & a18064;
assign a18192 = ~a18190 & a18188;
assign a18194 = a18192 & a18178;
assign a18196 = ~a18194 & ~l666;
assign a18198 = ~a18196 & ~a18156;
assign a18200 = l1686 & ~l888;
assign a18202 = a18200 & a18088;
assign a18204 = l1686 & ~l892;
assign a18206 = a18204 & a2370;
assign a18208 = a18206 & ~a2270;
assign a18210 = ~a18208 & ~a18202;
assign a18212 = l1686 & ~l880;
assign a18214 = a18212 & l612;
assign a18216 = a18214 & a18074;
assign a18218 = l1686 & ~l898;
assign a18220 = a18218 & a6648;
assign a18222 = ~a18220 & ~a18216;
assign a18224 = l1686 & ~l896;
assign a18226 = a18224 & a18040;
assign a18228 = a18226 & ~a2270;
assign a18230 = ~a18228 & a18222;
assign a18232 = l1686 & ~l894;
assign a18234 = a18232 & a18042;
assign a18236 = l1686 & ~l884;
assign a18238 = a18236 & a17906;
assign a18240 = ~a18238 & ~a18234;
assign a18242 = a18240 & a18230;
assign a18244 = a18242 & a18210;
assign a18246 = l1686 & ~l890;
assign a18248 = a18246 & a2338;
assign a18250 = a18248 & ~a2270;
assign a18252 = l1686 & ~l882;
assign a18254 = a18252 & a18036;
assign a18256 = l1686 & ~l886;
assign a18258 = a18256 & l612;
assign a18260 = a18258 & a17890;
assign a18262 = ~a18260 & ~a18254;
assign a18264 = a18262 & ~a18250;
assign a18266 = a18264 & a18244;
assign a18268 = ~a18266 & l666;
assign a18270 = a18218 & a18076;
assign a18272 = a18226 & a2270;
assign a18274 = ~a18272 & ~a18270;
assign a18276 = a18232 & a18082;
assign a18278 = ~a18276 & a18274;
assign a18280 = ~a18248 & ~a18206;
assign a18282 = ~a18280 & a2270;
assign a18284 = ~a18282 & a18278;
assign a18286 = a18200 & a6648;
assign a18288 = a18258 & a17886;
assign a18290 = ~a18288 & ~a18286;
assign a18292 = a18236 & a18058;
assign a18294 = ~a18292 & a18290;
assign a18296 = a18252 & a17906;
assign a18298 = a18214 & a18048;
assign a18300 = ~a18298 & ~a18296;
assign a18302 = a18300 & a18294;
assign a18304 = a18302 & a18284;
assign a18306 = ~a18304 & ~l666;
assign a18308 = ~a18306 & ~a18268;
assign a18310 = ~a18308 & a8042;
assign a18312 = a18308 & ~a8042;
assign a18314 = ~a18312 & ~a18310;
assign a18316 = l1686 & ~l734;
assign a18318 = a18316 & a18088;
assign a18320 = l1686 & ~l738;
assign a18322 = a18320 & a2370;
assign a18324 = a18322 & ~a2270;
assign a18326 = ~a18324 & ~a18318;
assign a18328 = l1686 & ~l726;
assign a18330 = a18328 & l612;
assign a18332 = a18330 & a18074;
assign a18334 = l1686 & ~l744;
assign a18336 = a18334 & a6648;
assign a18338 = ~a18336 & ~a18332;
assign a18340 = l1686 & ~l742;
assign a18342 = a18340 & a18040;
assign a18344 = a18342 & ~a2270;
assign a18346 = ~a18344 & a18338;
assign a18348 = l1686 & ~l740;
assign a18350 = a18348 & a18042;
assign a18352 = l1686 & ~l730;
assign a18354 = a18352 & a17906;
assign a18356 = ~a18354 & ~a18350;
assign a18358 = a18356 & a18346;
assign a18360 = a18358 & a18326;
assign a18362 = ~a8506 & ~l1686;
assign a18364 = l1686 & l736;
assign a18366 = ~a18364 & ~a18362;
assign a18368 = a18366 & a2338;
assign a18370 = a18368 & ~a2270;
assign a18372 = l1686 & ~l728;
assign a18374 = a18372 & a18036;
assign a18376 = l1686 & ~l732;
assign a18378 = a18376 & l612;
assign a18380 = a18378 & a17890;
assign a18382 = ~a18380 & ~a18374;
assign a18384 = a18382 & ~a18370;
assign a18386 = a18384 & a18360;
assign a18388 = ~a18386 & l666;
assign a18390 = a18334 & a18076;
assign a18392 = a18342 & a2270;
assign a18394 = ~a18392 & ~a18390;
assign a18396 = a18348 & a18082;
assign a18398 = ~a18396 & a18394;
assign a18400 = ~a18368 & ~a18322;
assign a18402 = ~a18400 & a2270;
assign a18404 = ~a18402 & a18398;
assign a18406 = a18316 & a6648;
assign a18408 = a18378 & a17886;
assign a18410 = ~a18408 & ~a18406;
assign a18412 = a18352 & a18058;
assign a18414 = ~a18412 & a18410;
assign a18416 = a18372 & a17906;
assign a18418 = a18330 & a18048;
assign a18420 = ~a18418 & ~a18416;
assign a18422 = a18420 & a18414;
assign a18424 = a18422 & a18404;
assign a18426 = ~a18424 & ~l666;
assign a18428 = ~a18426 & ~a18388;
assign a18430 = a18428 & ~a16052;
assign a18432 = ~a18430 & a18314;
assign a18434 = l1686 & ~l866;
assign a18436 = a18434 & a18088;
assign a18438 = l1686 & ~l870;
assign a18440 = a18438 & a2370;
assign a18442 = a18440 & ~a2270;
assign a18444 = ~a18442 & ~a18436;
assign a18446 = l1686 & l858;
assign a18448 = ~a18446 & ~a10154;
assign a18450 = a18448 & ~a2302;
assign a18452 = a18450 & a18074;
assign a18454 = l1686 & ~l876;
assign a18456 = a18454 & a6648;
assign a18458 = ~a18456 & ~a18452;
assign a18460 = l1686 & ~l874;
assign a18462 = a18460 & a18040;
assign a18464 = a18462 & ~a2270;
assign a18466 = ~a18464 & a18458;
assign a18468 = l1686 & ~l872;
assign a18470 = a18468 & a18042;
assign a18472 = l1686 & ~l862;
assign a18474 = a18472 & a17906;
assign a18476 = ~a18474 & ~a18470;
assign a18478 = a18476 & a18466;
assign a18480 = a18478 & a18444;
assign a18482 = ~a8094 & ~l1686;
assign a18484 = l1686 & l868;
assign a18486 = ~a18484 & ~a18482;
assign a18488 = a18486 & a2338;
assign a18490 = a18488 & ~a2270;
assign a18492 = l1686 & ~l860;
assign a18494 = a18492 & a18036;
assign a18496 = l1686 & ~l864;
assign a18498 = a18496 & l612;
assign a18500 = a18498 & a17890;
assign a18502 = ~a18500 & ~a18494;
assign a18504 = a18502 & ~a18490;
assign a18506 = a18504 & a18480;
assign a18508 = ~a18506 & l666;
assign a18510 = a18454 & a18076;
assign a18512 = a18462 & a2270;
assign a18514 = ~a18512 & ~a18510;
assign a18516 = a18468 & a18082;
assign a18518 = ~a18516 & a18514;
assign a18520 = ~a18488 & ~a18440;
assign a18522 = ~a18520 & a2270;
assign a18524 = ~a18522 & a18518;
assign a18526 = a18434 & a6648;
assign a18528 = a18498 & a17886;
assign a18530 = ~a18528 & ~a18526;
assign a18532 = a18472 & a18058;
assign a18534 = ~a18532 & a18530;
assign a18536 = a18492 & a17906;
assign a18538 = a18450 & a18048;
assign a18540 = ~a18538 & ~a18536;
assign a18542 = a18540 & a18534;
assign a18544 = a18542 & a18524;
assign a18546 = ~a18544 & ~l666;
assign a18548 = ~a18546 & ~a18508;
assign a18550 = ~a18548 & a16120;
assign a18552 = l1686 & ~l844;
assign a18554 = a18552 & a18088;
assign a18556 = l1686 & ~l848;
assign a18558 = a18556 & a2370;
assign a18560 = a18558 & ~a2270;
assign a18562 = ~a18560 & ~a18554;
assign a18564 = l1686 & l836;
assign a18566 = ~a18564 & ~a10200;
assign a18568 = a18566 & ~a2302;
assign a18570 = a18568 & a18074;
assign a18572 = l1686 & ~l854;
assign a18574 = a18572 & a6648;
assign a18576 = ~a18574 & ~a18570;
assign a18578 = l1686 & ~l852;
assign a18580 = a18578 & a18040;
assign a18582 = a18580 & ~a2270;
assign a18584 = ~a18582 & a18576;
assign a18586 = l1686 & ~l850;
assign a18588 = a18586 & a18042;
assign a18590 = l1686 & ~l840;
assign a18592 = a18590 & a17906;
assign a18594 = ~a18592 & ~a18588;
assign a18596 = a18594 & a18584;
assign a18598 = a18596 & a18562;
assign a18600 = ~a8108 & ~l1686;
assign a18602 = l1686 & l846;
assign a18604 = ~a18602 & ~a18600;
assign a18606 = a18604 & a2338;
assign a18608 = a18606 & ~a2270;
assign a18610 = l1686 & ~l838;
assign a18612 = a18610 & a18036;
assign a18614 = l1686 & ~l842;
assign a18616 = a18614 & l612;
assign a18618 = a18616 & a17890;
assign a18620 = ~a18618 & ~a18612;
assign a18622 = a18620 & ~a18608;
assign a18624 = a18622 & a18598;
assign a18626 = ~a18624 & l666;
assign a18628 = a18572 & a18076;
assign a18630 = a18580 & a2270;
assign a18632 = ~a18630 & ~a18628;
assign a18634 = a18586 & a18082;
assign a18636 = ~a18634 & a18632;
assign a18638 = ~a18606 & ~a18558;
assign a18640 = ~a18638 & a2270;
assign a18642 = ~a18640 & a18636;
assign a18644 = a18552 & a6648;
assign a18646 = a18616 & a17886;
assign a18648 = ~a18646 & ~a18644;
assign a18650 = a18590 & a18058;
assign a18652 = ~a18650 & a18648;
assign a18654 = a18610 & a17906;
assign a18656 = a18568 & a18048;
assign a18658 = ~a18656 & ~a18654;
assign a18660 = a18658 & a18652;
assign a18662 = a18660 & a18642;
assign a18664 = ~a18662 & ~l666;
assign a18666 = ~a18664 & ~a18626;
assign a18668 = ~a18666 & a16110;
assign a18670 = ~a18668 & ~a18550;
assign a18672 = a18666 & ~a16110;
assign a18674 = ~a18672 & ~a18670;
assign a18676 = l1686 & ~l822;
assign a18678 = a18676 & a18088;
assign a18680 = l1686 & ~l826;
assign a18682 = a18680 & a2370;
assign a18684 = a18682 & ~a2270;
assign a18686 = ~a18684 & ~a18678;
assign a18688 = l1686 & l814;
assign a18690 = ~a18688 & ~a10250;
assign a18692 = a18690 & ~a2302;
assign a18694 = a18692 & a18074;
assign a18696 = l1686 & ~l832;
assign a18698 = a18696 & a6648;
assign a18700 = ~a18698 & ~a18694;
assign a18702 = l1686 & ~l830;
assign a18704 = a18702 & a18040;
assign a18706 = a18704 & ~a2270;
assign a18708 = ~a18706 & a18700;
assign a18710 = l1686 & ~l828;
assign a18712 = a18710 & a18042;
assign a18714 = l1686 & ~l818;
assign a18716 = a18714 & a17906;
assign a18718 = ~a18716 & ~a18712;
assign a18720 = a18718 & a18708;
assign a18722 = a18720 & a18686;
assign a18724 = ~a8128 & ~l1686;
assign a18726 = l1686 & l824;
assign a18728 = ~a18726 & ~a18724;
assign a18730 = a18728 & a2338;
assign a18732 = a18730 & ~a2270;
assign a18734 = l1686 & ~l816;
assign a18736 = a18734 & a18036;
assign a18738 = l1686 & ~l820;
assign a18740 = a18738 & l612;
assign a18742 = a18740 & a17890;
assign a18744 = ~a18742 & ~a18736;
assign a18746 = a18744 & ~a18732;
assign a18748 = a18746 & a18722;
assign a18750 = ~a18748 & l666;
assign a18752 = a18696 & a18076;
assign a18754 = a18704 & a2270;
assign a18756 = ~a18754 & ~a18752;
assign a18758 = a18710 & a18082;
assign a18760 = ~a18758 & a18756;
assign a18762 = ~a18730 & ~a18682;
assign a18764 = ~a18762 & a2270;
assign a18766 = ~a18764 & a18760;
assign a18768 = a18676 & a6648;
assign a18770 = a18740 & a17886;
assign a18772 = ~a18770 & ~a18768;
assign a18774 = a18714 & a18058;
assign a18776 = ~a18774 & a18772;
assign a18778 = a18734 & a17906;
assign a18780 = a18692 & a18048;
assign a18782 = ~a18780 & ~a18778;
assign a18784 = a18782 & a18776;
assign a18786 = a18784 & a18766;
assign a18788 = ~a18786 & ~l666;
assign a18790 = ~a18788 & ~a18750;
assign a18792 = ~a18790 & a16100;
assign a18794 = ~a18792 & ~a18674;
assign a18796 = a18790 & ~a16100;
assign a18798 = ~a18796 & ~a18794;
assign a18800 = l1686 & ~l800;
assign a18802 = a18800 & a18088;
assign a18804 = l1686 & ~l804;
assign a18806 = a18804 & a2370;
assign a18808 = a18806 & ~a2270;
assign a18810 = ~a18808 & ~a18802;
assign a18812 = l1686 & l792;
assign a18814 = ~a18812 & ~a10312;
assign a18816 = a18814 & ~a2302;
assign a18818 = a18816 & a18074;
assign a18820 = l1686 & ~l810;
assign a18822 = a18820 & a6648;
assign a18824 = ~a18822 & ~a18818;
assign a18826 = l1686 & ~l808;
assign a18828 = a18826 & a18040;
assign a18830 = a18828 & ~a2270;
assign a18832 = ~a18830 & a18824;
assign a18834 = l1686 & ~l806;
assign a18836 = a18834 & a18042;
assign a18838 = l1686 & ~l796;
assign a18840 = a18838 & a17906;
assign a18842 = ~a18840 & ~a18836;
assign a18844 = a18842 & a18832;
assign a18846 = a18844 & a18810;
assign a18848 = ~a8150 & ~l1686;
assign a18850 = l1686 & l802;
assign a18852 = ~a18850 & ~a18848;
assign a18854 = a18852 & a2338;
assign a18856 = a18854 & ~a2270;
assign a18858 = l1686 & ~l794;
assign a18860 = a18858 & a18036;
assign a18862 = l1686 & ~l798;
assign a18864 = a18862 & l612;
assign a18866 = a18864 & a17890;
assign a18868 = ~a18866 & ~a18860;
assign a18870 = a18868 & ~a18856;
assign a18872 = a18870 & a18846;
assign a18874 = ~a18872 & l666;
assign a18876 = a18820 & a18076;
assign a18878 = a18828 & a2270;
assign a18880 = ~a18878 & ~a18876;
assign a18882 = a18834 & a18082;
assign a18884 = ~a18882 & a18880;
assign a18886 = ~a18854 & ~a18806;
assign a18888 = ~a18886 & a2270;
assign a18890 = ~a18888 & a18884;
assign a18892 = a18800 & a6648;
assign a18894 = a18864 & a17886;
assign a18896 = ~a18894 & ~a18892;
assign a18898 = a18838 & a18058;
assign a18900 = ~a18898 & a18896;
assign a18902 = a18858 & a17906;
assign a18904 = a18816 & a18048;
assign a18906 = ~a18904 & ~a18902;
assign a18908 = a18906 & a18900;
assign a18910 = a18908 & a18890;
assign a18912 = ~a18910 & ~l666;
assign a18914 = ~a18912 & ~a18874;
assign a18916 = ~a18914 & a16090;
assign a18918 = ~a18916 & ~a18798;
assign a18920 = a18914 & ~a16090;
assign a18922 = ~a18920 & ~a18918;
assign a18924 = l1686 & ~l778;
assign a18926 = a18924 & a18088;
assign a18928 = l1686 & ~l782;
assign a18930 = a18928 & a2370;
assign a18932 = a18930 & ~a2270;
assign a18934 = ~a18932 & ~a18926;
assign a18936 = l1686 & l770;
assign a18938 = ~a18936 & ~a10374;
assign a18940 = a18938 & ~a2302;
assign a18942 = a18940 & a18074;
assign a18944 = l1686 & ~l788;
assign a18946 = a18944 & a6648;
assign a18948 = ~a18946 & ~a18942;
assign a18950 = l1686 & ~l786;
assign a18952 = a18950 & a18040;
assign a18954 = a18952 & ~a2270;
assign a18956 = ~a18954 & a18948;
assign a18958 = l1686 & ~l784;
assign a18960 = a18958 & a18042;
assign a18962 = l1686 & ~l774;
assign a18964 = a18962 & a17906;
assign a18966 = ~a18964 & ~a18960;
assign a18968 = a18966 & a18956;
assign a18970 = a18968 & a18934;
assign a18972 = ~a8170 & ~l1686;
assign a18974 = l1686 & l780;
assign a18976 = ~a18974 & ~a18972;
assign a18978 = a18976 & a2338;
assign a18980 = a18978 & ~a2270;
assign a18982 = l1686 & ~l772;
assign a18984 = a18982 & a18036;
assign a18986 = l1686 & ~l776;
assign a18988 = a18986 & l612;
assign a18990 = a18988 & a17890;
assign a18992 = ~a18990 & ~a18984;
assign a18994 = a18992 & ~a18980;
assign a18996 = a18994 & a18970;
assign a18998 = ~a18996 & l666;
assign a19000 = a18944 & a18076;
assign a19002 = a18952 & a2270;
assign a19004 = ~a19002 & ~a19000;
assign a19006 = a18958 & a18082;
assign a19008 = ~a19006 & a19004;
assign a19010 = ~a18978 & ~a18930;
assign a19012 = ~a19010 & a2270;
assign a19014 = ~a19012 & a19008;
assign a19016 = a18924 & a6648;
assign a19018 = a18988 & a17886;
assign a19020 = ~a19018 & ~a19016;
assign a19022 = a18962 & a18058;
assign a19024 = ~a19022 & a19020;
assign a19026 = a18982 & a17906;
assign a19028 = a18940 & a18048;
assign a19030 = ~a19028 & ~a19026;
assign a19032 = a19030 & a19024;
assign a19034 = a19032 & a19014;
assign a19036 = ~a19034 & ~l666;
assign a19038 = ~a19036 & ~a18998;
assign a19040 = ~a19038 & a16080;
assign a19042 = ~a19040 & ~a18922;
assign a19044 = a19038 & ~a16080;
assign a19046 = ~a19044 & ~a19042;
assign a19048 = l1686 & ~l756;
assign a19050 = a19048 & a18088;
assign a19052 = l1686 & ~l760;
assign a19054 = a19052 & a2370;
assign a19056 = a19054 & ~a2270;
assign a19058 = ~a19056 & ~a19050;
assign a19060 = l1686 & l748;
assign a19062 = ~a19060 & ~a10436;
assign a19064 = a19062 & ~a2302;
assign a19066 = a19064 & a18074;
assign a19068 = l1686 & ~l766;
assign a19070 = a19068 & a6648;
assign a19072 = ~a19070 & ~a19066;
assign a19074 = l1686 & ~l764;
assign a19076 = a19074 & a18040;
assign a19078 = a19076 & ~a2270;
assign a19080 = ~a19078 & a19072;
assign a19082 = l1686 & ~l762;
assign a19084 = a19082 & a18042;
assign a19086 = l1686 & ~l752;
assign a19088 = a19086 & a17906;
assign a19090 = ~a19088 & ~a19084;
assign a19092 = a19090 & a19080;
assign a19094 = a19092 & a19058;
assign a19096 = ~a8190 & ~l1686;
assign a19098 = l1686 & l758;
assign a19100 = ~a19098 & ~a19096;
assign a19102 = a19100 & a2338;
assign a19104 = a19102 & ~a2270;
assign a19106 = l1686 & ~l750;
assign a19108 = a19106 & a18036;
assign a19110 = l1686 & ~l754;
assign a19112 = a19110 & l612;
assign a19114 = a19112 & a17890;
assign a19116 = ~a19114 & ~a19108;
assign a19118 = a19116 & ~a19104;
assign a19120 = a19118 & a19094;
assign a19122 = ~a19120 & l666;
assign a19124 = a19068 & a18076;
assign a19126 = a19076 & a2270;
assign a19128 = ~a19126 & ~a19124;
assign a19130 = a19082 & a18082;
assign a19132 = ~a19130 & a19128;
assign a19134 = ~a19102 & ~a19054;
assign a19136 = ~a19134 & a2270;
assign a19138 = ~a19136 & a19132;
assign a19140 = a19048 & a6648;
assign a19142 = a19112 & a17886;
assign a19144 = ~a19142 & ~a19140;
assign a19146 = a19086 & a18058;
assign a19148 = ~a19146 & a19144;
assign a19150 = a19106 & a17906;
assign a19152 = a19064 & a18048;
assign a19154 = ~a19152 & ~a19150;
assign a19156 = a19154 & a19148;
assign a19158 = a19156 & a19138;
assign a19160 = ~a19158 & ~l666;
assign a19162 = ~a19160 & ~a19122;
assign a19164 = ~a19162 & a16070;
assign a19166 = ~a19164 & ~a19046;
assign a19168 = a19162 & ~a16070;
assign a19170 = ~a19168 & ~a19166;
assign a19172 = ~a18428 & a16052;
assign a19174 = ~a19172 & ~a19170;
assign a19176 = ~a19174 & a18432;
assign a19178 = ~a19176 & ~a18198;
assign a19180 = ~a19172 & ~a18314;
assign a19182 = a18548 & ~a16120;
assign a19184 = ~a19182 & ~a18672;
assign a19186 = ~a19184 & ~a18668;
assign a19188 = ~a19186 & ~a18796;
assign a19190 = ~a19188 & ~a18792;
assign a19192 = ~a19190 & ~a18920;
assign a19194 = ~a19192 & ~a18916;
assign a19196 = ~a19194 & ~a19044;
assign a19198 = ~a19196 & ~a19040;
assign a19200 = ~a19198 & ~a19168;
assign a19202 = ~a19200 & ~a19164;
assign a19204 = ~a19202 & ~a18430;
assign a19206 = ~a19204 & a19180;
assign a19210 = i156 & ~i62;
assign a19212 = a19210 & ~l1686;
assign a19214 = l1686 & l698;
assign a19216 = ~a19214 & ~a19212;
assign a19218 = l1686 & ~l692;
assign a19220 = l1686 & l688;
assign a19222 = ~a19220 & ~a13698;
assign a19224 = l1686 & ~l690;
assign a19226 = ~a19224 & ~a19222;
assign a19228 = a19226 & a19218;
assign a19230 = l1686 & l694;
assign a19232 = ~a19230 & ~a13704;
assign a19234 = ~l1686 & i62;
assign a19236 = l1686 & l696;
assign a19238 = ~a19236 & ~a19234;
assign a19240 = ~a19238 & ~a19232;
assign a19242 = a19240 & a19228;
assign a19244 = a19242 & ~a19216;
assign a19246 = ~a19242 & a17934;
assign a19250 = ~a19238 & a19232;
assign a19252 = a19250 & ~a19218;
assign a19254 = a19252 & a19224;
assign a19256 = a19254 & a19222;
assign a19258 = a19256 & ~a19216;
assign a19260 = ~a19256 & a17944;
assign a19264 = a19240 & ~a19218;
assign a19266 = a19264 & ~a19222;
assign a19268 = a19266 & ~a19224;
assign a19270 = a19268 & ~a19216;
assign a19272 = ~a19268 & a17962;
assign a19276 = a19250 & a19228;
assign a19278 = a19276 & ~a19216;
assign a19280 = ~a19276 & a17992;
assign a19284 = a19264 & a19222;
assign a19286 = a19284 & ~a19224;
assign a19288 = a19286 & ~a19216;
assign a19290 = ~a19286 & a18012;
assign a19294 = a19254 & ~a19222;
assign a19296 = a19294 & ~a19216;
assign a19298 = ~a19294 & a17986;
assign a19302 = a19266 & a19224;
assign a19304 = a19302 & ~a19216;
assign a19306 = ~a19302 & a17926;
assign a19310 = a19252 & ~a19224;
assign a19312 = a19310 & ~a19222;
assign a19314 = a19312 & ~a19216;
assign a19316 = ~a19312 & a18004;
assign a19320 = a19284 & a19224;
assign a19322 = a19320 & ~a19216;
assign a19324 = ~a19320 & a17956;
assign a19328 = a19310 & a19222;
assign a19330 = a19328 & ~a19216;
assign a19332 = ~a19328 & a17976;
assign a19338 = a19336 & ~a16320;
assign a19340 = ~a19336 & a19222;
assign a19344 = a19336 & ~a16326;
assign a19346 = ~a19336 & a19224;
assign a19350 = a19336 & ~a16334;
assign a19352 = ~a19336 & a19218;
assign a19356 = a19336 & ~a16340;
assign a19358 = ~a19336 & a19232;
assign a19362 = l1686 & ~l702;
assign a19366 = ~a6902 & ~a5580;
assign a19368 = ~a19366 & a6714;
assign a19370 = l1686 & ~l1596;
assign a19372 = l1686 & ~l1594;
assign a19374 = l1686 & ~l1592;
assign a19376 = l1686 & ~l1590;
assign a19378 = l1686 & ~l1588;
assign a19380 = a19378 & i478;
assign a19382 = l1686 & ~l1586;
assign a19384 = a19382 & i476;
assign a19386 = l1686 & ~l1584;
assign a19388 = a19386 & i474;
assign a19390 = ~a19388 & ~a19384;
assign a19392 = ~a19382 & ~i476;
assign a19394 = ~a19392 & ~a19390;
assign a19396 = ~a19394 & ~a19380;
assign a19398 = ~a19378 & ~i478;
assign a19400 = ~a19398 & ~a19396;
assign a19402 = a19400 & a19376;
assign a19404 = a19402 & a19374;
assign a19406 = a19404 & a19372;
assign a19408 = ~a19406 & ~a19370;
assign a19410 = a19406 & a19370;
assign a19412 = ~a19410 & ~a19408;
assign a19414 = ~a19404 & ~a19372;
assign a19416 = ~a19414 & ~a19406;
assign a19418 = ~a19402 & ~a19374;
assign a19420 = ~a19418 & ~a19404;
assign a19422 = ~a19400 & ~a19376;
assign a19424 = ~a19422 & ~a19402;
assign a19426 = ~a19398 & ~a19380;
assign a19428 = ~a19426 & ~a19394;
assign a19430 = a19426 & a19394;
assign a19432 = ~a19430 & ~a19428;
assign a19434 = ~a19392 & ~a19384;
assign a19436 = ~a19434 & ~a19388;
assign a19438 = a19434 & a19388;
assign a19440 = ~a19438 & ~a19436;
assign a19442 = ~a19386 & i474;
assign a19444 = a19386 & ~i474;
assign a19446 = ~a19444 & ~a19442;
assign a19448 = ~a19446 & a19440;
assign a19450 = a19448 & a19432;
assign a19452 = a19450 & a19424;
assign a19454 = a19452 & a19420;
assign a19456 = a19454 & a19416;
assign a19458 = a19456 & ~a19412;
assign a19460 = ~a19456 & a19412;
assign a19462 = ~a19460 & ~a19458;
assign a19464 = ~a19462 & a19366;
assign a19466 = ~a19464 & ~a19368;
assign a19468 = ~a19466 & ~a6950;
assign a19470 = a2246 & i384;
assign a19472 = a4690 & ~a2246;
assign a19476 = a19474 & ~i478;
assign a19478 = ~a19474 & i478;
assign a19480 = a2246 & i382;
assign a19482 = a4672 & ~a2246;
assign a19486 = a19484 & ~i476;
assign a19488 = ~a19484 & i476;
assign a19490 = a2246 & i202;
assign a19492 = a4656 & ~a2246;
assign a19496 = ~a19494 & i474;
assign a19498 = ~a19496 & ~a19488;
assign a19500 = ~a19498 & ~a19486;
assign a19502 = ~a19500 & ~a19478;
assign a19504 = ~a19502 & ~a19476;
assign a19506 = a2246 & i386;
assign a19508 = a4706 & ~a2246;
assign a19512 = ~a19510 & a19504;
assign a19514 = a2246 & i388;
assign a19516 = a4722 & ~a2246;
assign a19520 = ~a19518 & a19512;
assign a19522 = a2246 & i390;
assign a19524 = a4738 & ~a2246;
assign a19528 = ~a19526 & a19520;
assign a19530 = a2246 & i354;
assign a19532 = a4752 & ~a2246;
assign a19536 = a19534 & ~a19528;
assign a19538 = ~a19534 & a19528;
assign a19540 = ~a19538 & ~a19536;
assign a19542 = a19540 & a6950;
assign a19544 = ~a19542 & ~a19468;
assign a19546 = ~a19544 & ~a6906;
assign a19548 = a6806 & i478;
assign a19550 = a6834 & i476;
assign a19552 = a6852 & i474;
assign a19554 = ~a19552 & ~a19550;
assign a19556 = ~a6834 & ~i476;
assign a19558 = ~a19556 & ~a19554;
assign a19560 = ~a19558 & ~a19548;
assign a19562 = ~a6806 & ~i478;
assign a19564 = ~a19562 & ~a19560;
assign a19566 = a19564 & a6744;
assign a19568 = a19566 & a6726;
assign a19570 = a19568 & a6720;
assign a19572 = ~a19570 & ~a6714;
assign a19574 = a19570 & a6714;
assign a19576 = ~a19574 & ~a19572;
assign a19578 = ~a19568 & ~a6720;
assign a19580 = ~a19578 & ~a19570;
assign a19582 = ~a19566 & ~a6726;
assign a19584 = ~a19582 & ~a19568;
assign a19586 = ~a19564 & ~a6744;
assign a19588 = ~a19586 & ~a19566;
assign a19590 = ~a19562 & ~a19548;
assign a19592 = ~a19590 & ~a19558;
assign a19594 = a19590 & a19558;
assign a19596 = ~a19594 & ~a19592;
assign a19598 = ~a19556 & ~a19550;
assign a19600 = ~a19598 & ~a19552;
assign a19602 = a19598 & a19552;
assign a19604 = ~a19602 & ~a19600;
assign a19606 = ~a6852 & i474;
assign a19608 = a6852 & ~i474;
assign a19610 = ~a19608 & ~a19606;
assign a19612 = ~a19610 & a19604;
assign a19614 = a19612 & a19596;
assign a19616 = a19614 & a19588;
assign a19618 = a19616 & a19584;
assign a19620 = a19618 & a19580;
assign a19622 = a19620 & ~a19576;
assign a19624 = ~a19620 & a19576;
assign a19626 = ~a19624 & ~a19622;
assign a19628 = ~a19626 & a6906;
assign a19632 = ~a19630 & ~a5396;
assign a19634 = a19630 & a5396;
assign a19636 = ~a19366 & a6720;
assign a19638 = ~a19454 & ~a19416;
assign a19640 = ~a19638 & ~a19456;
assign a19642 = a19640 & a19366;
assign a19644 = ~a19642 & ~a19636;
assign a19646 = ~a19644 & ~a6950;
assign a19648 = a19526 & ~a19520;
assign a19650 = ~a19648 & ~a19528;
assign a19652 = a19650 & a6950;
assign a19654 = ~a19652 & ~a19646;
assign a19656 = ~a19654 & ~a6906;
assign a19658 = ~a19618 & ~a19580;
assign a19660 = ~a19658 & ~a19620;
assign a19662 = a19660 & a6906;
assign a19666 = ~a19664 & ~a5394;
assign a19668 = a19664 & a5394;
assign a19670 = ~a19366 & a6726;
assign a19672 = ~a19452 & ~a19420;
assign a19674 = ~a19672 & ~a19454;
assign a19676 = a19674 & a19366;
assign a19678 = ~a19676 & ~a19670;
assign a19680 = ~a19678 & ~a6950;
assign a19682 = a19518 & ~a19512;
assign a19684 = ~a19682 & ~a19520;
assign a19686 = a19684 & a6950;
assign a19688 = ~a19686 & ~a19680;
assign a19690 = ~a19688 & ~a6906;
assign a19692 = ~a19616 & ~a19584;
assign a19694 = ~a19692 & ~a19618;
assign a19696 = a19694 & a6906;
assign a19700 = ~a19698 & ~a5392;
assign a19702 = a19698 & a5392;
assign a19704 = ~a19366 & a6744;
assign a19706 = ~a19450 & ~a19424;
assign a19708 = ~a19706 & ~a19452;
assign a19710 = a19708 & a19366;
assign a19712 = ~a19710 & ~a19704;
assign a19714 = ~a19712 & ~a6950;
assign a19716 = a19510 & ~a19504;
assign a19718 = ~a19716 & ~a19512;
assign a19720 = a19718 & a6950;
assign a19722 = ~a19720 & ~a19714;
assign a19724 = ~a19722 & ~a6906;
assign a19726 = ~a19614 & ~a19588;
assign a19728 = ~a19726 & ~a19616;
assign a19730 = a19728 & a6906;
assign a19734 = ~a19732 & ~a5384;
assign a19736 = a19732 & a5384;
assign a19738 = ~a19366 & a6806;
assign a19740 = ~a19448 & ~a19432;
assign a19742 = ~a19740 & ~a19450;
assign a19744 = a19742 & a19366;
assign a19746 = ~a19744 & ~a19738;
assign a19748 = ~a19746 & ~a6950;
assign a19750 = ~a19478 & ~a19476;
assign a19752 = ~a19750 & a19500;
assign a19754 = a19750 & ~a19500;
assign a19756 = ~a19754 & ~a19752;
assign a19758 = ~a19756 & a6950;
assign a19760 = ~a19758 & ~a19748;
assign a19762 = ~a19760 & ~a6906;
assign a19764 = ~a19612 & ~a19596;
assign a19766 = ~a19764 & ~a19614;
assign a19768 = a19766 & a6906;
assign a19772 = ~a19770 & ~a5376;
assign a19774 = a19770 & a5376;
assign a19776 = ~a19366 & a6834;
assign a19778 = a19446 & ~a19440;
assign a19780 = ~a19778 & ~a19448;
assign a19782 = a19780 & a19366;
assign a19784 = ~a19782 & ~a19776;
assign a19786 = ~a19784 & ~a6950;
assign a19788 = ~a19488 & ~a19486;
assign a19790 = ~a19788 & a19496;
assign a19792 = a19788 & ~a19496;
assign a19794 = ~a19792 & ~a19790;
assign a19796 = ~a19794 & a6950;
assign a19798 = ~a19796 & ~a19786;
assign a19800 = ~a19798 & ~a6906;
assign a19802 = a19610 & ~a19604;
assign a19804 = ~a19802 & ~a19612;
assign a19806 = a19804 & a6906;
assign a19810 = ~a19808 & ~a5368;
assign a19812 = a19808 & a5368;
assign a19814 = ~a19366 & a6852;
assign a19816 = a19446 & a19366;
assign a19818 = ~a19816 & ~a19814;
assign a19820 = ~a19818 & ~a6950;
assign a19822 = a19494 & ~i474;
assign a19824 = ~a19822 & ~a19496;
assign a19826 = a19824 & a6950;
assign a19828 = ~a19826 & ~a19820;
assign a19830 = ~a19828 & ~a6906;
assign a19832 = a19610 & a6906;
assign a19836 = a19834 & a5514;
assign a19838 = ~a19836 & ~a19812;
assign a19840 = ~a19838 & ~a19810;
assign a19842 = ~a19840 & ~a19774;
assign a19844 = ~a19842 & ~a19772;
assign a19846 = ~a19844 & ~a19736;
assign a19848 = ~a19846 & ~a19734;
assign a19850 = ~a19848 & ~a19702;
assign a19852 = ~a19850 & ~a19700;
assign a19854 = ~a19852 & ~a19668;
assign a19856 = ~a19854 & ~a19666;
assign a19858 = ~a19856 & ~a19634;
assign a19860 = ~a19858 & ~a19632;
assign a19862 = ~a19366 & a6882;
assign a19864 = l1686 & ~l1598;
assign a19866 = a19456 & ~a19408;
assign a19868 = ~a19866 & ~a19410;
assign a19870 = ~a19868 & a19864;
assign a19872 = a19868 & ~a19864;
assign a19874 = ~a19872 & ~a19870;
assign a19876 = a19874 & a19366;
assign a19878 = ~a19876 & ~a19862;
assign a19880 = ~a19878 & ~a6950;
assign a19882 = a2246 & i200;
assign a19884 = a4760 & ~a2246;
assign a19888 = a19886 & a19538;
assign a19890 = ~a19886 & ~a19538;
assign a19892 = ~a19890 & ~a19888;
assign a19894 = ~a19892 & a6950;
assign a19896 = ~a19894 & ~a19880;
assign a19898 = ~a19896 & ~a6906;
assign a19900 = a19620 & ~a19572;
assign a19902 = ~a19900 & ~a19574;
assign a19904 = ~a19902 & a6882;
assign a19906 = a19902 & ~a6882;
assign a19908 = ~a19906 & ~a19904;
assign a19910 = a19908 & a6906;
assign a19914 = a19912 & a5398;
assign a19916 = ~a19912 & ~a5398;
assign a19918 = ~a19916 & ~a19914;
assign a19920 = ~a19918 & ~a19860;
assign a19922 = a19918 & a19860;
assign a19928 = a8500 & ~l1686;
assign a19930 = l1686 & l1582;
assign a19932 = ~a19930 & ~a19928;
assign a19934 = a19932 & a19312;
assign a19936 = ~a19312 & a18328;
assign a19940 = a19932 & a19302;
assign a19942 = ~a19302 & a18372;
assign a19946 = a19932 & a19294;
assign a19948 = ~a19294 & a18352;
assign a19952 = a19932 & a19328;
assign a19954 = ~a19328 & a18376;
assign a19958 = a19932 & a19276;
assign a19960 = ~a19276 & a18316;
assign a19964 = a19932 & a19286;
assign a19966 = ~a19286 & a18366;
assign a19970 = a19932 & a19242;
assign a19972 = ~a19242 & a18320;
assign a19976 = a19932 & a19256;
assign a19978 = ~a19256 & a18348;
assign a19982 = a19932 & a19320;
assign a19984 = ~a19320 & a18340;
assign a19988 = a19932 & a19268;
assign a19990 = ~a19268 & a18334;
assign a19994 = a8460 & ~l1686;
assign a19996 = l1686 & l1580;
assign a19998 = ~a19996 & ~a19994;
assign a20000 = a19998 & a19312;
assign a20002 = ~a19312 & a19062;
assign a20006 = a19998 & a19302;
assign a20008 = ~a19302 & a19106;
assign a20012 = a19998 & a19294;
assign a20014 = ~a19294 & a19086;
assign a20018 = a19998 & a19328;
assign a20020 = ~a19328 & a19110;
assign a20024 = a19998 & a19276;
assign a20026 = ~a19276 & a19048;
assign a20030 = a19998 & a19286;
assign a20032 = ~a19286 & a19100;
assign a20036 = a19998 & a19242;
assign a20038 = ~a19242 & a19052;
assign a20042 = a19998 & a19256;
assign a20044 = ~a19256 & a19082;
assign a20048 = a19998 & a19320;
assign a20050 = ~a19320 & a19074;
assign a20054 = a19998 & a19268;
assign a20056 = ~a19268 & a19068;
assign a20062 = a8420 & ~l1686;
assign a20064 = l1686 & l1578;
assign a20066 = ~a20064 & ~a20062;
assign a20068 = a20066 & a19312;
assign a20070 = ~a19312 & a18938;
assign a20074 = a20066 & a19302;
assign a20076 = ~a19302 & a18982;
assign a20080 = a20066 & a19294;
assign a20082 = ~a19294 & a18962;
assign a20086 = a20066 & a19328;
assign a20088 = ~a19328 & a18986;
assign a20092 = a20066 & a19276;
assign a20094 = ~a19276 & a18924;
assign a20098 = a20066 & a19286;
assign a20100 = ~a19286 & a18976;
assign a20104 = a20066 & a19242;
assign a20106 = ~a19242 & a18928;
assign a20110 = a20066 & a19256;
assign a20112 = ~a19256 & a18958;
assign a20116 = a20066 & a19320;
assign a20118 = ~a19320 & a18950;
assign a20122 = a20066 & a19268;
assign a20124 = ~a19268 & a18944;
assign a20130 = a8380 & ~l1686;
assign a20132 = l1686 & l1576;
assign a20134 = ~a20132 & ~a20130;
assign a20136 = a20134 & a19312;
assign a20138 = ~a19312 & a18814;
assign a20142 = a20134 & a19302;
assign a20144 = ~a19302 & a18858;
assign a20148 = a20134 & a19294;
assign a20150 = ~a19294 & a18838;
assign a20154 = a20134 & a19328;
assign a20156 = ~a19328 & a18862;
assign a20160 = a20134 & a19276;
assign a20162 = ~a19276 & a18800;
assign a20166 = a20134 & a19286;
assign a20168 = ~a19286 & a18852;
assign a20172 = a20134 & a19242;
assign a20174 = ~a19242 & a18804;
assign a20178 = a20134 & a19256;
assign a20180 = ~a19256 & a18834;
assign a20184 = a20134 & a19320;
assign a20186 = ~a19320 & a18826;
assign a20190 = a20134 & a19268;
assign a20192 = ~a19268 & a18820;
assign a20198 = a6778 & ~l1686;
assign a20200 = l1686 & l1574;
assign a20202 = ~a20200 & ~a20198;
assign a20204 = a20202 & a19312;
assign a20206 = ~a19312 & a18690;
assign a20210 = a20202 & a19302;
assign a20212 = ~a19302 & a18734;
assign a20216 = a20202 & a19294;
assign a20218 = ~a19294 & a18714;
assign a20222 = a20202 & a19328;
assign a20224 = ~a19328 & a18738;
assign a20228 = a20202 & a19276;
assign a20230 = ~a19276 & a18676;
assign a20234 = a20202 & a19286;
assign a20236 = ~a19286 & a18728;
assign a20240 = a20202 & a19242;
assign a20242 = ~a19242 & a18680;
assign a20246 = a20202 & a19256;
assign a20248 = ~a19256 & a18710;
assign a20252 = a20202 & a19320;
assign a20254 = ~a19320 & a18702;
assign a20258 = a20202 & a19268;
assign a20260 = ~a19268 & a18696;
assign a20266 = a6756 & ~l1686;
assign a20268 = l1686 & l1572;
assign a20270 = ~a20268 & ~a20266;
assign a20272 = a20270 & a19312;
assign a20274 = ~a19312 & a18566;
assign a20278 = a20270 & a19302;
assign a20280 = ~a19302 & a18610;
assign a20284 = a20270 & a19294;
assign a20286 = ~a19294 & a18590;
assign a20290 = a20270 & a19328;
assign a20292 = ~a19328 & a18614;
assign a20296 = a20270 & a19276;
assign a20298 = ~a19276 & a18552;
assign a20302 = a20270 & a19286;
assign a20304 = ~a19286 & a18604;
assign a20308 = a20270 & a19242;
assign a20310 = ~a19242 & a18556;
assign a20314 = a20270 & a19256;
assign a20316 = ~a19256 & a18586;
assign a20320 = a20270 & a19320;
assign a20322 = ~a19320 & a18578;
assign a20326 = a20270 & a19268;
assign a20328 = ~a19268 & a18572;
assign a20334 = a6764 & ~l1686;
assign a20336 = l1686 & l938;
assign a20338 = ~a20336 & ~a20334;
assign a20340 = a20338 & a19312;
assign a20342 = ~a19312 & a18448;
assign a20346 = a20338 & a19302;
assign a20348 = ~a19302 & a18492;
assign a20352 = a20338 & a19294;
assign a20354 = ~a19294 & a18472;
assign a20358 = a20338 & a19328;
assign a20360 = ~a19328 & a18496;
assign a20364 = a20338 & a19276;
assign a20366 = ~a19276 & a18434;
assign a20370 = a20338 & a19286;
assign a20372 = ~a19286 & a18486;
assign a20376 = a20338 & a19242;
assign a20378 = ~a19242 & a18438;
assign a20382 = a20338 & a19256;
assign a20384 = ~a19256 & a18468;
assign a20388 = a20338 & a19320;
assign a20390 = ~a19320 & a18460;
assign a20394 = a20338 & a19268;
assign a20396 = ~a19268 & a18454;
assign a20400 = i198 & ~i62;
assign a20402 = ~a20400 & ~l1686;
assign a20404 = l1686 & l936;
assign a20406 = ~a20404 & ~a20402;
assign a20408 = a20406 & a19312;
assign a20410 = ~a19312 & a18212;
assign a20414 = a20406 & a19302;
assign a20416 = ~a19302 & a18252;
assign a20420 = a20406 & a19294;
assign a20422 = ~a19294 & a18236;
assign a20426 = a20406 & a19328;
assign a20428 = ~a19328 & a18256;
assign a20432 = a20406 & a19276;
assign a20434 = ~a19276 & a18200;
assign a20438 = a20406 & a19286;
assign a20440 = ~a19286 & a18246;
assign a20444 = a20406 & a19242;
assign a20446 = ~a19242 & a18204;
assign a20450 = a20406 & a19256;
assign a20452 = ~a19256 & a18232;
assign a20456 = a20406 & a19320;
assign a20458 = ~a19320 & a18224;
assign a20462 = a20406 & a19268;
assign a20464 = ~a19268 & a18218;
assign a20468 = ~a19286 & a18126;
assign a20470 = ~a20468 & ~l494;
assign a20472 = a18036 & l666;
assign a20474 = ~a20472 & a20470;
assign a20476 = l1686 & ~l926;
assign a20478 = ~a20476 & a19222;
assign a20480 = a20478 & ~a19224;
assign a20482 = l1686 & ~l924;
assign a20484 = a20482 & l690;
assign a20486 = a20484 & a19222;
assign a20488 = ~a20486 & ~a20480;
assign a20490 = a20476 & a19222;
assign a20492 = l1686 & ~l920;
assign a20494 = a20492 & ~a19232;
assign a20496 = a20494 & ~a20482;
assign a20498 = a20496 & ~a19224;
assign a20500 = a20498 & a20490;
assign a20502 = ~a20500 & a20488;
assign a20504 = l1686 & ~l922;
assign a20506 = ~a20504 & ~a20476;
assign a20508 = a20506 & a19218;
assign a20510 = ~a20492 & ~a20482;
assign a20512 = a20510 & a20508;
assign a20514 = a20504 & a19218;
assign a20516 = a20514 & a20494;
assign a20518 = ~a20516 & ~a20512;
assign a20520 = a19232 & a19218;
assign a20522 = ~a20482 & ~a20476;
assign a20524 = a20522 & ~a20504;
assign a20526 = a20524 & a20520;
assign a20528 = ~a20526 & a20518;
assign a20530 = a20482 & a19224;
assign a20532 = a20530 & a20494;
assign a20534 = a20532 & a20490;
assign a20536 = a20476 & ~a19222;
assign a20538 = a20536 & a20530;
assign a20540 = ~a20538 & ~a20534;
assign a20542 = a20532 & ~a19222;
assign a20544 = a20542 & ~a20476;
assign a20546 = ~a20544 & a20540;
assign a20548 = a20546 & a20528;
assign a20550 = a20522 & a19224;
assign a20552 = a20506 & a20496;
assign a20554 = a20552 & ~a19222;
assign a20556 = ~a20554 & ~a20550;
assign a20558 = a20556 & a20548;
assign a20560 = a20558 & a20502;
assign a20562 = ~a20560 & a6710;
assign a20566 = ~a19256 & ~l902;
assign a20568 = ~a20566 & ~l494;
assign a20570 = a2370 & l666;
assign a20572 = a20570 & a2270;
assign a20574 = ~a20572 & a20568;
assign a20576 = a20482 & l920;
assign a20578 = a20576 & a20536;
assign a20580 = a20576 & ~a19224;
assign a20582 = ~a20580 & ~a20578;
assign a20584 = ~a20492 & a19232;
assign a20586 = a20584 & a19222;
assign a20588 = a20586 & a20482;
assign a20590 = ~a20588 & a20582;
assign a20592 = a19224 & l924;
assign a20594 = a20592 & a19222;
assign a20596 = a20478 & a19224;
assign a20598 = ~a20596 & ~a20594;
assign a20600 = ~a20598 & a19232;
assign a20602 = ~a20600 & a20590;
assign a20604 = a20484 & ~a20476;
assign a20606 = ~a20604 & ~a20544;
assign a20608 = ~a20504 & ~a19222;
assign a20610 = a20608 & a20498;
assign a20612 = a20536 & ~a19224;
assign a20614 = a20612 & a20510;
assign a20616 = ~a20614 & ~a20610;
assign a20618 = a20616 & a20528;
assign a20620 = a19232 & a19226;
assign a20622 = a20476 & l924;
assign a20624 = a20622 & a20620;
assign a20626 = ~a20624 & ~a20500;
assign a20628 = a20626 & a20618;
assign a20630 = a20628 & a20606;
assign a20632 = a20630 & a20602;
assign a20634 = ~a20632 & a6710;
assign a20638 = ~a19328 & ~l904;
assign a20640 = ~a20638 & ~l494;
assign a20642 = a17906 & l666;
assign a20644 = ~a20642 & a20640;
assign a20646 = a20480 & a19232;
assign a20648 = a20510 & a19224;
assign a20650 = ~a20648 & ~a20614;
assign a20652 = a20650 & ~a20646;
assign a20654 = a20586 & ~a19224;
assign a20656 = a20486 & a19232;
assign a20658 = ~a20656 & ~a20654;
assign a20660 = a20658 & a20652;
assign a20662 = a20660 & a20558;
assign a20664 = ~a20662 & a6710;
assign a20668 = ~a19276 & ~l906;
assign a20670 = ~a20668 & ~l494;
assign a20672 = a2270 & l666;
assign a20674 = a20672 & ~a2302;
assign a20676 = a20674 & a2296;
assign a20678 = ~a20676 & a20670;
assign a20680 = a20484 & a19232;
assign a20682 = a20504 & l692;
assign a20684 = a20682 & ~a20492;
assign a20686 = ~a20684 & ~a20680;
assign a20688 = a20686 & ~a20526;
assign a20690 = a20584 & a19218;
assign a20692 = ~a20690 & ~a20624;
assign a20694 = a20692 & a20688;
assign a20696 = a20608 & a20494;
assign a20698 = a20696 & ~a19224;
assign a20700 = ~a20698 & ~a20484;
assign a20702 = ~a20700 & ~a19218;
assign a20704 = a20612 & ~a19218;
assign a20706 = ~a20704 & ~a20702;
assign a20708 = a20546 & ~a20500;
assign a20710 = a20708 & a20706;
assign a20712 = a20710 & a20694;
assign a20714 = ~a20712 & a6710;
assign a20718 = ~a19312 & a18104;
assign a20720 = ~a20718 & ~l494;
assign a20722 = a20674 & a17888;
assign a20724 = ~a20722 & a20720;
assign a20726 = a19232 & ~a19218;
assign a20728 = ~a20726 & a19226;
assign a20730 = ~a20728 & a20504;
assign a20732 = ~a20730 & ~a20486;
assign a20734 = ~a20492 & ~a20476;
assign a20736 = a20734 & ~a19224;
assign a20738 = ~a20736 & ~a20484;
assign a20740 = ~a20738 & a20726;
assign a20742 = ~a20740 & a20732;
assign a20744 = a20648 & ~a20476;
assign a20746 = a20736 & a19222;
assign a20748 = ~a20746 & ~a20744;
assign a20750 = a20748 & a20742;
assign a20752 = a20704 & a19232;
assign a20754 = ~a20752 & a20518;
assign a20756 = a20754 & a20708;
assign a20758 = a20756 & a20750;
assign a20760 = ~a20758 & a6710;
assign a20764 = ~a19294 & ~l910;
assign a20766 = ~a20764 & ~l494;
assign a20768 = a20672 & a18040;
assign a20770 = ~a20768 & a20766;
assign a20772 = a20580 & ~a20476;
assign a20774 = ~a20772 & ~a20534;
assign a20776 = a20596 & ~a20492;
assign a20778 = ~a20776 & a20774;
assign a20780 = ~a20536 & a20482;
assign a20782 = ~a20780 & a19232;
assign a20784 = a20782 & a19224;
assign a20786 = a19224 & ~a19222;
assign a20788 = a20786 & a20584;
assign a20790 = ~a20788 & ~a20594;
assign a20792 = a20790 & ~a20784;
assign a20794 = a20792 & a20778;
assign a20796 = a20794 & a20628;
assign a20798 = ~a20796 & a6710;
assign a20802 = ~a19320 & ~l912;
assign a20804 = ~a20802 & ~l494;
assign a20806 = a20570 & ~a2270;
assign a20808 = ~a20806 & a20804;
assign a20810 = a20598 & ~a20534;
assign a20812 = a20810 & a20630;
assign a20814 = ~a20812 & a6710;
assign a20818 = ~a19242 & ~a18144;
assign a20820 = a6648 & l666;
assign a20822 = ~a20820 & ~a20818;
assign a20824 = a20476 & a19218;
assign a20826 = ~a20824 & ~a20484;
assign a20828 = a20826 & ~a20526;
assign a20830 = a20828 & a20616;
assign a20832 = a20830 & a20756;
assign a20834 = ~a20832 & a6710;
assign a20838 = ~a19302 & ~l916;
assign a20840 = ~a20838 & ~l494;
assign a20842 = ~a2270 & l666;
assign a20844 = a20842 & a18040;
assign a20846 = ~a20844 & a20840;
assign a20848 = ~a20592 & a20546;
assign a20850 = a20848 & a20628;
assign a20852 = ~a20850 & a6710;
assign a20856 = ~a19268 & a18136;
assign a20858 = ~a20856 & ~l494;
assign a20860 = a20842 & a2338;
assign a20862 = ~a20860 & a20858;
assign a20864 = ~a20682 & ~a20516;
assign a20866 = a20864 & a20710;
assign a20868 = ~a20866 & a6710;
assign a20872 = l1686 & ~l934;
assign a20874 = l1686 & ~l932;
assign a20876 = l1686 & ~l930;
assign a20878 = l1686 & ~l928;
assign a20880 = ~a1698 & i466;
assign a20882 = a20880 & a6666;
assign a20884 = a20882 & ~l1686;
assign a20886 = l1686 & l1566;
assign a20888 = ~a20886 & ~a20884;
assign a20890 = ~a16262 & ~a13508;
assign a20892 = a20890 & ~a20888;
assign a20894 = a20892 & a16256;
assign a20896 = a20894 & a15340;
assign a20900 = ~a5130 & ~a5128;
assign a20902 = a20900 & a18366;
assign a20904 = a5124 & l498;
assign a20906 = a20904 & a20902;
assign a20908 = a18372 & l502;
assign a20910 = a20908 & a6602;
assign a20912 = ~a20910 & ~a20906;
assign a20914 = a5126 & l502;
assign a20916 = a20914 & a5130;
assign a20918 = a20916 & a5124;
assign a20920 = a20918 & a18320;
assign a20922 = ~a20920 & a20912;
assign a20924 = a5130 & l502;
assign a20926 = a20924 & a18340;
assign a20928 = a20926 & a20904;
assign a20930 = a20914 & ~a5130;
assign a20932 = a20930 & a18376;
assign a20934 = a20932 & ~a5124;
assign a20936 = ~a20934 & ~a20928;
assign a20938 = a20936 & a20922;
assign a20940 = a5130 & l498;
assign a20942 = a20940 & a18352;
assign a20944 = a20916 & a18348;
assign a20946 = ~a20944 & ~a20942;
assign a20948 = a5128 & l496;
assign a20950 = a20948 & a18316;
assign a20952 = a6558 & ~a5130;
assign a20954 = a20952 & a18328;
assign a20956 = ~a20954 & ~a20950;
assign a20958 = a20956 & a20946;
assign a20960 = ~a20958 & ~a5124;
assign a20962 = a18334 & l496;
assign a20964 = a20962 & a6434;
assign a20966 = ~a20964 & ~a20960;
assign a20968 = a20966 & a20938;
assign a20970 = a20968 & ~a16298;
assign a20972 = ~a20968 & a16298;
assign a20974 = a20900 & a19100;
assign a20976 = a20974 & a20904;
assign a20978 = a19106 & l502;
assign a20980 = a20978 & a6602;
assign a20982 = ~a20980 & ~a20976;
assign a20984 = a20918 & a19052;
assign a20986 = ~a20984 & a20982;
assign a20988 = a20924 & a19074;
assign a20990 = a20988 & a20904;
assign a20992 = a20930 & a19110;
assign a20994 = a20992 & ~a5124;
assign a20996 = ~a20994 & ~a20990;
assign a20998 = a20996 & a20986;
assign a21000 = a20940 & a19086;
assign a21002 = a20916 & a19082;
assign a21004 = ~a21002 & ~a21000;
assign a21006 = a20948 & a19048;
assign a21008 = a20952 & a19062;
assign a21010 = ~a21008 & ~a21006;
assign a21012 = a21010 & a21004;
assign a21014 = ~a21012 & ~a5124;
assign a21016 = a19068 & l496;
assign a21018 = a21016 & a6434;
assign a21020 = ~a21018 & ~a21014;
assign a21022 = a21020 & a20998;
assign a21024 = a21022 & ~a16292;
assign a21026 = ~a21022 & a16292;
assign a21028 = a20900 & a18976;
assign a21030 = a21028 & a20904;
assign a21032 = a18982 & l502;
assign a21034 = a21032 & a6602;
assign a21036 = ~a21034 & ~a21030;
assign a21038 = a20918 & a18928;
assign a21040 = ~a21038 & a21036;
assign a21042 = a20924 & a18950;
assign a21044 = a21042 & a20904;
assign a21046 = a20930 & a18986;
assign a21048 = a21046 & ~a5124;
assign a21050 = ~a21048 & ~a21044;
assign a21052 = a21050 & a21040;
assign a21054 = a20940 & a18962;
assign a21056 = a20916 & a18958;
assign a21058 = ~a21056 & ~a21054;
assign a21060 = a20948 & a18924;
assign a21062 = a20952 & a18938;
assign a21064 = ~a21062 & ~a21060;
assign a21066 = a21064 & a21058;
assign a21068 = ~a21066 & ~a5124;
assign a21070 = a18944 & l496;
assign a21072 = a21070 & a6434;
assign a21074 = ~a21072 & ~a21068;
assign a21076 = a21074 & a21052;
assign a21078 = a21076 & ~a16286;
assign a21080 = ~a21076 & a16286;
assign a21082 = a20900 & a18852;
assign a21084 = a21082 & a20904;
assign a21086 = a18858 & l502;
assign a21088 = a21086 & a6602;
assign a21090 = ~a21088 & ~a21084;
assign a21092 = a20918 & a18804;
assign a21094 = ~a21092 & a21090;
assign a21096 = a20924 & a18826;
assign a21098 = a21096 & a20904;
assign a21100 = a20930 & a18862;
assign a21102 = a21100 & ~a5124;
assign a21104 = ~a21102 & ~a21098;
assign a21106 = a21104 & a21094;
assign a21108 = a20940 & a18838;
assign a21110 = a20916 & a18834;
assign a21112 = ~a21110 & ~a21108;
assign a21114 = a20948 & a18800;
assign a21116 = a20952 & a18814;
assign a21118 = ~a21116 & ~a21114;
assign a21120 = a21118 & a21112;
assign a21122 = ~a21120 & ~a5124;
assign a21124 = a18820 & l496;
assign a21126 = a21124 & a6434;
assign a21128 = ~a21126 & ~a21122;
assign a21130 = a21128 & a21106;
assign a21132 = a21130 & ~a16280;
assign a21134 = ~a21130 & a16280;
assign a21136 = a20900 & a18728;
assign a21138 = a21136 & a20904;
assign a21140 = a18734 & l502;
assign a21142 = a21140 & a6602;
assign a21144 = ~a21142 & ~a21138;
assign a21146 = a20918 & a18680;
assign a21148 = ~a21146 & a21144;
assign a21150 = a20924 & a18702;
assign a21152 = a21150 & a20904;
assign a21154 = a20930 & a18738;
assign a21156 = a21154 & ~a5124;
assign a21158 = ~a21156 & ~a21152;
assign a21160 = a21158 & a21148;
assign a21162 = a20940 & a18714;
assign a21164 = a20916 & a18710;
assign a21166 = ~a21164 & ~a21162;
assign a21168 = a20948 & a18676;
assign a21170 = a20952 & a18690;
assign a21172 = ~a21170 & ~a21168;
assign a21174 = a21172 & a21166;
assign a21176 = ~a21174 & ~a5124;
assign a21178 = a18696 & l496;
assign a21180 = a21178 & a6434;
assign a21182 = ~a21180 & ~a21176;
assign a21184 = a21182 & a21160;
assign a21186 = a21184 & ~a16274;
assign a21188 = ~a21184 & a16274;
assign a21190 = a20924 & a18578;
assign a21192 = a21190 & a20904;
assign a21194 = a20940 & a18590;
assign a21196 = a21194 & ~a5124;
assign a21198 = ~a21196 & ~a21192;
assign a21200 = a18610 & l502;
assign a21202 = a21200 & a6602;
assign a21204 = a20900 & a18604;
assign a21206 = a21204 & a20904;
assign a21208 = ~a21206 & ~a21202;
assign a21210 = a21208 & a21198;
assign a21212 = a20918 & a18556;
assign a21214 = a20916 & a18586;
assign a21216 = a21214 & ~a5124;
assign a21218 = ~a21216 & ~a21212;
assign a21220 = a21218 & a21210;
assign a21222 = a20952 & a18566;
assign a21224 = a20930 & a18614;
assign a21226 = ~a21224 & ~a21222;
assign a21228 = ~a21226 & ~a5124;
assign a21230 = a18572 & l496;
assign a21232 = a21230 & a6434;
assign a21234 = a20948 & ~a5124;
assign a21236 = a21234 & a18552;
assign a21238 = ~a21236 & ~a21232;
assign a21240 = a21238 & ~a21228;
assign a21242 = a21240 & a21220;
assign a21244 = a21242 & ~a16268;
assign a21246 = ~a21242 & a16268;
assign a21248 = a20924 & a18460;
assign a21250 = a21248 & a20904;
assign a21252 = a20940 & a18472;
assign a21254 = a21252 & ~a5124;
assign a21256 = ~a21254 & ~a21250;
assign a21258 = a18492 & l502;
assign a21260 = a21258 & a6602;
assign a21262 = a20900 & a18486;
assign a21264 = a21262 & a20904;
assign a21266 = ~a21264 & ~a21260;
assign a21268 = a21266 & a21256;
assign a21270 = a20918 & a18438;
assign a21272 = a20916 & a18468;
assign a21274 = a21272 & ~a5124;
assign a21276 = ~a21274 & ~a21270;
assign a21278 = a21276 & a21268;
assign a21280 = a20952 & a18448;
assign a21282 = a20930 & a18496;
assign a21284 = ~a21282 & ~a21280;
assign a21286 = ~a21284 & ~a5124;
assign a21288 = a18454 & l496;
assign a21290 = a21288 & a6434;
assign a21292 = a21234 & a18434;
assign a21294 = ~a21292 & ~a21290;
assign a21296 = a21294 & ~a21286;
assign a21298 = a21296 & a21278;
assign a21300 = ~a21298 & a16310;
assign a21302 = ~a21300 & ~a21246;
assign a21304 = ~a21302 & ~a21244;
assign a21306 = ~a21304 & ~a21188;
assign a21308 = ~a21306 & ~a21186;
assign a21310 = ~a21308 & ~a21134;
assign a21312 = ~a21310 & ~a21132;
assign a21314 = ~a21312 & ~a21080;
assign a21316 = ~a21314 & ~a21078;
assign a21318 = ~a21316 & ~a21026;
assign a21320 = ~a21318 & ~a21024;
assign a21322 = ~a21320 & ~a20972;
assign a21324 = ~a21322 & ~a20970;
assign a21326 = a18252 & l502;
assign a21328 = a20940 & ~a5124;
assign a21330 = a21328 & a21326;
assign a21332 = a21234 & a18204;
assign a21334 = ~a21332 & ~a21330;
assign a21336 = a20900 & a18246;
assign a21338 = a21336 & a6556;
assign a21340 = a18218 & l496;
assign a21342 = a6558 & ~a5124;
assign a21344 = a21342 & a21340;
assign a21346 = ~a21344 & ~a21338;
assign a21348 = a21346 & a21334;
assign a21350 = a20940 & a18236;
assign a21352 = a20916 & a18232;
assign a21354 = ~a21352 & ~a21350;
assign a21356 = ~a21354 & a5124;
assign a21358 = ~a21356 & a21348;
assign a21360 = a18200 & a6436;
assign a21362 = a20924 & a18224;
assign a21364 = a21362 & a6556;
assign a21366 = ~a21364 & ~a21360;
assign a21368 = a20952 & a18212;
assign a21370 = a20930 & a18256;
assign a21372 = ~a21370 & ~a21368;
assign a21374 = ~a21372 & a5124;
assign a21376 = ~a21374 & a21366;
assign a21378 = a21376 & a21358;
assign a21380 = ~a21378 & a16304;
assign a21382 = a21378 & ~a16304;
assign a21384 = ~a21382 & ~a21380;
assign a21386 = a21328 & a20908;
assign a21388 = a21234 & a18320;
assign a21390 = ~a21388 & ~a21386;
assign a21392 = a20902 & a6556;
assign a21394 = a21342 & a20962;
assign a21396 = ~a21394 & ~a21392;
assign a21398 = a21396 & a21390;
assign a21400 = ~a20946 & a5124;
assign a21402 = ~a21400 & a21398;
assign a21404 = a20956 & ~a20932;
assign a21406 = ~a21404 & a5124;
assign a21408 = a20926 & a6556;
assign a21410 = ~a21408 & ~a21406;
assign a21412 = a21410 & a21402;
assign a21414 = a21412 & ~a16298;
assign a21416 = ~a21412 & a16298;
assign a21418 = a21328 & a20978;
assign a21420 = a21234 & a19052;
assign a21422 = ~a21420 & ~a21418;
assign a21424 = a20974 & a6556;
assign a21426 = a21342 & a21016;
assign a21428 = ~a21426 & ~a21424;
assign a21430 = a21428 & a21422;
assign a21432 = ~a21004 & a5124;
assign a21434 = ~a21432 & a21430;
assign a21436 = a21010 & ~a20992;
assign a21438 = ~a21436 & a5124;
assign a21440 = a20988 & a6556;
assign a21442 = ~a21440 & ~a21438;
assign a21444 = a21442 & a21434;
assign a21446 = a21444 & ~a16292;
assign a21448 = ~a21444 & a16292;
assign a21450 = a21328 & a21032;
assign a21452 = a21234 & a18928;
assign a21454 = ~a21452 & ~a21450;
assign a21456 = a21028 & a6556;
assign a21458 = a21342 & a21070;
assign a21460 = ~a21458 & ~a21456;
assign a21462 = a21460 & a21454;
assign a21464 = ~a21058 & a5124;
assign a21466 = ~a21464 & a21462;
assign a21468 = a21064 & ~a21046;
assign a21470 = ~a21468 & a5124;
assign a21472 = a21042 & a6556;
assign a21474 = ~a21472 & ~a21470;
assign a21476 = a21474 & a21466;
assign a21478 = a21476 & ~a16286;
assign a21480 = ~a21476 & a16286;
assign a21482 = a21328 & a21086;
assign a21484 = a21234 & a18804;
assign a21486 = ~a21484 & ~a21482;
assign a21488 = a21082 & a6556;
assign a21490 = a21342 & a21124;
assign a21492 = ~a21490 & ~a21488;
assign a21494 = a21492 & a21486;
assign a21496 = ~a21112 & a5124;
assign a21498 = ~a21496 & a21494;
assign a21500 = a21118 & ~a21100;
assign a21502 = ~a21500 & a5124;
assign a21504 = a21096 & a6556;
assign a21506 = ~a21504 & ~a21502;
assign a21508 = a21506 & a21498;
assign a21510 = a21508 & ~a16280;
assign a21512 = ~a21508 & a16280;
assign a21514 = a21328 & a21140;
assign a21516 = a21234 & a18680;
assign a21518 = ~a21516 & ~a21514;
assign a21520 = a21136 & a6556;
assign a21522 = a21342 & a21178;
assign a21524 = ~a21522 & ~a21520;
assign a21526 = a21524 & a21518;
assign a21528 = ~a21166 & a5124;
assign a21530 = ~a21528 & a21526;
assign a21532 = a21172 & ~a21154;
assign a21534 = ~a21532 & a5124;
assign a21536 = a21150 & a6556;
assign a21538 = ~a21536 & ~a21534;
assign a21540 = a21538 & a21530;
assign a21542 = a21540 & ~a16274;
assign a21544 = ~a21540 & a16274;
assign a21546 = a21328 & a21200;
assign a21548 = a21234 & a18556;
assign a21550 = ~a21548 & ~a21546;
assign a21552 = a21204 & a6556;
assign a21554 = a21342 & a21230;
assign a21556 = ~a21554 & ~a21552;
assign a21558 = a21556 & a21550;
assign a21560 = ~a21214 & ~a21194;
assign a21562 = ~a21560 & a5124;
assign a21564 = ~a21562 & a21558;
assign a21566 = a18552 & a6436;
assign a21568 = a21190 & a6556;
assign a21570 = ~a21568 & ~a21566;
assign a21572 = ~a21226 & a5124;
assign a21574 = ~a21572 & a21570;
assign a21576 = a21574 & a21564;
assign a21578 = a21576 & ~a16268;
assign a21580 = ~a21576 & a16268;
assign a21582 = a21328 & a21258;
assign a21584 = a21234 & a18438;
assign a21586 = ~a21584 & ~a21582;
assign a21588 = a21262 & a6556;
assign a21590 = a21342 & a21288;
assign a21592 = ~a21590 & ~a21588;
assign a21594 = a21592 & a21586;
assign a21596 = ~a21272 & ~a21252;
assign a21598 = ~a21596 & a5124;
assign a21600 = ~a21598 & a21594;
assign a21602 = a18434 & a6436;
assign a21604 = a21248 & a6556;
assign a21606 = ~a21604 & ~a21602;
assign a21608 = ~a21284 & a5124;
assign a21610 = ~a21608 & a21606;
assign a21612 = a21610 & a21600;
assign a21614 = ~a21612 & a16310;
assign a21616 = ~a21614 & ~a21580;
assign a21618 = ~a21616 & ~a21578;
assign a21620 = ~a21618 & ~a21544;
assign a21622 = ~a21620 & ~a21542;
assign a21624 = ~a21622 & ~a21512;
assign a21626 = ~a21624 & ~a21510;
assign a21628 = ~a21626 & ~a21480;
assign a21630 = ~a21628 & ~a21478;
assign a21632 = ~a21630 & ~a21448;
assign a21634 = ~a21632 & ~a21446;
assign a21636 = ~a21634 & ~a21416;
assign a21638 = ~a21636 & ~a21414;
assign a21640 = ~a21638 & a21384;
assign a21642 = a21640 & a21324;
assign a21644 = a21362 & a20904;
assign a21646 = a21326 & a6602;
assign a21648 = ~a21646 & ~a21644;
assign a21650 = a21336 & a20904;
assign a21652 = a21340 & a6434;
assign a21654 = ~a21652 & ~a21650;
assign a21656 = a21654 & a21648;
assign a21658 = ~a21354 & ~a5124;
assign a21660 = ~a21658 & a21656;
assign a21662 = a21234 & a18200;
assign a21664 = a20918 & a18204;
assign a21666 = ~a21664 & ~a21662;
assign a21668 = ~a21372 & ~a5124;
assign a21670 = ~a21668 & a21666;
assign a21672 = a21670 & a21660;
assign a21674 = ~a21672 & a16304;
assign a21676 = a21672 & ~a16304;
assign a21678 = ~a21676 & ~a21674;
assign a21680 = a21678 & a21324;
assign a21682 = ~a21680 & ~a21640;
assign a21684 = ~a21672 & a21378;
assign a21686 = a21672 & ~a21378;
assign a21688 = ~a21686 & ~a21684;
assign a21690 = ~a21688 & ~a21682;
assign a21692 = ~a21690 & ~a21642;
assign a21694 = l1686 & ~l1488;
assign a21696 = a21694 & ~a16262;
assign a21700 = a21698 & a21692;
assign a21702 = a5130 & l690;
assign a21704 = a19232 & ~a5124;
assign a21706 = ~a21704 & ~a21702;
assign a21708 = ~a19222 & a5126;
assign a21710 = ~a19232 & a5124;
assign a21712 = ~a21710 & ~a21708;
assign a21714 = a21712 & a21706;
assign a21716 = a19222 & ~a5126;
assign a21718 = a19224 & l496;
assign a21720 = ~a21718 & ~a21716;
assign a21722 = a19218 & l502;
assign a21724 = a5128 & l692;
assign a21726 = ~a21724 & ~a21722;
assign a21728 = a21726 & a21720;
assign a21730 = a21728 & a21714;
assign a21732 = ~a21730 & a21700;
assign a21734 = a20924 & l912;
assign a21736 = a21734 & a20904;
assign a21738 = ~a5128 & l916;
assign a21740 = a21738 & a6602;
assign a21742 = ~a21740 & ~a21736;
assign a21744 = a20900 & ~a18126;
assign a21746 = a21744 & a20904;
assign a21748 = ~a18136 & ~a5130;
assign a21750 = a21748 & a6434;
assign a21752 = ~a21750 & ~a21746;
assign a21754 = a21752 & a21742;
assign a21756 = a20940 & l910;
assign a21758 = a20916 & l902;
assign a21760 = ~a21758 & ~a21756;
assign a21762 = ~a21760 & ~a5124;
assign a21764 = ~a21762 & a21754;
assign a21766 = a20948 & l906;
assign a21768 = a20952 & ~a18104;
assign a21770 = a20930 & l904;
assign a21772 = ~a21770 & ~a21768;
assign a21774 = a21772 & ~a21766;
assign a21776 = ~a21774 & ~a5124;
assign a21778 = a20918 & a18144;
assign a21780 = ~a21778 & ~a21776;
assign a21782 = a21780 & a21764;
assign a21784 = ~a21782 & a21732;
assign a21786 = a21738 & a21328;
assign a21788 = a21234 & a18144;
assign a21790 = ~a21788 & ~a21786;
assign a21792 = a21744 & a6556;
assign a21794 = a21748 & a21342;
assign a21796 = ~a21794 & ~a21792;
assign a21798 = a21796 & a21790;
assign a21800 = ~a21760 & a5124;
assign a21802 = ~a21800 & a21798;
assign a21804 = ~a21774 & a5124;
assign a21806 = a21734 & a6556;
assign a21808 = ~a21806 & ~a21804;
assign a21810 = a21808 & a21802;
assign a21812 = ~a21810 & ~a21784;
assign a21814 = ~a10802 & ~l972;
assign a21816 = ~l1496 & ~l988;
assign a21818 = a10826 & a10744;
assign a21820 = ~a21818 & ~a10748;
assign a21822 = a21820 & i436;
assign a21824 = a10828 & ~a8032;
assign a21826 = ~a21824 & a21822;
assign a21828 = ~a10948 & ~a8054;
assign a21830 = ~a10862 & ~a8864;
assign a21832 = ~a21830 & ~a21828;
assign a21834 = a10948 & a8054;
assign a21836 = ~a10906 & ~a8052;
assign a21838 = ~a21836 & ~a21834;
assign a21840 = a21838 & a21832;
assign a21842 = a10798 & a8050;
assign a21844 = ~a10798 & ~a8050;
assign a21846 = ~a21844 & ~a21842;
assign a21848 = a10862 & a8864;
assign a21850 = a10906 & a8052;
assign a21852 = ~a21850 & ~a21848;
assign a21854 = a21852 & a21846;
assign a21856 = a21854 & a21840;
assign a21858 = ~a21856 & a21814;
assign a21860 = ~a21858 & ~a21826;
assign a21862 = a21858 & a10498;
assign a21864 = ~a21858 & i434;
assign a21866 = ~a21864 & ~a21862;
assign a21868 = ~a21866 & ~a8032;
assign a21870 = a10478 & a8032;
assign a21872 = ~a21870 & ~a21868;
assign a21874 = ~a21872 & a11614;
assign a21876 = a21872 & ~a11614;
assign a21878 = a21858 & a10440;
assign a21880 = ~a21858 & i432;
assign a21882 = ~a21880 & ~a21878;
assign a21884 = ~a21882 & ~a8032;
assign a21886 = a10416 & a8032;
assign a21888 = ~a21886 & ~a21884;
assign a21890 = ~a21888 & a11600;
assign a21892 = a21888 & ~a11600;
assign a21894 = a21858 & a10378;
assign a21896 = ~a21858 & i430;
assign a21898 = ~a21896 & ~a21894;
assign a21900 = ~a21898 & ~a8032;
assign a21902 = a10354 & a8032;
assign a21904 = ~a21902 & ~a21900;
assign a21906 = ~a21904 & a11586;
assign a21908 = a21904 & ~a11586;
assign a21910 = a21858 & a10316;
assign a21912 = ~a21858 & i428;
assign a21914 = ~a21912 & ~a21910;
assign a21916 = ~a21914 & ~a8032;
assign a21918 = a10292 & a8032;
assign a21920 = ~a21918 & ~a21916;
assign a21922 = ~a21920 & a11572;
assign a21924 = a21920 & ~a11572;
assign a21926 = a21858 & a10254;
assign a21928 = ~a21858 & i426;
assign a21930 = ~a21928 & ~a21926;
assign a21932 = ~a21930 & ~a8032;
assign a21934 = a10230 & a8032;
assign a21936 = ~a21934 & ~a21932;
assign a21938 = ~a21936 & a11558;
assign a21940 = a21936 & ~a11558;
assign a21942 = a21858 & a10204;
assign a21944 = ~a21858 & i424;
assign a21946 = ~a21944 & ~a21942;
assign a21948 = ~a21946 & ~a8032;
assign a21950 = a10188 & a8032;
assign a21952 = ~a21950 & ~a21948;
assign a21954 = ~a21952 & a11538;
assign a21956 = a21952 & ~a11538;
assign a21958 = a21858 & a10158;
assign a21960 = ~a21858 & i422;
assign a21962 = ~a21960 & ~a21958;
assign a21964 = ~a21962 & ~a8032;
assign a21966 = a10180 & a8032;
assign a21968 = ~a21966 & ~a21964;
assign a21970 = a21968 & ~a11544;
assign a21972 = ~a21970 & ~a21956;
assign a21974 = ~a21972 & ~a21954;
assign a21976 = ~a21974 & ~a21940;
assign a21978 = ~a21976 & ~a21938;
assign a21980 = ~a21978 & ~a21924;
assign a21982 = ~a21980 & ~a21922;
assign a21984 = ~a21982 & ~a21908;
assign a21986 = ~a21984 & ~a21906;
assign a21988 = ~a21986 & ~a21892;
assign a21990 = ~a21988 & ~a21890;
assign a21992 = ~a21990 & ~a21876;
assign a21994 = ~a21992 & ~a21874;
assign a21996 = a21858 & a8870;
assign a21998 = ~a21858 & i420;
assign a22000 = ~a21998 & ~a21996;
assign a22002 = ~a22000 & ~a8032;
assign a22004 = a8872 & a8032;
assign a22006 = ~a22004 & ~a22002;
assign a22008 = a22006 & ~a13194;
assign a22010 = ~a22006 & a13194;
assign a22012 = ~a22010 & ~a22008;
assign a22014 = ~a22012 & ~a21994;
assign a22016 = a22012 & a21994;
assign a22018 = ~a22016 & ~a22014;
assign a22020 = a11056 & ~a10906;
assign a22022 = ~a11056 & a10906;
assign a22024 = ~a22022 & ~a22020;
assign a22026 = ~a11066 & a10948;
assign a22028 = ~a22026 & a22024;
assign a22030 = ~a11076 & a10798;
assign a22032 = ~a22030 & a22028;
assign a22034 = a11088 & ~a10862;
assign a22036 = ~a11088 & a10862;
assign a22038 = ~a22036 & ~a22034;
assign a22040 = a11066 & ~a10948;
assign a22042 = ~a22040 & a22038;
assign a22044 = a11076 & ~a10798;
assign a22046 = ~a22044 & a22042;
assign a22048 = a22046 & a22032;
assign a22050 = a22048 & ~a22018;
assign a22052 = ~a21872 & a15956;
assign a22054 = a21872 & ~a15956;
assign a22056 = ~a21888 & a15858;
assign a22058 = a21888 & ~a15858;
assign a22060 = ~a21904 & a15760;
assign a22062 = a21904 & ~a15760;
assign a22064 = ~a21920 & a15656;
assign a22066 = a21920 & ~a15656;
assign a22068 = ~a21936 & a15552;
assign a22070 = a21936 & ~a15552;
assign a22072 = ~a21952 & a15448;
assign a22074 = a21952 & ~a15448;
assign a22076 = a21968 & ~a11380;
assign a22078 = ~a22076 & ~a22074;
assign a22080 = ~a22078 & ~a22072;
assign a22082 = ~a22080 & ~a22070;
assign a22084 = ~a22082 & ~a22068;
assign a22086 = ~a22084 & ~a22066;
assign a22088 = ~a22086 & ~a22064;
assign a22090 = ~a22088 & ~a22062;
assign a22092 = ~a22090 & ~a22060;
assign a22094 = ~a22092 & ~a22058;
assign a22096 = ~a22094 & ~a22056;
assign a22098 = ~a22096 & ~a22054;
assign a22100 = ~a22098 & ~a22052;
assign a22102 = a22006 & ~a11278;
assign a22104 = ~a22006 & a11278;
assign a22106 = ~a22104 & ~a22102;
assign a22108 = ~a22106 & ~a22100;
assign a22110 = a22106 & a22100;
assign a22112 = ~a22110 & ~a22108;
assign a22114 = ~a22112 & ~a22048;
assign a22116 = ~a22114 & ~a22050;
assign a22118 = a11752 & a10920;
assign a22120 = a11756 & ~a10920;
assign a22122 = ~a22120 & ~a22118;
assign a22124 = ~a22122 & a10962;
assign a22126 = a11768 & a10920;
assign a22128 = a11776 & ~a10920;
assign a22130 = ~a22128 & ~a22126;
assign a22132 = ~a22130 & ~a10962;
assign a22134 = ~a22132 & ~a22124;
assign a22136 = ~a22134 & a10816;
assign a22138 = a11788 & a10920;
assign a22140 = a11792 & ~a10920;
assign a22142 = ~a22140 & ~a22138;
assign a22144 = ~a22142 & a10962;
assign a22146 = a11800 & a10920;
assign a22148 = a11804 & ~a10920;
assign a22150 = ~a22148 & ~a22146;
assign a22152 = ~a22150 & ~a10962;
assign a22154 = ~a22152 & ~a22144;
assign a22156 = ~a22154 & ~a10816;
assign a22158 = ~a22156 & ~a22136;
assign a22160 = ~a22158 & a10876;
assign a22162 = a11820 & a10920;
assign a22164 = a11824 & ~a10920;
assign a22166 = ~a22164 & ~a22162;
assign a22168 = a10962 & a10878;
assign a22170 = a22168 & ~a22166;
assign a22174 = a22172 & ~a21872;
assign a22176 = ~a22172 & a21872;
assign a22178 = a12008 & a10920;
assign a22180 = a12016 & ~a10920;
assign a22182 = ~a22180 & ~a22178;
assign a22184 = ~a22182 & a10962;
assign a22186 = a12028 & a10920;
assign a22188 = a12036 & ~a10920;
assign a22190 = ~a22188 & ~a22186;
assign a22192 = ~a22190 & ~a10962;
assign a22194 = ~a22192 & ~a22184;
assign a22196 = ~a22194 & a10816;
assign a22198 = a12048 & a10920;
assign a22200 = a12052 & ~a10920;
assign a22202 = ~a22200 & ~a22198;
assign a22204 = ~a22202 & a10962;
assign a22206 = a12060 & a10920;
assign a22208 = a12064 & ~a10920;
assign a22210 = ~a22208 & ~a22206;
assign a22212 = ~a22210 & ~a10962;
assign a22214 = ~a22212 & ~a22204;
assign a22216 = ~a22214 & ~a10816;
assign a22218 = ~a22216 & ~a22196;
assign a22220 = ~a22218 & a10876;
assign a22222 = a12080 & a10920;
assign a22224 = a12084 & ~a10920;
assign a22226 = ~a22224 & ~a22222;
assign a22228 = ~a22226 & a22168;
assign a22232 = a22230 & ~a21888;
assign a22234 = ~a22230 & a21888;
assign a22236 = a12196 & a10920;
assign a22238 = a12204 & ~a10920;
assign a22240 = ~a22238 & ~a22236;
assign a22242 = ~a22240 & a10962;
assign a22244 = a12216 & a10920;
assign a22246 = a12224 & ~a10920;
assign a22248 = ~a22246 & ~a22244;
assign a22250 = ~a22248 & ~a10962;
assign a22252 = ~a22250 & ~a22242;
assign a22254 = ~a22252 & a10816;
assign a22256 = a12236 & a10920;
assign a22258 = a12240 & ~a10920;
assign a22260 = ~a22258 & ~a22256;
assign a22262 = ~a22260 & a10962;
assign a22264 = a12248 & a10920;
assign a22266 = a12252 & ~a10920;
assign a22268 = ~a22266 & ~a22264;
assign a22270 = ~a22268 & ~a10962;
assign a22272 = ~a22270 & ~a22262;
assign a22274 = ~a22272 & ~a10816;
assign a22276 = ~a22274 & ~a22254;
assign a22278 = ~a22276 & a10876;
assign a22280 = a12268 & a10920;
assign a22282 = a12272 & ~a10920;
assign a22284 = ~a22282 & ~a22280;
assign a22286 = ~a22284 & a22168;
assign a22290 = a22288 & ~a21904;
assign a22292 = ~a22288 & a21904;
assign a22294 = a12396 & a10920;
assign a22296 = a12404 & ~a10920;
assign a22298 = ~a22296 & ~a22294;
assign a22300 = ~a22298 & a10962;
assign a22302 = a12416 & a10920;
assign a22304 = a12424 & ~a10920;
assign a22306 = ~a22304 & ~a22302;
assign a22308 = ~a22306 & ~a10962;
assign a22310 = ~a22308 & ~a22300;
assign a22312 = ~a22310 & a10816;
assign a22314 = a12436 & a10920;
assign a22316 = a12440 & ~a10920;
assign a22318 = ~a22316 & ~a22314;
assign a22320 = ~a22318 & a10962;
assign a22322 = a12448 & a10920;
assign a22324 = a12452 & ~a10920;
assign a22326 = ~a22324 & ~a22322;
assign a22328 = ~a22326 & ~a10962;
assign a22330 = ~a22328 & ~a22320;
assign a22332 = ~a22330 & ~a10816;
assign a22334 = ~a22332 & ~a22312;
assign a22336 = ~a22334 & a10876;
assign a22338 = a12468 & a10920;
assign a22340 = a12472 & ~a10920;
assign a22342 = ~a22340 & ~a22338;
assign a22344 = ~a22342 & a22168;
assign a22348 = a22346 & ~a21920;
assign a22350 = ~a22346 & a21920;
assign a22352 = a12596 & a10920;
assign a22354 = a12604 & ~a10920;
assign a22356 = ~a22354 & ~a22352;
assign a22358 = ~a22356 & a10962;
assign a22360 = a12616 & a10920;
assign a22362 = a12624 & ~a10920;
assign a22364 = ~a22362 & ~a22360;
assign a22366 = ~a22364 & ~a10962;
assign a22368 = ~a22366 & ~a22358;
assign a22370 = ~a22368 & a10816;
assign a22372 = a12636 & a10920;
assign a22374 = a12640 & ~a10920;
assign a22376 = ~a22374 & ~a22372;
assign a22378 = ~a22376 & a10962;
assign a22380 = a12648 & a10920;
assign a22382 = a12652 & ~a10920;
assign a22384 = ~a22382 & ~a22380;
assign a22386 = ~a22384 & ~a10962;
assign a22388 = ~a22386 & ~a22378;
assign a22390 = ~a22388 & ~a10816;
assign a22392 = ~a22390 & ~a22370;
assign a22394 = ~a22392 & a10876;
assign a22396 = a12668 & a10920;
assign a22398 = a12672 & ~a10920;
assign a22400 = ~a22398 & ~a22396;
assign a22402 = ~a22400 & a22168;
assign a22406 = a22404 & ~a21936;
assign a22408 = ~a22404 & a21936;
assign a22410 = a12796 & a10920;
assign a22412 = a12804 & ~a10920;
assign a22414 = ~a22412 & ~a22410;
assign a22416 = ~a22414 & a10962;
assign a22418 = a12816 & a10920;
assign a22420 = a12824 & ~a10920;
assign a22422 = ~a22420 & ~a22418;
assign a22424 = ~a22422 & ~a10962;
assign a22426 = ~a22424 & ~a22416;
assign a22428 = ~a22426 & a10816;
assign a22430 = a12836 & a10920;
assign a22432 = a12840 & ~a10920;
assign a22434 = ~a22432 & ~a22430;
assign a22436 = ~a22434 & a10962;
assign a22438 = a12848 & a10920;
assign a22440 = a12852 & ~a10920;
assign a22442 = ~a22440 & ~a22438;
assign a22444 = ~a22442 & ~a10962;
assign a22446 = ~a22444 & ~a22436;
assign a22448 = ~a22446 & ~a10816;
assign a22450 = ~a22448 & ~a22428;
assign a22452 = ~a22450 & a10876;
assign a22454 = a12868 & a10920;
assign a22456 = a12872 & ~a10920;
assign a22458 = ~a22456 & ~a22454;
assign a22460 = ~a22458 & a22168;
assign a22464 = a22462 & ~a21952;
assign a22466 = ~a22462 & a21952;
assign a22468 = a11304 & a10920;
assign a22470 = a11316 & ~a10920;
assign a22472 = ~a22470 & ~a22468;
assign a22474 = ~a22472 & a10962;
assign a22476 = a11328 & a10920;
assign a22478 = a11336 & ~a10920;
assign a22480 = ~a22478 & ~a22476;
assign a22482 = ~a22480 & ~a10962;
assign a22484 = ~a22482 & ~a22474;
assign a22486 = ~a22484 & a10816;
assign a22488 = a11348 & a10920;
assign a22490 = a11352 & ~a10920;
assign a22492 = ~a22490 & ~a22488;
assign a22494 = ~a22492 & a10962;
assign a22496 = a11360 & a10920;
assign a22498 = a11364 & ~a10920;
assign a22500 = ~a22498 & ~a22496;
assign a22502 = ~a22500 & ~a10962;
assign a22504 = ~a22502 & ~a22494;
assign a22506 = ~a22504 & ~a10816;
assign a22508 = ~a22506 & ~a22486;
assign a22510 = ~a22508 & a10876;
assign a22512 = a11292 & a10920;
assign a22514 = a11296 & ~a10920;
assign a22516 = ~a22514 & ~a22512;
assign a22518 = ~a22516 & a22168;
assign a22522 = ~a22520 & a21968;
assign a22524 = ~a22522 & ~a22466;
assign a22526 = ~a22524 & ~a22464;
assign a22528 = ~a22526 & ~a22408;
assign a22530 = ~a22528 & ~a22406;
assign a22532 = ~a22530 & ~a22350;
assign a22534 = ~a22532 & ~a22348;
assign a22536 = ~a22534 & ~a22292;
assign a22538 = ~a22536 & ~a22290;
assign a22540 = ~a22538 & ~a22234;
assign a22542 = ~a22540 & ~a22232;
assign a22544 = ~a22542 & ~a22176;
assign a22546 = ~a22544 & ~a22174;
assign a22548 = a11214 & a10920;
assign a22550 = a11222 & ~a10920;
assign a22552 = ~a22550 & ~a22548;
assign a22554 = ~a22552 & a10962;
assign a22556 = a11230 & a10920;
assign a22558 = a11234 & ~a10920;
assign a22560 = ~a22558 & ~a22556;
assign a22562 = ~a22560 & ~a10962;
assign a22564 = ~a22562 & ~a22554;
assign a22566 = ~a22564 & a10816;
assign a22568 = a11246 & a10920;
assign a22570 = a11250 & ~a10920;
assign a22572 = ~a22570 & ~a22568;
assign a22574 = ~a22572 & a10962;
assign a22576 = a11258 & a10920;
assign a22578 = a11262 & ~a10920;
assign a22580 = ~a22578 & ~a22576;
assign a22582 = ~a22580 & ~a10962;
assign a22584 = ~a22582 & ~a22574;
assign a22586 = ~a22584 & ~a10816;
assign a22588 = ~a22586 & ~a22566;
assign a22590 = ~a22588 & a10876;
assign a22592 = a11202 & a10920;
assign a22594 = a11206 & ~a10920;
assign a22596 = ~a22594 & ~a22592;
assign a22598 = ~a22596 & a22168;
assign a22602 = ~a22600 & a22006;
assign a22604 = a22600 & ~a22006;
assign a22606 = ~a22604 & ~a22602;
assign a22608 = ~a22606 & a22546;
assign a22610 = a22606 & ~a22546;
assign a22612 = ~a22610 & ~a22608;
assign a22614 = ~a22612 & ~a22116;
assign a22616 = a22614 & ~a8032;
assign a22618 = a22616 & i418;
assign a22620 = ~a22618 & a21860;
assign a22622 = ~a22620 & a21816;
assign a22624 = a22622 & ~a8068;
assign a22626 = ~a22624 & a8032;
assign a22628 = ~a22626 & a21814;
assign a22632 = a15336 & l958;
assign a22634 = a22624 & ~a8048;
assign a22636 = ~a22634 & a15320;
assign a22640 = a15328 & l958;
assign a22642 = ~a15328 & ~l958;
assign a22644 = ~a22642 & ~a22640;
assign a22646 = ~a22644 & ~a15338;
assign a22648 = ~a15320 & a15298;
assign a22650 = a22648 & a13508;
assign a22652 = a22650 & i352;
assign a22654 = a22652 & a15338;
assign a22658 = ~a22642 & l954;
assign a22660 = a22642 & ~l954;
assign a22662 = ~a22660 & ~a22658;
assign a22666 = ~a22660 & a15332;
assign a22672 = ~a22654 & a15990;
assign a22674 = a22654 & a8868;
assign a22678 = a13508 & i438;
assign a22680 = a22678 & a15298;
assign a22682 = ~a11388 & a10778;
assign a22684 = ~a22682 & ~a22680;
assign a22690 = ~a10800 & ~a10784;
assign a22692 = ~a22690 & ~a11388;
assign a22694 = ~a22692 & ~a22680;
assign a22698 = ~a10800 & l984;
assign a22700 = a10800 & ~l984;
assign a22702 = ~a22700 & ~a22698;
assign a22704 = ~a22702 & ~a11388;
assign a22708 = ~a22700 & ~a10774;
assign a22710 = ~a22708 & ~a22680;
assign a22714 = a21816 & i464;
assign a22716 = ~i454 & ~i452;
assign a22718 = ~a22716 & i456;
assign a22720 = a22718 & i450;
assign a22722 = a22720 & i448;
assign a22724 = a22722 & i446;
assign a22726 = a22724 & i444;
assign a22728 = ~a22726 & ~i442;
assign a22730 = ~a13508 & a11432;
assign a22732 = ~a22730 & ~a13516;
assign a22734 = ~a22732 & a21814;
assign a22736 = ~a21814 & ~a15314;
assign a22738 = ~a22736 & ~a22734;
assign a22740 = ~a22738 & ~l1494;
assign a22742 = a15350 & l1494;
assign a22744 = ~a22742 & ~a22740;
assign a22746 = ~a22744 & a13494;
assign a22748 = ~a13494 & a5514;
assign a22752 = ~a22750 & a13162;
assign a22754 = a22750 & ~a13162;
assign a22756 = ~a22754 & ~a22752;
assign a22758 = ~a13508 & a11486;
assign a22760 = ~a22758 & ~a13630;
assign a22762 = ~a22760 & a21814;
assign a22764 = ~a21814 & ~a15884;
assign a22766 = ~a22764 & ~a22762;
assign a22768 = ~a22766 & ~l1494;
assign a22770 = a15892 & l1494;
assign a22772 = ~a22770 & ~a22768;
assign a22774 = ~a22772 & a13494;
assign a22776 = ~a13494 & a5396;
assign a22780 = ~a22778 & a12002;
assign a22782 = a22778 & ~a12002;
assign a22784 = ~a22782 & ~a22780;
assign a22786 = ~a13508 & a11478;
assign a22788 = ~a22786 & ~a13610;
assign a22790 = ~a22788 & a21814;
assign a22792 = ~a21814 & ~a15786;
assign a22794 = ~a22792 & ~a22790;
assign a22796 = ~a22794 & ~l1494;
assign a22798 = a15794 & l1494;
assign a22800 = ~a22798 & ~a22796;
assign a22802 = ~a22800 & a13494;
assign a22804 = ~a13494 & a5394;
assign a22808 = ~a22806 & a12190;
assign a22810 = a22806 & ~a12190;
assign a22812 = ~a22810 & ~a22808;
assign a22814 = ~a13508 & a11472;
assign a22816 = ~a22814 & ~a13590;
assign a22818 = ~a22816 & a21814;
assign a22820 = ~a21814 & ~a15682;
assign a22822 = ~a22820 & ~a22818;
assign a22824 = ~a22822 & ~l1494;
assign a22826 = a15696 & l1494;
assign a22828 = ~a22826 & ~a22824;
assign a22830 = ~a22828 & a13494;
assign a22832 = ~a13494 & a5392;
assign a22836 = ~a22834 & a12390;
assign a22838 = a22834 & ~a12390;
assign a22840 = ~a22838 & ~a22836;
assign a22842 = ~a13508 & a11462;
assign a22844 = ~a22842 & ~a13570;
assign a22846 = ~a22844 & a21814;
assign a22848 = ~a21814 & ~a15578;
assign a22850 = ~a22848 & ~a22846;
assign a22852 = ~a22850 & ~l1494;
assign a22854 = a15592 & l1494;
assign a22856 = ~a22854 & ~a22852;
assign a22858 = ~a22856 & a13494;
assign a22860 = ~a13494 & a5384;
assign a22864 = ~a22862 & a12590;
assign a22866 = a22862 & ~a12590;
assign a22868 = ~a22866 & ~a22864;
assign a22870 = ~a13508 & a11452;
assign a22872 = ~a22870 & ~a13550;
assign a22874 = ~a22872 & a21814;
assign a22876 = ~a21814 & ~a15474;
assign a22878 = ~a22876 & ~a22874;
assign a22880 = ~a22878 & ~l1494;
assign a22882 = a15488 & l1494;
assign a22884 = ~a22882 & ~a22880;
assign a22886 = ~a22884 & a13494;
assign a22888 = ~a13494 & a5376;
assign a22892 = ~a22890 & a12790;
assign a22894 = a22890 & ~a12790;
assign a22896 = ~a22894 & ~a22892;
assign a22898 = ~a13508 & a11442;
assign a22900 = ~a22898 & ~a13530;
assign a22902 = ~a22900 & a21814;
assign a22904 = ~a21814 & ~a15370;
assign a22906 = ~a22904 & ~a22902;
assign a22908 = ~a22906 & ~l1494;
assign a22910 = a15384 & l1494;
assign a22912 = ~a22910 & ~a22908;
assign a22914 = ~a22912 & a13494;
assign a22916 = ~a13494 & a5368;
assign a22920 = ~a22918 & a12990;
assign a22922 = a22918 & ~a12990;
assign a22924 = ~a22922 & ~a22920;
assign a22926 = ~a13508 & a11490;
assign a22928 = ~a22926 & ~a13650;
assign a22930 = ~a22928 & a21814;
assign a22932 = ~a21814 & ~a15982;
assign a22934 = ~a22932 & ~a22930;
assign a22936 = ~a22934 & ~l1494;
assign a22938 = a15990 & l1494;
assign a22940 = ~a22938 & ~a22936;
assign a22942 = ~a22940 & a13494;
assign a22944 = ~a13494 & a5398;
assign a22948 = ~a22946 & a13336;
assign a22950 = a22946 & ~a13336;
assign a22952 = ~a22950 & ~a22948;
assign a22954 = ~a22952 & a22756;
assign a22956 = a22954 & a22924;
assign a22958 = a22956 & a22896;
assign a22960 = a22958 & a22868;
assign a22962 = a22960 & a22840;
assign a22964 = a22962 & a22812;
assign a22966 = a22964 & a22784;
assign a22968 = i458 & i442;
assign a22970 = a22968 & i460;
assign a22972 = ~a22968 & ~i460;
assign a22974 = ~a22972 & ~a22970;
assign a22976 = a22974 & ~a22726;
assign a22978 = a22970 & i462;
assign a22980 = a22978 & i454;
assign a22982 = ~a22978 & ~i454;
assign a22984 = ~a22982 & ~a22980;
assign a22986 = ~a22984 & ~a22726;
assign a22988 = ~a22920 & ~a22752;
assign a22990 = ~a22988 & ~a22922;
assign a22992 = ~a22990 & ~a22892;
assign a22994 = ~a22992 & ~a22894;
assign a22996 = ~a22994 & ~a22864;
assign a22998 = ~a22996 & ~a22866;
assign a23000 = ~a22998 & ~a22836;
assign a23002 = ~a23000 & ~a22838;
assign a23004 = ~a23002 & ~a22808;
assign a23006 = ~a23004 & ~a22810;
assign a23008 = a23006 & a22784;
assign a23010 = ~a23006 & ~a22784;
assign a23012 = ~a23010 & ~a23008;
assign a23014 = a22980 & i452;
assign a23016 = a23014 & i456;
assign a23018 = a23016 & i450;
assign a23020 = a23018 & i448;
assign a23022 = a23020 & i446;
assign a23024 = ~a23022 & i444;
assign a23026 = a23022 & ~i444;
assign a23028 = ~a23026 & ~a23024;
assign a23030 = a23028 & ~a22726;
assign a23032 = a22924 & a22752;
assign a23034 = ~a22924 & ~a22752;
assign a23036 = ~a23034 & ~a23032;
assign a23038 = a22990 & a22896;
assign a23040 = ~a22990 & ~a22896;
assign a23042 = ~a23040 & ~a23038;
assign a23044 = a22994 & a22868;
assign a23046 = ~a22994 & ~a22868;
assign a23048 = ~a23046 & ~a23044;
assign a23050 = a22998 & a22840;
assign a23052 = ~a22998 & ~a22840;
assign a23054 = ~a23052 & ~a23050;
assign a23056 = a23002 & a22812;
assign a23058 = ~a23002 & ~a22812;
assign a23060 = ~a23058 & ~a23056;
assign a23062 = a23012 & ~a22756;
assign a23064 = a23062 & a23060;
assign a23066 = a23064 & a23054;
assign a23068 = a23066 & a23048;
assign a23070 = a23068 & a23042;
assign a23072 = a23070 & a23036;
assign a23074 = ~a23072 & ~a23030;
assign a23076 = ~a23036 & a23012;
assign a23078 = a23076 & a23060;
assign a23080 = a23078 & a23054;
assign a23082 = a23080 & a23048;
assign a23084 = a23074 & a23036;
assign a23086 = ~a23074 & ~a23036;
assign a23088 = ~a23020 & ~i446;
assign a23090 = ~a23088 & ~a23022;
assign a23092 = ~a23090 & ~a22726;
assign a23094 = a23092 & ~a22756;
assign a23096 = ~a23094 & ~a23086;
assign a23098 = ~a23096 & ~a23084;
assign a23100 = ~a23098 & a23082;
assign a23102 = a23100 & a23042;
assign a23104 = ~a23102 & a23074;
assign a23106 = ~a23042 & a23012;
assign a23108 = a23106 & a23060;
assign a23110 = a23108 & a23054;
assign a23112 = a23104 & a23042;
assign a23114 = ~a23104 & ~a23042;
assign a23116 = ~a23098 & a23070;
assign a23118 = ~a23116 & ~a23092;
assign a23120 = a23118 & a23036;
assign a23122 = ~a23118 & ~a23036;
assign a23124 = ~a23018 & ~i448;
assign a23126 = ~a23124 & ~a23020;
assign a23128 = ~a23126 & ~a22726;
assign a23130 = a23128 & ~a22756;
assign a23132 = ~a23130 & ~a23122;
assign a23134 = ~a23132 & ~a23120;
assign a23136 = ~a23134 & ~a23114;
assign a23138 = ~a23136 & ~a23112;
assign a23140 = ~a23138 & a23110;
assign a23142 = a23140 & a23048;
assign a23144 = ~a23138 & a23082;
assign a23146 = a23144 & ~a23118;
assign a23148 = ~a23146 & ~a23142;
assign a23150 = a23148 & a23104;
assign a23152 = ~a23138 & a23068;
assign a23154 = a23152 & a23128;
assign a23156 = ~a23152 & ~a23128;
assign a23158 = ~a23156 & ~a23154;
assign a23160 = a23150 & a23048;
assign a23162 = ~a23150 & ~a23048;
assign a23164 = ~a23144 & a23118;
assign a23166 = ~a23164 & ~a23146;
assign a23168 = ~a23166 & ~a23154;
assign a23170 = a23168 & a23042;
assign a23172 = ~a23168 & ~a23042;
assign a23174 = ~a23158 & a23036;
assign a23176 = a23158 & ~a23036;
assign a23178 = ~a23016 & ~i450;
assign a23180 = ~a23178 & ~a23018;
assign a23182 = ~a23180 & ~a22726;
assign a23184 = a23182 & ~a22756;
assign a23186 = ~a23184 & ~a23176;
assign a23188 = ~a23186 & ~a23174;
assign a23190 = ~a23188 & ~a23172;
assign a23192 = ~a23190 & ~a23170;
assign a23194 = ~a23192 & ~a23162;
assign a23196 = ~a23194 & ~a23160;
assign a23198 = ~a23196 & a23080;
assign a23200 = a23198 & a23158;
assign a23202 = ~a23196 & a23066;
assign a23204 = a23202 & a23182;
assign a23206 = ~a23204 & ~a23200;
assign a23208 = ~a23198 & ~a23158;
assign a23210 = ~a23208 & ~a23206;
assign a23212 = ~a23196 & a23110;
assign a23214 = a23212 & ~a23168;
assign a23216 = ~a23214 & ~a23210;
assign a23218 = ~a23212 & a23168;
assign a23220 = ~a23218 & ~a23216;
assign a23222 = ~a23048 & a23012;
assign a23224 = a23222 & a23060;
assign a23226 = a23224 & ~a23196;
assign a23228 = a23226 & a23054;
assign a23230 = ~a23228 & ~a23220;
assign a23232 = a23230 & a23150;
assign a23234 = ~a23202 & ~a23182;
assign a23236 = ~a23234 & ~a23204;
assign a23238 = a23232 & a23054;
assign a23240 = ~a23232 & ~a23054;
assign a23242 = ~a23218 & ~a23214;
assign a23244 = a23242 & a23210;
assign a23246 = ~a23242 & ~a23210;
assign a23248 = ~a23246 & ~a23244;
assign a23250 = ~a23248 & a23048;
assign a23252 = a23248 & ~a23048;
assign a23254 = ~a23208 & ~a23200;
assign a23256 = a23254 & a23204;
assign a23258 = ~a23254 & ~a23204;
assign a23260 = ~a23258 & ~a23256;
assign a23262 = ~a23260 & a23042;
assign a23264 = a23260 & ~a23042;
assign a23266 = ~a23236 & a23036;
assign a23268 = a23236 & ~a23036;
assign a23270 = ~a23014 & ~i456;
assign a23272 = ~a23270 & ~a23016;
assign a23274 = ~a23272 & ~a22726;
assign a23276 = a23274 & ~a22756;
assign a23278 = ~a23276 & ~a23268;
assign a23280 = ~a23278 & ~a23266;
assign a23282 = ~a23280 & ~a23264;
assign a23284 = ~a23282 & ~a23262;
assign a23286 = ~a23284 & ~a23252;
assign a23288 = ~a23286 & ~a23250;
assign a23290 = ~a23288 & ~a23240;
assign a23292 = ~a23290 & ~a23238;
assign a23294 = ~a23292 & a23078;
assign a23296 = a23294 & a23236;
assign a23298 = ~a23292 & a23064;
assign a23300 = a23298 & a23274;
assign a23302 = ~a23300 & ~a23296;
assign a23304 = ~a23294 & ~a23236;
assign a23306 = ~a23304 & ~a23302;
assign a23308 = ~a23292 & a23108;
assign a23310 = a23308 & a23260;
assign a23312 = ~a23310 & ~a23306;
assign a23314 = ~a23308 & ~a23260;
assign a23316 = ~a23314 & ~a23312;
assign a23318 = ~a23292 & a23224;
assign a23320 = a23318 & a23248;
assign a23322 = ~a23320 & ~a23316;
assign a23324 = ~a23318 & ~a23248;
assign a23326 = ~a23324 & ~a23322;
assign a23328 = ~a23054 & a23012;
assign a23330 = a23328 & ~a23292;
assign a23332 = a23330 & a23060;
assign a23334 = ~a23332 & ~a23326;
assign a23336 = a23334 & a23232;
assign a23338 = ~a23298 & ~a23274;
assign a23340 = ~a23338 & ~a23300;
assign a23342 = a23336 & a23060;
assign a23344 = ~a23336 & ~a23060;
assign a23346 = ~a23324 & ~a23320;
assign a23348 = a23346 & a23316;
assign a23350 = ~a23346 & ~a23316;
assign a23352 = ~a23350 & ~a23348;
assign a23354 = ~a23352 & a23054;
assign a23356 = a23352 & ~a23054;
assign a23358 = ~a23314 & ~a23310;
assign a23360 = a23358 & a23306;
assign a23362 = ~a23358 & ~a23306;
assign a23364 = ~a23362 & ~a23360;
assign a23366 = ~a23364 & a23048;
assign a23368 = a23364 & ~a23048;
assign a23370 = ~a23304 & ~a23296;
assign a23372 = a23370 & a23300;
assign a23374 = ~a23370 & ~a23300;
assign a23376 = ~a23374 & ~a23372;
assign a23378 = ~a23376 & a23042;
assign a23380 = a23376 & ~a23042;
assign a23382 = ~a23340 & a23036;
assign a23384 = a23340 & ~a23036;
assign a23386 = ~a22980 & ~i452;
assign a23388 = ~a23386 & ~a23014;
assign a23390 = a23388 & ~a22726;
assign a23392 = ~a23390 & ~a22756;
assign a23394 = ~a23392 & ~a23384;
assign a23396 = ~a23394 & ~a23382;
assign a23398 = ~a23396 & ~a23380;
assign a23400 = ~a23398 & ~a23378;
assign a23402 = ~a23400 & ~a23368;
assign a23404 = ~a23402 & ~a23366;
assign a23406 = ~a23404 & ~a23356;
assign a23408 = ~a23406 & ~a23354;
assign a23410 = ~a23408 & ~a23344;
assign a23412 = ~a23410 & ~a23342;
assign a23414 = ~a23412 & a23076;
assign a23416 = a23414 & a23340;
assign a23418 = ~a23412 & a23062;
assign a23420 = a23418 & ~a23390;
assign a23422 = ~a23420 & ~a23416;
assign a23424 = ~a23414 & ~a23340;
assign a23426 = ~a23424 & ~a23422;
assign a23428 = ~a23412 & a23106;
assign a23430 = a23428 & a23376;
assign a23432 = ~a23430 & ~a23426;
assign a23434 = ~a23428 & ~a23376;
assign a23436 = ~a23434 & ~a23432;
assign a23438 = ~a23412 & a23222;
assign a23440 = a23438 & a23364;
assign a23442 = ~a23440 & ~a23436;
assign a23444 = ~a23438 & ~a23364;
assign a23446 = ~a23444 & ~a23442;
assign a23448 = ~a23412 & a23328;
assign a23450 = a23448 & a23352;
assign a23452 = ~a23450 & ~a23446;
assign a23454 = ~a23448 & ~a23352;
assign a23456 = ~a23454 & ~a23452;
assign a23458 = ~a23412 & ~a23060;
assign a23460 = a23458 & a23012;
assign a23462 = ~a23460 & ~a23456;
assign a23464 = a23462 & a23336;
assign a23466 = a23464 & a23012;
assign a23468 = ~a23464 & ~a23012;
assign a23470 = ~a23454 & ~a23450;
assign a23472 = a23470 & a23446;
assign a23474 = ~a23470 & ~a23446;
assign a23476 = ~a23474 & ~a23472;
assign a23478 = ~a23476 & a23060;
assign a23480 = a23476 & ~a23060;
assign a23482 = ~a23444 & ~a23440;
assign a23484 = a23482 & a23436;
assign a23486 = ~a23482 & ~a23436;
assign a23488 = ~a23486 & ~a23484;
assign a23490 = ~a23488 & a23054;
assign a23492 = a23488 & ~a23054;
assign a23494 = ~a23434 & ~a23430;
assign a23496 = a23494 & a23426;
assign a23498 = ~a23494 & ~a23426;
assign a23500 = ~a23498 & ~a23496;
assign a23502 = ~a23500 & a23048;
assign a23504 = a23500 & ~a23048;
assign a23506 = ~a23424 & ~a23416;
assign a23508 = a23506 & a23420;
assign a23510 = ~a23506 & ~a23420;
assign a23512 = ~a23510 & ~a23508;
assign a23514 = ~a23512 & a23042;
assign a23516 = a23512 & ~a23042;
assign a23518 = ~a23418 & a23390;
assign a23520 = ~a23518 & ~a23420;
assign a23522 = ~a23520 & a23036;
assign a23524 = a23520 & ~a23036;
assign a23526 = a22986 & ~a22756;
assign a23528 = ~a23526 & ~a23524;
assign a23530 = ~a23528 & ~a23522;
assign a23532 = ~a23530 & ~a23516;
assign a23534 = ~a23532 & ~a23514;
assign a23536 = ~a23534 & ~a23504;
assign a23538 = ~a23536 & ~a23502;
assign a23540 = ~a23538 & ~a23492;
assign a23542 = ~a23540 & ~a23490;
assign a23544 = ~a23542 & ~a23480;
assign a23546 = ~a23544 & ~a23478;
assign a23548 = ~a23546 & ~a23468;
assign a23550 = ~a23548 & ~a23466;
assign a23552 = ~a23550 & ~a22756;
assign a23554 = a23552 & a22986;
assign a23556 = ~a23552 & ~a22986;
assign a23558 = ~a23556 & ~a23554;
assign a23560 = ~a23550 & ~a23036;
assign a23562 = a23560 & a23520;
assign a23564 = ~a23562 & ~a23554;
assign a23566 = ~a23560 & ~a23520;
assign a23568 = ~a23566 & ~a23564;
assign a23570 = ~a23550 & ~a23042;
assign a23572 = a23570 & a23512;
assign a23574 = ~a23572 & ~a23568;
assign a23576 = ~a23570 & ~a23512;
assign a23578 = ~a23576 & ~a23574;
assign a23580 = ~a23550 & ~a23048;
assign a23582 = a23580 & a23500;
assign a23584 = ~a23582 & ~a23578;
assign a23586 = ~a23580 & ~a23500;
assign a23588 = ~a23586 & ~a23584;
assign a23590 = ~a23550 & ~a23054;
assign a23592 = a23590 & a23488;
assign a23594 = ~a23592 & ~a23588;
assign a23596 = ~a23590 & ~a23488;
assign a23598 = ~a23596 & ~a23594;
assign a23600 = ~a23550 & ~a23060;
assign a23602 = a23600 & a23476;
assign a23604 = ~a23602 & ~a23598;
assign a23606 = ~a23600 & ~a23476;
assign a23608 = ~a23606 & ~a23604;
assign a23610 = ~a23550 & ~a23012;
assign a23612 = ~a23610 & ~a23608;
assign a23614 = a23612 & a23464;
assign a23616 = a23614 & ~a22966;
assign a23618 = ~a23614 & a22966;
assign a23620 = ~a23606 & ~a23602;
assign a23622 = a23620 & a23598;
assign a23624 = ~a23620 & ~a23598;
assign a23626 = ~a23624 & ~a23622;
assign a23628 = ~a23626 & a23012;
assign a23630 = a23626 & ~a23012;
assign a23632 = ~a23596 & ~a23592;
assign a23634 = a23632 & a23588;
assign a23636 = ~a23632 & ~a23588;
assign a23638 = ~a23636 & ~a23634;
assign a23640 = ~a23638 & a23060;
assign a23642 = a23638 & ~a23060;
assign a23644 = ~a23586 & ~a23582;
assign a23646 = a23644 & a23578;
assign a23648 = ~a23644 & ~a23578;
assign a23650 = ~a23648 & ~a23646;
assign a23652 = ~a23650 & a23054;
assign a23654 = a23650 & ~a23054;
assign a23656 = ~a23576 & ~a23572;
assign a23658 = a23656 & a23568;
assign a23660 = ~a23656 & ~a23568;
assign a23662 = ~a23660 & ~a23658;
assign a23664 = ~a23662 & a23048;
assign a23666 = a23662 & ~a23048;
assign a23668 = ~a23566 & ~a23562;
assign a23670 = a23668 & a23554;
assign a23672 = ~a23668 & ~a23554;
assign a23674 = ~a23672 & ~a23670;
assign a23676 = ~a23674 & a23042;
assign a23678 = a23674 & ~a23042;
assign a23680 = ~a23558 & a23036;
assign a23682 = a23558 & ~a23036;
assign a23684 = ~a22970 & ~i462;
assign a23686 = ~a23684 & ~a22978;
assign a23688 = a23686 & ~a22726;
assign a23690 = ~a23688 & ~a22756;
assign a23692 = ~a23690 & ~a23682;
assign a23694 = ~a23692 & ~a23680;
assign a23696 = ~a23694 & ~a23678;
assign a23698 = ~a23696 & ~a23676;
assign a23700 = ~a23698 & ~a23666;
assign a23702 = ~a23700 & ~a23664;
assign a23704 = ~a23702 & ~a23654;
assign a23706 = ~a23704 & ~a23652;
assign a23708 = ~a23706 & ~a23642;
assign a23710 = ~a23708 & ~a23640;
assign a23712 = ~a23710 & ~a23630;
assign a23714 = ~a23712 & ~a23628;
assign a23716 = ~a23714 & ~a23618;
assign a23718 = ~a23716 & ~a23616;
assign a23720 = ~a23718 & ~a23036;
assign a23722 = a23720 & a23558;
assign a23724 = ~a23718 & ~a22756;
assign a23726 = a23724 & ~a23688;
assign a23728 = ~a23726 & ~a23722;
assign a23730 = ~a23720 & ~a23558;
assign a23732 = ~a23730 & ~a23728;
assign a23734 = ~a23718 & ~a23042;
assign a23736 = a23734 & a23674;
assign a23738 = ~a23736 & ~a23732;
assign a23740 = ~a23734 & ~a23674;
assign a23742 = ~a23740 & ~a23738;
assign a23744 = ~a23718 & ~a23048;
assign a23746 = a23744 & a23662;
assign a23748 = ~a23746 & ~a23742;
assign a23750 = ~a23744 & ~a23662;
assign a23752 = ~a23750 & ~a23748;
assign a23754 = ~a23718 & ~a23054;
assign a23756 = a23754 & a23650;
assign a23758 = ~a23756 & ~a23752;
assign a23760 = ~a23754 & ~a23650;
assign a23762 = ~a23760 & ~a23758;
assign a23764 = ~a23718 & ~a23060;
assign a23766 = a23764 & a23638;
assign a23768 = ~a23766 & ~a23762;
assign a23770 = ~a23764 & ~a23638;
assign a23772 = ~a23770 & ~a23768;
assign a23774 = ~a23718 & ~a23012;
assign a23776 = a23774 & a23626;
assign a23778 = ~a23774 & ~a23626;
assign a23780 = ~a23778 & ~a23776;
assign a23782 = a23780 & a23772;
assign a23784 = ~a23780 & ~a23772;
assign a23786 = ~a23784 & ~a23782;
assign a23788 = ~a23786 & ~a22966;
assign a23790 = a23786 & a22966;
assign a23792 = ~a23770 & ~a23766;
assign a23794 = a23792 & a23762;
assign a23796 = ~a23792 & ~a23762;
assign a23798 = ~a23796 & ~a23794;
assign a23800 = ~a23798 & a23012;
assign a23802 = a23798 & ~a23012;
assign a23804 = ~a23760 & ~a23756;
assign a23806 = a23804 & a23752;
assign a23808 = ~a23804 & ~a23752;
assign a23810 = ~a23808 & ~a23806;
assign a23812 = ~a23810 & a23060;
assign a23814 = a23810 & ~a23060;
assign a23816 = ~a23750 & ~a23746;
assign a23818 = a23816 & a23742;
assign a23820 = ~a23816 & ~a23742;
assign a23822 = ~a23820 & ~a23818;
assign a23824 = ~a23822 & a23054;
assign a23826 = a23822 & ~a23054;
assign a23828 = ~a23740 & ~a23736;
assign a23830 = a23828 & a23732;
assign a23832 = ~a23828 & ~a23732;
assign a23834 = ~a23832 & ~a23830;
assign a23836 = ~a23834 & a23048;
assign a23838 = a23834 & ~a23048;
assign a23840 = ~a23730 & ~a23722;
assign a23842 = a23840 & a23726;
assign a23844 = ~a23840 & ~a23726;
assign a23846 = ~a23844 & ~a23842;
assign a23848 = ~a23846 & a23042;
assign a23850 = a23846 & ~a23042;
assign a23852 = ~a23724 & a23688;
assign a23854 = ~a23852 & ~a23726;
assign a23856 = ~a23854 & a23036;
assign a23858 = a23854 & ~a23036;
assign a23860 = ~a22976 & ~a22756;
assign a23862 = ~a23860 & ~a23858;
assign a23864 = ~a23862 & ~a23856;
assign a23866 = ~a23864 & ~a23850;
assign a23868 = ~a23866 & ~a23848;
assign a23870 = ~a23868 & ~a23838;
assign a23872 = ~a23870 & ~a23836;
assign a23874 = ~a23872 & ~a23826;
assign a23876 = ~a23874 & ~a23824;
assign a23878 = ~a23876 & ~a23814;
assign a23880 = ~a23878 & ~a23812;
assign a23882 = ~a23880 & ~a23802;
assign a23884 = ~a23882 & ~a23800;
assign a23886 = ~a23884 & ~a23790;
assign a23888 = ~a23886 & ~a23788;
assign a23890 = ~a23888 & ~a22756;
assign a23892 = a23890 & ~a22976;
assign a23894 = ~a23890 & a22976;
assign a23896 = ~a23894 & ~a23892;
assign a23898 = ~a23888 & ~a23036;
assign a23900 = a23898 & a23854;
assign a23902 = ~a23900 & ~a23892;
assign a23904 = ~a23898 & ~a23854;
assign a23906 = ~a23904 & ~a23902;
assign a23908 = ~a23888 & ~a23042;
assign a23910 = a23908 & a23846;
assign a23912 = ~a23910 & ~a23906;
assign a23914 = ~a23908 & ~a23846;
assign a23916 = ~a23914 & ~a23912;
assign a23918 = ~a23888 & ~a23048;
assign a23920 = a23918 & a23834;
assign a23922 = ~a23920 & ~a23916;
assign a23924 = ~a23918 & ~a23834;
assign a23926 = ~a23924 & ~a23922;
assign a23928 = ~a23888 & ~a23054;
assign a23930 = a23928 & a23822;
assign a23932 = ~a23930 & ~a23926;
assign a23934 = ~a23928 & ~a23822;
assign a23936 = ~a23934 & ~a23932;
assign a23938 = ~a23888 & ~a23060;
assign a23940 = a23938 & a23810;
assign a23942 = ~a23940 & ~a23936;
assign a23944 = ~a23938 & ~a23810;
assign a23946 = ~a23944 & ~a23942;
assign a23948 = ~a23888 & ~a23012;
assign a23950 = a23948 & a23798;
assign a23952 = ~a23948 & ~a23798;
assign a23954 = ~a23952 & ~a23950;
assign a23956 = a23954 & a23946;
assign a23958 = ~a23954 & ~a23946;
assign a23960 = ~a23958 & ~a23956;
assign a23962 = ~a23960 & ~a22966;
assign a23964 = a23960 & a22966;
assign a23966 = ~a23944 & ~a23940;
assign a23968 = a23966 & a23936;
assign a23970 = ~a23966 & ~a23936;
assign a23972 = ~a23970 & ~a23968;
assign a23974 = ~a23972 & a23012;
assign a23976 = a23972 & ~a23012;
assign a23978 = ~a23934 & ~a23930;
assign a23980 = a23978 & a23926;
assign a23982 = ~a23978 & ~a23926;
assign a23984 = ~a23982 & ~a23980;
assign a23986 = ~a23984 & a23060;
assign a23988 = a23984 & ~a23060;
assign a23990 = ~a23924 & ~a23920;
assign a23992 = a23990 & a23916;
assign a23994 = ~a23990 & ~a23916;
assign a23996 = ~a23994 & ~a23992;
assign a23998 = ~a23996 & a23054;
assign a24000 = a23996 & ~a23054;
assign a24002 = ~a23914 & ~a23910;
assign a24004 = a24002 & a23906;
assign a24006 = ~a24002 & ~a23906;
assign a24008 = ~a24006 & ~a24004;
assign a24010 = ~a24008 & a23048;
assign a24012 = a24008 & ~a23048;
assign a24014 = ~a23904 & ~a23900;
assign a24016 = a24014 & a23892;
assign a24018 = ~a24014 & ~a23892;
assign a24020 = ~a24018 & ~a24016;
assign a24022 = ~a24020 & a23042;
assign a24024 = a24020 & ~a23042;
assign a24026 = ~a23896 & a23036;
assign a24028 = a23896 & ~a23036;
assign a24030 = ~i458 & ~i442;
assign a24032 = ~a24030 & ~a22968;
assign a24034 = a24032 & ~a22726;
assign a24036 = ~a24034 & ~a22756;
assign a24038 = ~a24036 & ~a24028;
assign a24040 = ~a24038 & ~a24026;
assign a24042 = ~a24040 & ~a24024;
assign a24044 = ~a24042 & ~a24022;
assign a24046 = ~a24044 & ~a24012;
assign a24048 = ~a24046 & ~a24010;
assign a24050 = ~a24048 & ~a24000;
assign a24052 = ~a24050 & ~a23998;
assign a24054 = ~a24052 & ~a23988;
assign a24056 = ~a24054 & ~a23986;
assign a24058 = ~a24056 & ~a23976;
assign a24060 = ~a24058 & ~a23974;
assign a24062 = ~a24060 & ~a23964;
assign a24064 = ~a24062 & ~a23962;
assign a24066 = ~a24064 & ~a23036;
assign a24068 = a24066 & a23896;
assign a24070 = ~a24064 & ~a22756;
assign a24072 = a24070 & ~a24034;
assign a24074 = ~a24072 & ~a24068;
assign a24076 = ~a24066 & ~a23896;
assign a24078 = ~a24076 & ~a24074;
assign a24080 = ~a24064 & ~a23042;
assign a24082 = a24080 & a24020;
assign a24084 = ~a24082 & ~a24078;
assign a24086 = ~a24080 & ~a24020;
assign a24088 = ~a24086 & ~a24084;
assign a24090 = ~a24064 & ~a23048;
assign a24092 = a24090 & a24008;
assign a24094 = ~a24092 & ~a24088;
assign a24096 = ~a24090 & ~a24008;
assign a24098 = ~a24096 & ~a24094;
assign a24100 = ~a24064 & ~a23054;
assign a24102 = a24100 & a23996;
assign a24104 = ~a24102 & ~a24098;
assign a24106 = ~a24100 & ~a23996;
assign a24108 = ~a24106 & ~a24104;
assign a24110 = ~a24064 & ~a23060;
assign a24112 = a24110 & a23984;
assign a24114 = ~a24112 & ~a24108;
assign a24116 = ~a24110 & ~a23984;
assign a24118 = ~a24116 & ~a24114;
assign a24120 = ~a24064 & ~a23012;
assign a24122 = a24120 & a23972;
assign a24124 = ~a24120 & ~a23972;
assign a24126 = ~a24124 & ~a24122;
assign a24128 = a24126 & a24118;
assign a24130 = ~a24126 & ~a24118;
assign a24132 = ~a24130 & ~a24128;
assign a24134 = ~a24132 & ~a22966;
assign a24136 = a24132 & a22966;
assign a24138 = ~a24116 & ~a24112;
assign a24140 = a24138 & a24108;
assign a24142 = ~a24138 & ~a24108;
assign a24144 = ~a24142 & ~a24140;
assign a24146 = ~a24144 & a23012;
assign a24148 = a24144 & ~a23012;
assign a24150 = ~a24106 & ~a24102;
assign a24152 = a24150 & a24098;
assign a24154 = ~a24150 & ~a24098;
assign a24156 = ~a24154 & ~a24152;
assign a24158 = ~a24156 & a23060;
assign a24160 = a24156 & ~a23060;
assign a24162 = ~a24096 & ~a24092;
assign a24164 = a24162 & a24088;
assign a24166 = ~a24162 & ~a24088;
assign a24168 = ~a24166 & ~a24164;
assign a24170 = ~a24168 & a23054;
assign a24172 = a24168 & ~a23054;
assign a24174 = ~a24086 & ~a24082;
assign a24176 = a24174 & a24078;
assign a24178 = ~a24174 & ~a24078;
assign a24180 = ~a24178 & ~a24176;
assign a24182 = ~a24180 & a23048;
assign a24184 = a24180 & ~a23048;
assign a24186 = ~a24076 & ~a24068;
assign a24188 = a24186 & a24072;
assign a24190 = ~a24186 & ~a24072;
assign a24192 = ~a24190 & ~a24188;
assign a24194 = ~a24192 & a23042;
assign a24196 = a24192 & ~a23042;
assign a24198 = ~a24070 & a24034;
assign a24200 = ~a24198 & ~a24072;
assign a24202 = ~a24200 & a23036;
assign a24204 = a24200 & ~a23036;
assign a24206 = ~a22756 & ~a22728;
assign a24208 = ~a24206 & ~a24204;
assign a24210 = ~a24208 & ~a24202;
assign a24212 = ~a24210 & ~a24196;
assign a24214 = ~a24212 & ~a24194;
assign a24216 = ~a24214 & ~a24184;
assign a24218 = ~a24216 & ~a24182;
assign a24220 = ~a24218 & ~a24172;
assign a24222 = ~a24220 & ~a24170;
assign a24224 = ~a24222 & ~a24160;
assign a24226 = ~a24224 & ~a24158;
assign a24228 = ~a24226 & ~a24148;
assign a24230 = ~a24228 & ~a24146;
assign a24232 = ~a24230 & ~a24136;
assign a24234 = ~a24232 & ~a24134;
assign a24236 = ~a24234 & ~a22756;
assign a24238 = a24236 & ~a22728;
assign a24240 = ~a24236 & a22728;
assign a24242 = ~a24240 & ~a24238;
assign a24244 = ~a22966 & a22756;
assign a24246 = a24244 & a23036;
assign a24248 = a24246 & a23042;
assign a24250 = a24248 & a23048;
assign a24252 = a24250 & a23054;
assign a24254 = a24252 & a23060;
assign a24256 = a24254 & a23012;
assign a24258 = ~a24256 & a24242;
assign a24260 = ~a24258 & a11426;
assign a24262 = ~a24234 & ~a23036;
assign a24264 = a24262 & a24200;
assign a24266 = ~a24262 & ~a24200;
assign a24268 = ~a24266 & ~a24264;
assign a24270 = a24268 & a24238;
assign a24272 = ~a24268 & ~a24238;
assign a24274 = ~a24272 & ~a24270;
assign a24276 = a24274 & a24242;
assign a24278 = ~a24274 & ~a24242;
assign a24280 = ~a24278 & ~a24276;
assign a24282 = a24280 & ~a24256;
assign a24284 = ~a24282 & a24260;
assign a24286 = ~a24264 & ~a24238;
assign a24288 = ~a24286 & ~a24266;
assign a24290 = ~a24234 & ~a23042;
assign a24292 = a24290 & a24192;
assign a24294 = ~a24290 & ~a24192;
assign a24296 = ~a24294 & ~a24292;
assign a24298 = a24296 & a24288;
assign a24300 = ~a24296 & ~a24288;
assign a24302 = ~a24300 & ~a24298;
assign a24304 = a24302 & ~a24278;
assign a24306 = ~a24302 & a24278;
assign a24308 = ~a24306 & ~a24304;
assign a24310 = a24308 & ~a24256;
assign a24312 = ~a24310 & a24284;
assign a24314 = ~a24292 & ~a24288;
assign a24316 = ~a24314 & ~a24294;
assign a24318 = ~a24234 & ~a23048;
assign a24320 = a24318 & a24180;
assign a24322 = ~a24318 & ~a24180;
assign a24324 = ~a24322 & ~a24320;
assign a24326 = a24324 & a24316;
assign a24328 = ~a24324 & ~a24316;
assign a24330 = ~a24328 & ~a24326;
assign a24332 = a24330 & ~a24306;
assign a24334 = ~a24330 & a24306;
assign a24336 = ~a24334 & ~a24332;
assign a24338 = a24336 & ~a24256;
assign a24340 = ~a24338 & a24312;
assign a24342 = ~a24320 & ~a24316;
assign a24344 = ~a24342 & ~a24322;
assign a24346 = ~a24234 & ~a23054;
assign a24348 = a24346 & a24168;
assign a24350 = ~a24346 & ~a24168;
assign a24352 = ~a24350 & ~a24348;
assign a24354 = a24352 & a24344;
assign a24356 = ~a24352 & ~a24344;
assign a24358 = ~a24356 & ~a24354;
assign a24360 = a24358 & ~a24334;
assign a24362 = ~a24358 & a24334;
assign a24364 = ~a24362 & ~a24360;
assign a24366 = a24364 & ~a24256;
assign a24368 = ~a24366 & a24340;
assign a24370 = ~a24348 & ~a24344;
assign a24372 = ~a24370 & ~a24350;
assign a24374 = ~a24234 & ~a23060;
assign a24376 = a24374 & a24156;
assign a24378 = ~a24374 & ~a24156;
assign a24380 = ~a24378 & ~a24376;
assign a24382 = a24380 & a24372;
assign a24384 = ~a24380 & ~a24372;
assign a24386 = ~a24384 & ~a24382;
assign a24388 = a24386 & ~a24362;
assign a24390 = ~a24386 & a24362;
assign a24392 = ~a24390 & ~a24388;
assign a24394 = a24392 & ~a24256;
assign a24396 = ~a24394 & a24368;
assign a24398 = ~a24376 & ~a24372;
assign a24400 = ~a24398 & ~a24378;
assign a24402 = ~a24234 & ~a23012;
assign a24404 = a24402 & a24144;
assign a24406 = ~a24402 & ~a24144;
assign a24408 = ~a24406 & ~a24404;
assign a24410 = a24408 & a24400;
assign a24412 = ~a24408 & ~a24400;
assign a24414 = ~a24412 & ~a24410;
assign a24416 = a24414 & ~a24390;
assign a24418 = ~a24414 & a24390;
assign a24420 = ~a24418 & ~a24416;
assign a24422 = a24420 & ~a24256;
assign a24424 = ~a24422 & a24396;
assign a24426 = ~a24404 & ~a24400;
assign a24428 = ~a24426 & ~a24406;
assign a24430 = ~a24428 & a24134;
assign a24432 = ~a24430 & a24418;
assign a24434 = a24430 & ~a24418;
assign a24436 = ~a24434 & ~a24432;
assign a24438 = ~a24436 & ~a24256;
assign a24440 = ~a24438 & a24424;
assign a24444 = a24422 & a8874;
assign a24446 = a24394 & a10044;
assign a24448 = a24366 & a10074;
assign a24450 = a24338 & a10100;
assign a24452 = a24310 & a10126;
assign a24454 = a24282 & a10152;
assign a24456 = a24258 & a10178;
assign a24458 = ~a24456 & ~a24454;
assign a24460 = ~a24282 & ~a10152;
assign a24462 = ~a24460 & ~a24458;
assign a24464 = ~a24462 & ~a24452;
assign a24466 = ~a24310 & ~a10126;
assign a24468 = ~a24466 & ~a24464;
assign a24470 = ~a24468 & ~a24450;
assign a24472 = ~a24338 & ~a10100;
assign a24474 = ~a24472 & ~a24470;
assign a24476 = ~a24474 & ~a24448;
assign a24478 = ~a24366 & ~a10074;
assign a24480 = ~a24478 & ~a24476;
assign a24482 = ~a24480 & ~a24446;
assign a24484 = ~a24394 & ~a10044;
assign a24486 = ~a24484 & ~a24482;
assign a24488 = ~a24486 & ~a24444;
assign a24490 = ~a24422 & ~a8874;
assign a24492 = ~a24490 & ~a24488;
assign a24494 = ~a24492 & ~a24438;
assign a24496 = a24492 & a24438;
assign a24498 = ~a24496 & ~a24494;
assign a24500 = a24498 & a13508;
assign a24502 = ~a24500 & a8868;
assign a24504 = a24500 & ~a8868;
assign a24506 = ~a24504 & ~a24502;
assign a24508 = l1686 & ~l1492;
assign a24510 = a10782 & a10776;
assign a24512 = a24510 & a11386;
assign a24514 = ~a24512 & ~a11524;
assign a24516 = a24514 & ~a8032;
assign a24518 = a24516 & ~a24508;
assign a24520 = a24518 & ~a24506;
assign a24522 = a24422 & a11486;
assign a24524 = a24394 & a11478;
assign a24526 = a24366 & a11472;
assign a24528 = a24338 & a11462;
assign a24530 = a24310 & a11452;
assign a24532 = a24282 & a11442;
assign a24534 = a24258 & a11432;
assign a24536 = ~a24534 & ~a24532;
assign a24538 = ~a24282 & ~a11442;
assign a24540 = ~a24538 & ~a24536;
assign a24542 = ~a24540 & ~a24530;
assign a24544 = ~a24310 & ~a11452;
assign a24546 = ~a24544 & ~a24542;
assign a24548 = ~a24546 & ~a24528;
assign a24550 = ~a24338 & ~a11462;
assign a24552 = ~a24550 & ~a24548;
assign a24554 = ~a24552 & ~a24526;
assign a24556 = ~a24366 & ~a11472;
assign a24558 = ~a24556 & ~a24554;
assign a24560 = ~a24558 & ~a24524;
assign a24562 = ~a24394 & ~a11478;
assign a24564 = ~a24562 & ~a24560;
assign a24566 = ~a24564 & ~a24522;
assign a24568 = ~a24422 & ~a11486;
assign a24570 = ~a24568 & ~a24566;
assign a24572 = a24438 & ~a11490;
assign a24574 = ~a24438 & a11490;
assign a24576 = ~a24574 & ~a24572;
assign a24578 = a24576 & a24570;
assign a24580 = ~a24576 & ~a24570;
assign a24582 = ~a24580 & ~a24578;
assign a24584 = ~a24582 & ~a24518;
assign a24586 = ~a24584 & ~a24520;
assign a24588 = ~a24586 & ~l1494;
assign a24590 = a24422 & a15892;
assign a24592 = a24394 & a15794;
assign a24594 = a24366 & a15696;
assign a24596 = a24338 & a15592;
assign a24598 = a24310 & a15488;
assign a24600 = a24282 & a15384;
assign a24602 = a24258 & a15350;
assign a24604 = ~a24602 & ~a24600;
assign a24606 = ~a24282 & ~a15384;
assign a24608 = ~a24606 & ~a24604;
assign a24610 = ~a24608 & ~a24598;
assign a24612 = ~a24310 & ~a15488;
assign a24614 = ~a24612 & ~a24610;
assign a24616 = ~a24614 & ~a24596;
assign a24618 = ~a24338 & ~a15592;
assign a24620 = ~a24618 & ~a24616;
assign a24622 = ~a24620 & ~a24594;
assign a24624 = ~a24366 & ~a15696;
assign a24626 = ~a24624 & ~a24622;
assign a24628 = ~a24626 & ~a24592;
assign a24630 = ~a24394 & ~a15794;
assign a24632 = ~a24630 & ~a24628;
assign a24634 = ~a24632 & ~a24590;
assign a24636 = ~a24422 & ~a15892;
assign a24638 = ~a24636 & ~a24634;
assign a24640 = a24438 & ~a15990;
assign a24642 = ~a24438 & a15990;
assign a24644 = ~a24642 & ~a24640;
assign a24646 = a24644 & a24638;
assign a24648 = ~a24644 & ~a24638;
assign a24650 = ~a24648 & ~a24646;
assign a24652 = ~a24650 & l1494;
assign a24654 = ~a24652 & ~a24588;
assign a24656 = ~a24654 & a13494;
assign a24658 = ~a13494 & a11490;
assign a24662 = ~a12186 & i378;
assign a24664 = i380 & ~i378;
assign a24666 = a24664 & i376;
assign a24668 = a24666 & i374;
assign a24670 = a24668 & i372;
assign a24672 = ~a24670 & i370;
assign a24674 = ~a24672 & ~a13158;
assign a24676 = ~a24674 & i372;
assign a24678 = ~a24676 & ~a12986;
assign a24680 = a24674 & ~i372;
assign a24682 = ~a24680 & ~a24678;
assign a24684 = ~a24682 & ~i374;
assign a24686 = ~a24684 & a12786;
assign a24688 = a24682 & i374;
assign a24690 = ~a24688 & ~a24686;
assign a24692 = ~a24690 & i376;
assign a24694 = ~a24692 & ~a12586;
assign a24696 = a24690 & ~i376;
assign a24698 = ~a24696 & ~a24694;
assign a24700 = ~a24698 & ~i380;
assign a24702 = ~a24700 & a12386;
assign a24704 = a24698 & i380;
assign a24706 = ~a24704 & ~a24702;
assign a24708 = ~a24706 & ~a24662;
assign a24710 = a12186 & ~i378;
assign a24712 = ~a24710 & ~a24708;
assign a24714 = a5580 & a4760;
assign a24716 = ~a16462 & a11214;
assign a24718 = ~a19886 & a16462;
assign a24722 = ~a24720 & ~a10706;
assign a24724 = ~a16344 & a11222;
assign a24726 = ~a19886 & a16344;
assign a24730 = ~a24728 & a10706;
assign a24732 = ~a24730 & ~a24722;
assign a24734 = ~a24732 & ~a8860;
assign a24736 = ~a16668 & a11230;
assign a24738 = ~a19886 & a16668;
assign a24742 = ~a24740 & ~a10706;
assign a24744 = ~a16802 & a11234;
assign a24746 = ~a19886 & a16802;
assign a24750 = ~a24748 & a10706;
assign a24752 = ~a24750 & ~a24742;
assign a24754 = ~a24752 & a8860;
assign a24756 = ~a24754 & ~a24734;
assign a24758 = ~a24756 & ~a8862;
assign a24760 = ~a16944 & a11246;
assign a24762 = ~a19886 & a16944;
assign a24766 = ~a24764 & ~a10706;
assign a24768 = ~a17076 & a11250;
assign a24770 = ~a19886 & a17076;
assign a24774 = ~a24772 & a10706;
assign a24776 = ~a24774 & ~a24766;
assign a24778 = ~a24776 & ~a8860;
assign a24780 = ~a17210 & a11258;
assign a24782 = ~a19886 & a17210;
assign a24786 = ~a24784 & ~a10706;
assign a24788 = ~a17344 & a11262;
assign a24790 = ~a19886 & a17344;
assign a24794 = ~a24792 & a10706;
assign a24796 = ~a24794 & ~a24786;
assign a24798 = ~a24796 & a8860;
assign a24800 = ~a24798 & ~a24778;
assign a24802 = ~a24800 & a8862;
assign a24804 = ~a24802 & ~a24758;
assign a24806 = ~a24804 & ~a8866;
assign a24808 = ~a17482 & a11202;
assign a24810 = ~a19886 & a17482;
assign a24814 = ~a24812 & ~a10706;
assign a24816 = ~a17720 & a11206;
assign a24818 = ~a19886 & a17720;
assign a24822 = ~a24820 & a10706;
assign a24824 = ~a24822 & ~a24814;
assign a24826 = ~a24824 & a8866;
assign a24828 = ~a24826 & ~a24806;
assign a24830 = ~a24828 & ~a5580;
assign a24832 = ~a24830 & ~a24714;
assign a24834 = a24832 & a13332;
assign a24836 = ~a24832 & ~a13332;
assign a24838 = ~a24836 & ~a24834;
assign a24840 = a5580 & a4752;
assign a24842 = ~a16462 & a11752;
assign a24844 = ~a19534 & a16462;
assign a24848 = ~a24846 & ~a10706;
assign a24850 = ~a16344 & a11756;
assign a24852 = ~a19534 & a16344;
assign a24856 = ~a24854 & a10706;
assign a24858 = ~a24856 & ~a24848;
assign a24860 = ~a24858 & ~a8860;
assign a24862 = ~a16668 & a11768;
assign a24864 = ~a19534 & a16668;
assign a24868 = ~a24866 & ~a10706;
assign a24870 = ~a16802 & a11776;
assign a24872 = ~a19534 & a16802;
assign a24876 = ~a24874 & a10706;
assign a24878 = ~a24876 & ~a24868;
assign a24880 = ~a24878 & a8860;
assign a24882 = ~a24880 & ~a24860;
assign a24884 = ~a24882 & ~a8862;
assign a24886 = ~a16944 & a11788;
assign a24888 = ~a19534 & a16944;
assign a24892 = ~a24890 & ~a10706;
assign a24894 = ~a17076 & a11792;
assign a24896 = ~a19534 & a17076;
assign a24900 = ~a24898 & a10706;
assign a24902 = ~a24900 & ~a24892;
assign a24904 = ~a24902 & ~a8860;
assign a24906 = ~a17210 & a11800;
assign a24908 = ~a19534 & a17210;
assign a24912 = ~a24910 & ~a10706;
assign a24914 = ~a17344 & a11804;
assign a24916 = ~a19534 & a17344;
assign a24920 = ~a24918 & a10706;
assign a24922 = ~a24920 & ~a24912;
assign a24924 = ~a24922 & a8860;
assign a24926 = ~a24924 & ~a24904;
assign a24928 = ~a24926 & a8862;
assign a24930 = ~a24928 & ~a24884;
assign a24932 = ~a24930 & ~a8866;
assign a24934 = ~a17482 & a11820;
assign a24936 = ~a19534 & a17482;
assign a24940 = ~a24938 & ~a10706;
assign a24942 = ~a17720 & a11824;
assign a24944 = ~a19534 & a17720;
assign a24948 = ~a24946 & a10706;
assign a24950 = ~a24948 & ~a24940;
assign a24952 = ~a24950 & a8866;
assign a24954 = ~a24952 & ~a24932;
assign a24956 = ~a24954 & ~a5580;
assign a24958 = ~a24956 & ~a24840;
assign a24960 = a24958 & a11998;
assign a24962 = ~a24958 & ~a11998;
assign a24964 = a5580 & a4738;
assign a24966 = ~a16462 & a12008;
assign a24968 = ~a19526 & a16462;
assign a24972 = ~a24970 & ~a10706;
assign a24974 = ~a16344 & a12016;
assign a24976 = ~a19526 & a16344;
assign a24980 = ~a24978 & a10706;
assign a24982 = ~a24980 & ~a24972;
assign a24984 = ~a24982 & ~a8860;
assign a24986 = ~a16668 & a12028;
assign a24988 = ~a19526 & a16668;
assign a24992 = ~a24990 & ~a10706;
assign a24994 = ~a16802 & a12036;
assign a24996 = ~a19526 & a16802;
assign a25000 = ~a24998 & a10706;
assign a25002 = ~a25000 & ~a24992;
assign a25004 = ~a25002 & a8860;
assign a25006 = ~a25004 & ~a24984;
assign a25008 = ~a25006 & ~a8862;
assign a25010 = ~a16944 & a12048;
assign a25012 = ~a19526 & a16944;
assign a25016 = ~a25014 & ~a10706;
assign a25018 = ~a17076 & a12052;
assign a25020 = ~a19526 & a17076;
assign a25024 = ~a25022 & a10706;
assign a25026 = ~a25024 & ~a25016;
assign a25028 = ~a25026 & ~a8860;
assign a25030 = ~a17210 & a12060;
assign a25032 = ~a19526 & a17210;
assign a25036 = ~a25034 & ~a10706;
assign a25038 = ~a17344 & a12064;
assign a25040 = ~a19526 & a17344;
assign a25044 = ~a25042 & a10706;
assign a25046 = ~a25044 & ~a25036;
assign a25048 = ~a25046 & a8860;
assign a25050 = ~a25048 & ~a25028;
assign a25052 = ~a25050 & a8862;
assign a25054 = ~a25052 & ~a25008;
assign a25056 = ~a25054 & ~a8866;
assign a25058 = ~a17482 & a12080;
assign a25060 = ~a19526 & a17482;
assign a25064 = ~a25062 & ~a10706;
assign a25066 = ~a17720 & a12084;
assign a25068 = ~a19526 & a17720;
assign a25072 = ~a25070 & a10706;
assign a25074 = ~a25072 & ~a25064;
assign a25076 = ~a25074 & a8866;
assign a25078 = ~a25076 & ~a25056;
assign a25080 = ~a25078 & ~a5580;
assign a25082 = ~a25080 & ~a24964;
assign a25084 = a25082 & ~a12186;
assign a25086 = ~a25082 & a12186;
assign a25088 = a5580 & a4722;
assign a25090 = ~a16462 & a12196;
assign a25092 = ~a19518 & a16462;
assign a25096 = ~a25094 & ~a10706;
assign a25098 = ~a16344 & a12204;
assign a25100 = ~a19518 & a16344;
assign a25104 = ~a25102 & a10706;
assign a25106 = ~a25104 & ~a25096;
assign a25108 = ~a25106 & ~a8860;
assign a25110 = ~a16668 & a12216;
assign a25112 = ~a19518 & a16668;
assign a25116 = ~a25114 & ~a10706;
assign a25118 = ~a16802 & a12224;
assign a25120 = ~a19518 & a16802;
assign a25124 = ~a25122 & a10706;
assign a25126 = ~a25124 & ~a25116;
assign a25128 = ~a25126 & a8860;
assign a25130 = ~a25128 & ~a25108;
assign a25132 = ~a25130 & ~a8862;
assign a25134 = ~a16944 & a12236;
assign a25136 = ~a19518 & a16944;
assign a25140 = ~a25138 & ~a10706;
assign a25142 = ~a17076 & a12240;
assign a25144 = ~a19518 & a17076;
assign a25148 = ~a25146 & a10706;
assign a25150 = ~a25148 & ~a25140;
assign a25152 = ~a25150 & ~a8860;
assign a25154 = ~a17210 & a12248;
assign a25156 = ~a19518 & a17210;
assign a25160 = ~a25158 & ~a10706;
assign a25162 = ~a17344 & a12252;
assign a25164 = ~a19518 & a17344;
assign a25168 = ~a25166 & a10706;
assign a25170 = ~a25168 & ~a25160;
assign a25172 = ~a25170 & a8860;
assign a25174 = ~a25172 & ~a25152;
assign a25176 = ~a25174 & a8862;
assign a25178 = ~a25176 & ~a25132;
assign a25180 = ~a25178 & ~a8866;
assign a25182 = ~a17482 & a12268;
assign a25184 = ~a19518 & a17482;
assign a25188 = ~a25186 & ~a10706;
assign a25190 = ~a17720 & a12272;
assign a25192 = ~a19518 & a17720;
assign a25196 = ~a25194 & a10706;
assign a25198 = ~a25196 & ~a25188;
assign a25200 = ~a25198 & a8866;
assign a25202 = ~a25200 & ~a25180;
assign a25204 = ~a25202 & ~a5580;
assign a25206 = ~a25204 & ~a25088;
assign a25208 = a25206 & ~a12386;
assign a25210 = ~a25206 & a12386;
assign a25212 = a5580 & a4706;
assign a25214 = ~a16462 & a12396;
assign a25216 = ~a19510 & a16462;
assign a25220 = ~a25218 & ~a10706;
assign a25222 = ~a16344 & a12404;
assign a25224 = ~a19510 & a16344;
assign a25228 = ~a25226 & a10706;
assign a25230 = ~a25228 & ~a25220;
assign a25232 = ~a25230 & ~a8860;
assign a25234 = ~a16668 & a12416;
assign a25236 = ~a19510 & a16668;
assign a25240 = ~a25238 & ~a10706;
assign a25242 = ~a16802 & a12424;
assign a25244 = ~a19510 & a16802;
assign a25248 = ~a25246 & a10706;
assign a25250 = ~a25248 & ~a25240;
assign a25252 = ~a25250 & a8860;
assign a25254 = ~a25252 & ~a25232;
assign a25256 = ~a25254 & ~a8862;
assign a25258 = ~a16944 & a12436;
assign a25260 = ~a19510 & a16944;
assign a25264 = ~a25262 & ~a10706;
assign a25266 = ~a17076 & a12440;
assign a25268 = ~a19510 & a17076;
assign a25272 = ~a25270 & a10706;
assign a25274 = ~a25272 & ~a25264;
assign a25276 = ~a25274 & ~a8860;
assign a25278 = ~a17210 & a12448;
assign a25280 = ~a19510 & a17210;
assign a25284 = ~a25282 & ~a10706;
assign a25286 = ~a17344 & a12452;
assign a25288 = ~a19510 & a17344;
assign a25292 = ~a25290 & a10706;
assign a25294 = ~a25292 & ~a25284;
assign a25296 = ~a25294 & a8860;
assign a25298 = ~a25296 & ~a25276;
assign a25300 = ~a25298 & a8862;
assign a25302 = ~a25300 & ~a25256;
assign a25304 = ~a25302 & ~a8866;
assign a25306 = ~a17482 & a12468;
assign a25308 = ~a19510 & a17482;
assign a25312 = ~a25310 & ~a10706;
assign a25314 = ~a17720 & a12472;
assign a25316 = ~a19510 & a17720;
assign a25320 = ~a25318 & a10706;
assign a25322 = ~a25320 & ~a25312;
assign a25324 = ~a25322 & a8866;
assign a25326 = ~a25324 & ~a25304;
assign a25328 = ~a25326 & ~a5580;
assign a25330 = ~a25328 & ~a25212;
assign a25332 = a25330 & ~a12586;
assign a25334 = ~a25330 & a12586;
assign a25336 = a5580 & a4690;
assign a25338 = ~a16462 & a12596;
assign a25340 = ~a19474 & a16462;
assign a25344 = ~a25342 & ~a10706;
assign a25346 = ~a16344 & a12604;
assign a25348 = ~a19474 & a16344;
assign a25352 = ~a25350 & a10706;
assign a25354 = ~a25352 & ~a25344;
assign a25356 = ~a25354 & ~a8860;
assign a25358 = ~a16668 & a12616;
assign a25360 = ~a19474 & a16668;
assign a25364 = ~a25362 & ~a10706;
assign a25366 = ~a16802 & a12624;
assign a25368 = ~a19474 & a16802;
assign a25372 = ~a25370 & a10706;
assign a25374 = ~a25372 & ~a25364;
assign a25376 = ~a25374 & a8860;
assign a25378 = ~a25376 & ~a25356;
assign a25380 = ~a25378 & ~a8862;
assign a25382 = ~a16944 & a12636;
assign a25384 = ~a19474 & a16944;
assign a25388 = ~a25386 & ~a10706;
assign a25390 = ~a17076 & a12640;
assign a25392 = ~a19474 & a17076;
assign a25396 = ~a25394 & a10706;
assign a25398 = ~a25396 & ~a25388;
assign a25400 = ~a25398 & ~a8860;
assign a25402 = ~a17210 & a12648;
assign a25404 = ~a19474 & a17210;
assign a25408 = ~a25406 & ~a10706;
assign a25410 = ~a17344 & a12652;
assign a25412 = ~a19474 & a17344;
assign a25416 = ~a25414 & a10706;
assign a25418 = ~a25416 & ~a25408;
assign a25420 = ~a25418 & a8860;
assign a25422 = ~a25420 & ~a25400;
assign a25424 = ~a25422 & a8862;
assign a25426 = ~a25424 & ~a25380;
assign a25428 = ~a25426 & ~a8866;
assign a25430 = ~a17482 & a12668;
assign a25432 = ~a19474 & a17482;
assign a25436 = ~a25434 & ~a10706;
assign a25438 = ~a17720 & a12672;
assign a25440 = ~a19474 & a17720;
assign a25444 = ~a25442 & a10706;
assign a25446 = ~a25444 & ~a25436;
assign a25448 = ~a25446 & a8866;
assign a25450 = ~a25448 & ~a25428;
assign a25452 = ~a25450 & ~a5580;
assign a25454 = ~a25452 & ~a25336;
assign a25456 = a25454 & ~a12786;
assign a25458 = ~a25454 & a12786;
assign a25460 = a5580 & a4672;
assign a25462 = ~a16462 & a12796;
assign a25464 = ~a19484 & a16462;
assign a25468 = ~a25466 & ~a10706;
assign a25470 = ~a16344 & a12804;
assign a25472 = ~a19484 & a16344;
assign a25476 = ~a25474 & a10706;
assign a25478 = ~a25476 & ~a25468;
assign a25480 = ~a25478 & ~a8860;
assign a25482 = ~a16668 & a12816;
assign a25484 = ~a19484 & a16668;
assign a25488 = ~a25486 & ~a10706;
assign a25490 = ~a16802 & a12824;
assign a25492 = ~a19484 & a16802;
assign a25496 = ~a25494 & a10706;
assign a25498 = ~a25496 & ~a25488;
assign a25500 = ~a25498 & a8860;
assign a25502 = ~a25500 & ~a25480;
assign a25504 = ~a25502 & ~a8862;
assign a25506 = ~a16944 & a12836;
assign a25508 = ~a19484 & a16944;
assign a25512 = ~a25510 & ~a10706;
assign a25514 = ~a17076 & a12840;
assign a25516 = ~a19484 & a17076;
assign a25520 = ~a25518 & a10706;
assign a25522 = ~a25520 & ~a25512;
assign a25524 = ~a25522 & ~a8860;
assign a25526 = ~a17210 & a12848;
assign a25528 = ~a19484 & a17210;
assign a25532 = ~a25530 & ~a10706;
assign a25534 = ~a17344 & a12852;
assign a25536 = ~a19484 & a17344;
assign a25540 = ~a25538 & a10706;
assign a25542 = ~a25540 & ~a25532;
assign a25544 = ~a25542 & a8860;
assign a25546 = ~a25544 & ~a25524;
assign a25548 = ~a25546 & a8862;
assign a25550 = ~a25548 & ~a25504;
assign a25552 = ~a25550 & ~a8866;
assign a25554 = ~a17482 & a12868;
assign a25556 = ~a19484 & a17482;
assign a25560 = ~a25558 & ~a10706;
assign a25562 = ~a17720 & a12872;
assign a25564 = ~a19484 & a17720;
assign a25568 = ~a25566 & a10706;
assign a25570 = ~a25568 & ~a25560;
assign a25572 = ~a25570 & a8866;
assign a25574 = ~a25572 & ~a25552;
assign a25576 = ~a25574 & ~a5580;
assign a25578 = ~a25576 & ~a25460;
assign a25580 = a25578 & ~a12986;
assign a25582 = ~a25578 & a12986;
assign a25584 = a5580 & a4656;
assign a25586 = ~a16462 & a11304;
assign a25588 = ~a19494 & a16462;
assign a25592 = ~a25590 & ~a10706;
assign a25594 = ~a16344 & a11316;
assign a25596 = ~a19494 & a16344;
assign a25600 = ~a25598 & a10706;
assign a25602 = ~a25600 & ~a25592;
assign a25604 = ~a25602 & ~a8860;
assign a25606 = ~a16668 & a11328;
assign a25608 = ~a19494 & a16668;
assign a25612 = ~a25610 & ~a10706;
assign a25614 = ~a16802 & a11336;
assign a25616 = ~a19494 & a16802;
assign a25620 = ~a25618 & a10706;
assign a25622 = ~a25620 & ~a25612;
assign a25624 = ~a25622 & a8860;
assign a25626 = ~a25624 & ~a25604;
assign a25628 = ~a25626 & ~a8862;
assign a25630 = ~a16944 & a11348;
assign a25632 = ~a19494 & a16944;
assign a25636 = ~a25634 & ~a10706;
assign a25638 = ~a17076 & a11352;
assign a25640 = ~a19494 & a17076;
assign a25644 = ~a25642 & a10706;
assign a25646 = ~a25644 & ~a25636;
assign a25648 = ~a25646 & ~a8860;
assign a25650 = ~a17210 & a11360;
assign a25652 = ~a19494 & a17210;
assign a25656 = ~a25654 & ~a10706;
assign a25658 = ~a17344 & a11364;
assign a25660 = ~a19494 & a17344;
assign a25664 = ~a25662 & a10706;
assign a25666 = ~a25664 & ~a25656;
assign a25668 = ~a25666 & a8860;
assign a25670 = ~a25668 & ~a25648;
assign a25672 = ~a25670 & a8862;
assign a25674 = ~a25672 & ~a25628;
assign a25676 = ~a25674 & ~a8866;
assign a25678 = ~a17482 & a11292;
assign a25680 = ~a19494 & a17482;
assign a25684 = ~a25682 & ~a10706;
assign a25686 = ~a17720 & a11296;
assign a25688 = ~a19494 & a17720;
assign a25692 = ~a25690 & a10706;
assign a25694 = ~a25692 & ~a25684;
assign a25696 = ~a25694 & a8866;
assign a25698 = ~a25696 & ~a25676;
assign a25700 = ~a25698 & ~a5580;
assign a25702 = ~a25700 & ~a25584;
assign a25704 = ~a25702 & a13158;
assign a25706 = ~a25704 & ~a25582;
assign a25708 = ~a25706 & ~a25580;
assign a25710 = ~a25708 & ~a25458;
assign a25712 = ~a25710 & ~a25456;
assign a25714 = ~a25712 & ~a25334;
assign a25716 = ~a25714 & ~a25332;
assign a25718 = ~a25716 & ~a25210;
assign a25720 = ~a25718 & ~a25208;
assign a25722 = ~a25720 & ~a25086;
assign a25724 = ~a25722 & ~a25084;
assign a25726 = ~a25724 & ~a24962;
assign a25728 = ~a25726 & ~a24960;
assign a25730 = a25728 & a24838;
assign a25732 = a8300 & ~i356;
assign a25734 = a8296 & ~a8220;
assign a25736 = ~a25734 & ~a25732;
assign a25738 = a25736 & ~l1686;
assign a25740 = l1686 & l1498;
assign a25742 = ~a25740 & ~a25738;
assign a25744 = ~i360 & i358;
assign a25746 = a25744 & a8846;
assign a25748 = a25746 & ~l1686;
assign a25750 = l1686 & l1500;
assign a25752 = ~a25750 & ~a25748;
assign a25754 = ~a11986 & ~l494;
assign a25756 = a25754 & ~a25752;
assign a25758 = a25756 & ~a25742;
assign a25760 = ~a25758 & ~a25730;
assign a25762 = a10706 & ~a8860;
assign a25764 = a25762 & a8866;
assign a25766 = a25764 & ~a8862;
assign a25768 = a25766 & ~a24720;
assign a25770 = ~a24720 & a10706;
assign a25772 = ~a24728 & ~a10706;
assign a25774 = ~a25772 & ~a25770;
assign a25776 = ~a10706 & a8860;
assign a25778 = ~a25776 & ~a25762;
assign a25780 = a25778 & ~a25774;
assign a25782 = ~a24740 & a10706;
assign a25784 = ~a24748 & ~a10706;
assign a25786 = ~a25784 & ~a25782;
assign a25788 = ~a25786 & ~a25778;
assign a25790 = ~a25788 & ~a25780;
assign a25792 = a10706 & a8860;
assign a25794 = ~a25792 & ~a8862;
assign a25796 = a25792 & a8862;
assign a25798 = ~a25796 & ~a25794;
assign a25800 = ~a25798 & ~a25790;
assign a25802 = ~a24764 & a10706;
assign a25804 = ~a24772 & ~a10706;
assign a25806 = ~a25804 & ~a25802;
assign a25808 = ~a25806 & a25778;
assign a25810 = ~a24784 & a10706;
assign a25812 = ~a24792 & ~a10706;
assign a25814 = ~a25812 & ~a25810;
assign a25816 = ~a25814 & ~a25778;
assign a25818 = ~a25816 & ~a25808;
assign a25820 = ~a25818 & a25798;
assign a25822 = ~a25820 & ~a25800;
assign a25824 = a25796 & ~a8866;
assign a25826 = ~a25796 & a8866;
assign a25828 = ~a25826 & ~a25824;
assign a25830 = a25828 & ~a25822;
assign a25832 = ~a24812 & a10706;
assign a25834 = ~a24820 & ~a10706;
assign a25836 = ~a25834 & ~a25832;
assign a25838 = ~a25836 & ~a25828;
assign a25840 = ~a25838 & ~a25830;
assign a25842 = ~a25840 & ~a25766;
assign a25844 = ~a25842 & ~a25768;
assign a25846 = ~a10706 & ~a5542;
assign a25848 = a10706 & ~a5548;
assign a25850 = ~a25848 & ~a25846;
assign a25852 = ~a25850 & ~a8860;
assign a25854 = ~a10706 & ~a5556;
assign a25856 = a10706 & ~a5572;
assign a25858 = ~a25856 & ~a25854;
assign a25860 = ~a25858 & a8860;
assign a25862 = ~a25860 & ~a25852;
assign a25864 = ~a25862 & ~a8862;
assign a25866 = ~a10706 & l576;
assign a25868 = a10706 & l578;
assign a25870 = ~a25868 & ~a25866;
assign a25872 = ~a25870 & ~a8860;
assign a25874 = ~a10706 & l580;
assign a25876 = a10706 & l582;
assign a25878 = ~a25876 & ~a25874;
assign a25880 = ~a25878 & a8860;
assign a25882 = ~a25880 & ~a25872;
assign a25884 = ~a25882 & a8862;
assign a25886 = ~a25884 & ~a25864;
assign a25888 = ~a25886 & ~a8866;
assign a25890 = ~a10706 & l586;
assign a25892 = a10706 & l584;
assign a25894 = ~a25892 & ~a25890;
assign a25896 = ~a25894 & a8866;
assign a25898 = ~a25896 & ~a25888;
assign a25900 = ~a11056 & ~a10706;
assign a25902 = a11056 & a10706;
assign a25904 = ~a25902 & ~a25900;
assign a25906 = ~a11066 & ~a8860;
assign a25908 = ~a25906 & a25904;
assign a25910 = ~a11076 & ~a8862;
assign a25912 = ~a25910 & a25908;
assign a25914 = ~a11088 & ~a8866;
assign a25916 = a11088 & a8866;
assign a25918 = ~a25916 & ~a25914;
assign a25920 = a11066 & a8860;
assign a25922 = ~a25920 & a25918;
assign a25924 = a11076 & a8862;
assign a25926 = ~a25924 & a25922;
assign a25928 = a25926 & a25912;
assign a25930 = ~a25928 & ~a25898;
assign a25932 = a25930 & ~a25844;
assign a25934 = ~a25930 & a4760;
assign a25936 = ~a25934 & ~a25932;
assign a25938 = a25936 & ~a24832;
assign a25940 = ~a25938 & ~a24834;
assign a25942 = a25936 & a13332;
assign a25944 = ~a25942 & ~a25940;
assign a25946 = a25766 & ~a24846;
assign a25948 = ~a24846 & a10706;
assign a25950 = ~a24854 & ~a10706;
assign a25952 = ~a25950 & ~a25948;
assign a25954 = ~a25952 & a25778;
assign a25956 = ~a24866 & a10706;
assign a25958 = ~a24874 & ~a10706;
assign a25960 = ~a25958 & ~a25956;
assign a25962 = ~a25960 & ~a25778;
assign a25964 = ~a25962 & ~a25954;
assign a25966 = ~a25964 & ~a25798;
assign a25968 = ~a24890 & a10706;
assign a25970 = ~a24898 & ~a10706;
assign a25972 = ~a25970 & ~a25968;
assign a25974 = ~a25972 & a25778;
assign a25976 = ~a24910 & a10706;
assign a25978 = ~a24918 & ~a10706;
assign a25980 = ~a25978 & ~a25976;
assign a25982 = ~a25980 & ~a25778;
assign a25984 = ~a25982 & ~a25974;
assign a25986 = ~a25984 & a25798;
assign a25988 = ~a25986 & ~a25966;
assign a25990 = ~a25988 & a25828;
assign a25992 = ~a24938 & a10706;
assign a25994 = ~a24946 & ~a10706;
assign a25996 = ~a25994 & ~a25992;
assign a25998 = ~a25996 & ~a25828;
assign a26000 = ~a25998 & ~a25990;
assign a26002 = ~a26000 & ~a25766;
assign a26004 = ~a26002 & ~a25946;
assign a26006 = ~a26004 & a25930;
assign a26008 = ~a25930 & a4752;
assign a26010 = ~a26008 & ~a26006;
assign a26012 = a26010 & a11998;
assign a26014 = ~a26010 & ~a11998;
assign a26016 = a25766 & ~a24970;
assign a26018 = ~a24970 & a10706;
assign a26020 = ~a24978 & ~a10706;
assign a26022 = ~a26020 & ~a26018;
assign a26024 = ~a26022 & a25778;
assign a26026 = ~a24990 & a10706;
assign a26028 = ~a24998 & ~a10706;
assign a26030 = ~a26028 & ~a26026;
assign a26032 = ~a26030 & ~a25778;
assign a26034 = ~a26032 & ~a26024;
assign a26036 = ~a26034 & ~a25798;
assign a26038 = ~a25014 & a10706;
assign a26040 = ~a25022 & ~a10706;
assign a26042 = ~a26040 & ~a26038;
assign a26044 = ~a26042 & a25778;
assign a26046 = ~a25034 & a10706;
assign a26048 = ~a25042 & ~a10706;
assign a26050 = ~a26048 & ~a26046;
assign a26052 = ~a26050 & ~a25778;
assign a26054 = ~a26052 & ~a26044;
assign a26056 = ~a26054 & a25798;
assign a26058 = ~a26056 & ~a26036;
assign a26060 = ~a26058 & a25828;
assign a26062 = ~a25062 & a10706;
assign a26064 = ~a25070 & ~a10706;
assign a26066 = ~a26064 & ~a26062;
assign a26068 = ~a26066 & ~a25828;
assign a26070 = ~a26068 & ~a26060;
assign a26072 = ~a26070 & ~a25766;
assign a26074 = ~a26072 & ~a26016;
assign a26076 = ~a26074 & a25930;
assign a26078 = ~a25930 & a4738;
assign a26080 = ~a26078 & ~a26076;
assign a26082 = a26080 & ~a12186;
assign a26084 = ~a26080 & a12186;
assign a26086 = a25766 & ~a25094;
assign a26088 = ~a25094 & a10706;
assign a26090 = ~a25102 & ~a10706;
assign a26092 = ~a26090 & ~a26088;
assign a26094 = ~a26092 & a25778;
assign a26096 = ~a25114 & a10706;
assign a26098 = ~a25122 & ~a10706;
assign a26100 = ~a26098 & ~a26096;
assign a26102 = ~a26100 & ~a25778;
assign a26104 = ~a26102 & ~a26094;
assign a26106 = ~a26104 & ~a25798;
assign a26108 = ~a25138 & a10706;
assign a26110 = ~a25146 & ~a10706;
assign a26112 = ~a26110 & ~a26108;
assign a26114 = ~a26112 & a25778;
assign a26116 = ~a25158 & a10706;
assign a26118 = ~a25166 & ~a10706;
assign a26120 = ~a26118 & ~a26116;
assign a26122 = ~a26120 & ~a25778;
assign a26124 = ~a26122 & ~a26114;
assign a26126 = ~a26124 & a25798;
assign a26128 = ~a26126 & ~a26106;
assign a26130 = ~a26128 & a25828;
assign a26132 = ~a25186 & a10706;
assign a26134 = ~a25194 & ~a10706;
assign a26136 = ~a26134 & ~a26132;
assign a26138 = ~a26136 & ~a25828;
assign a26140 = ~a26138 & ~a26130;
assign a26142 = ~a26140 & ~a25766;
assign a26144 = ~a26142 & ~a26086;
assign a26146 = ~a26144 & a25930;
assign a26148 = ~a25930 & a4722;
assign a26150 = ~a26148 & ~a26146;
assign a26152 = a26150 & ~a12386;
assign a26154 = ~a26150 & a12386;
assign a26156 = a25766 & ~a25218;
assign a26158 = ~a25218 & a10706;
assign a26160 = ~a25226 & ~a10706;
assign a26162 = ~a26160 & ~a26158;
assign a26164 = ~a26162 & a25778;
assign a26166 = ~a25238 & a10706;
assign a26168 = ~a25246 & ~a10706;
assign a26170 = ~a26168 & ~a26166;
assign a26172 = ~a26170 & ~a25778;
assign a26174 = ~a26172 & ~a26164;
assign a26176 = ~a26174 & ~a25798;
assign a26178 = ~a25262 & a10706;
assign a26180 = ~a25270 & ~a10706;
assign a26182 = ~a26180 & ~a26178;
assign a26184 = ~a26182 & a25778;
assign a26186 = ~a25282 & a10706;
assign a26188 = ~a25290 & ~a10706;
assign a26190 = ~a26188 & ~a26186;
assign a26192 = ~a26190 & ~a25778;
assign a26194 = ~a26192 & ~a26184;
assign a26196 = ~a26194 & a25798;
assign a26198 = ~a26196 & ~a26176;
assign a26200 = ~a26198 & a25828;
assign a26202 = ~a25310 & a10706;
assign a26204 = ~a25318 & ~a10706;
assign a26206 = ~a26204 & ~a26202;
assign a26208 = ~a26206 & ~a25828;
assign a26210 = ~a26208 & ~a26200;
assign a26212 = ~a26210 & ~a25766;
assign a26214 = ~a26212 & ~a26156;
assign a26216 = ~a26214 & a25930;
assign a26218 = ~a25930 & a4706;
assign a26220 = ~a26218 & ~a26216;
assign a26222 = a26220 & ~a12586;
assign a26224 = ~a26220 & a12586;
assign a26226 = a25766 & ~a25342;
assign a26228 = ~a25342 & a10706;
assign a26230 = ~a25350 & ~a10706;
assign a26232 = ~a26230 & ~a26228;
assign a26234 = ~a26232 & a25778;
assign a26236 = ~a25362 & a10706;
assign a26238 = ~a25370 & ~a10706;
assign a26240 = ~a26238 & ~a26236;
assign a26242 = ~a26240 & ~a25778;
assign a26244 = ~a26242 & ~a26234;
assign a26246 = ~a26244 & ~a25798;
assign a26248 = ~a25386 & a10706;
assign a26250 = ~a25394 & ~a10706;
assign a26252 = ~a26250 & ~a26248;
assign a26254 = ~a26252 & a25778;
assign a26256 = ~a25406 & a10706;
assign a26258 = ~a25414 & ~a10706;
assign a26260 = ~a26258 & ~a26256;
assign a26262 = ~a26260 & ~a25778;
assign a26264 = ~a26262 & ~a26254;
assign a26266 = ~a26264 & a25798;
assign a26268 = ~a26266 & ~a26246;
assign a26270 = ~a26268 & a25828;
assign a26272 = ~a25434 & a10706;
assign a26274 = ~a25442 & ~a10706;
assign a26276 = ~a26274 & ~a26272;
assign a26278 = ~a26276 & ~a25828;
assign a26280 = ~a26278 & ~a26270;
assign a26282 = ~a26280 & ~a25766;
assign a26284 = ~a26282 & ~a26226;
assign a26286 = ~a26284 & a25930;
assign a26288 = ~a25930 & a4690;
assign a26290 = ~a26288 & ~a26286;
assign a26292 = a26290 & ~a12786;
assign a26294 = ~a26290 & a12786;
assign a26296 = a25766 & ~a25466;
assign a26298 = ~a25466 & a10706;
assign a26300 = ~a25474 & ~a10706;
assign a26302 = ~a26300 & ~a26298;
assign a26304 = ~a26302 & a25778;
assign a26306 = ~a25486 & a10706;
assign a26308 = ~a25494 & ~a10706;
assign a26310 = ~a26308 & ~a26306;
assign a26312 = ~a26310 & ~a25778;
assign a26314 = ~a26312 & ~a26304;
assign a26316 = ~a26314 & ~a25798;
assign a26318 = ~a25510 & a10706;
assign a26320 = ~a25518 & ~a10706;
assign a26322 = ~a26320 & ~a26318;
assign a26324 = ~a26322 & a25778;
assign a26326 = ~a25530 & a10706;
assign a26328 = ~a25538 & ~a10706;
assign a26330 = ~a26328 & ~a26326;
assign a26332 = ~a26330 & ~a25778;
assign a26334 = ~a26332 & ~a26324;
assign a26336 = ~a26334 & a25798;
assign a26338 = ~a26336 & ~a26316;
assign a26340 = ~a26338 & a25828;
assign a26342 = ~a25558 & a10706;
assign a26344 = ~a25566 & ~a10706;
assign a26346 = ~a26344 & ~a26342;
assign a26348 = ~a26346 & ~a25828;
assign a26350 = ~a26348 & ~a26340;
assign a26352 = ~a26350 & ~a25766;
assign a26354 = ~a26352 & ~a26296;
assign a26356 = ~a26354 & a25930;
assign a26358 = ~a25930 & a4672;
assign a26360 = ~a26358 & ~a26356;
assign a26362 = a26360 & ~a12986;
assign a26364 = ~a26360 & a12986;
assign a26366 = a25766 & ~a25590;
assign a26368 = ~a25590 & a10706;
assign a26370 = ~a25598 & ~a10706;
assign a26372 = ~a26370 & ~a26368;
assign a26374 = ~a26372 & a25778;
assign a26376 = ~a25610 & a10706;
assign a26378 = ~a25618 & ~a10706;
assign a26380 = ~a26378 & ~a26376;
assign a26382 = ~a26380 & ~a25778;
assign a26384 = ~a26382 & ~a26374;
assign a26386 = ~a26384 & ~a25798;
assign a26388 = ~a25634 & a10706;
assign a26390 = ~a25642 & ~a10706;
assign a26392 = ~a26390 & ~a26388;
assign a26394 = ~a26392 & a25778;
assign a26396 = ~a25654 & a10706;
assign a26398 = ~a25662 & ~a10706;
assign a26400 = ~a26398 & ~a26396;
assign a26402 = ~a26400 & ~a25778;
assign a26404 = ~a26402 & ~a26394;
assign a26406 = ~a26404 & a25798;
assign a26408 = ~a26406 & ~a26386;
assign a26410 = ~a26408 & a25828;
assign a26412 = ~a25682 & a10706;
assign a26414 = ~a25690 & ~a10706;
assign a26416 = ~a26414 & ~a26412;
assign a26418 = ~a26416 & ~a25828;
assign a26420 = ~a26418 & ~a26410;
assign a26422 = ~a26420 & ~a25766;
assign a26424 = ~a26422 & ~a26366;
assign a26426 = ~a26424 & a25930;
assign a26428 = ~a25930 & a4656;
assign a26430 = ~a26428 & ~a26426;
assign a26432 = ~a26430 & a13158;
assign a26434 = ~a26432 & ~a26364;
assign a26436 = ~a26434 & ~a26362;
assign a26438 = ~a26436 & ~a26294;
assign a26440 = ~a26438 & ~a26292;
assign a26442 = ~a26440 & ~a26224;
assign a26444 = ~a26442 & ~a26222;
assign a26446 = ~a26444 & ~a26154;
assign a26448 = ~a26446 & ~a26152;
assign a26450 = ~a26448 & ~a26084;
assign a26452 = ~a26450 & ~a26082;
assign a26454 = ~a26452 & ~a26014;
assign a26456 = ~a26454 & ~a26012;
assign a26458 = a26456 & a25944;
assign a26460 = ~a25728 & a24838;
assign a26462 = ~a26460 & ~a26458;
assign a26464 = ~a25936 & a24832;
assign a26466 = ~a26464 & ~a25938;
assign a26468 = a26466 & ~a26456;
assign a26470 = ~a26468 & ~a26462;
assign a26472 = a26470 & a25742;
assign a26474 = ~a11998 & a2548;
assign a26476 = a11998 & ~a2548;
assign a26478 = a12186 & a4404;
assign a26480 = ~a12186 & ~a4404;
assign a26482 = a12386 & a2566;
assign a26484 = ~a12386 & ~a2566;
assign a26486 = a12586 & a4428;
assign a26488 = ~a12586 & ~a4428;
assign a26490 = a12786 & a4464;
assign a26492 = ~a12786 & ~a4464;
assign a26494 = a12986 & a4500;
assign a26496 = ~a12986 & ~a4500;
assign a26498 = ~a13158 & ~a4536;
assign a26500 = ~a26498 & ~a26496;
assign a26502 = ~a26500 & ~a26494;
assign a26504 = ~a26502 & ~a26492;
assign a26506 = ~a26504 & ~a26490;
assign a26508 = ~a26506 & ~a26488;
assign a26510 = ~a26508 & ~a26486;
assign a26512 = ~a26510 & ~a26484;
assign a26514 = ~a26512 & ~a26482;
assign a26516 = ~a26514 & ~a26480;
assign a26518 = ~a26516 & ~a26478;
assign a26520 = ~a26518 & ~a26476;
assign a26522 = ~a26520 & ~a26474;
assign a26524 = a13332 & l532;
assign a26526 = a2268 & l994;
assign a26528 = ~a26526 & ~a26524;
assign a26530 = a26528 & ~a26522;
assign a26532 = ~a26530 & a26472;
assign a26534 = ~a26528 & a26522;
assign a26536 = ~a26534 & a26532;
assign a26538 = ~a26536 & a25760;
assign a26540 = ~a26538 & a24712;
assign a26542 = a26540 & a11998;
assign a26544 = ~a26542 & a13332;
assign a26546 = a26542 & ~a13332;
assign a26548 = ~a26546 & ~a26544;
assign a26550 = ~a26548 & ~a11986;
assign a26552 = ~a25082 & i378;
assign a26554 = a25206 & i380;
assign a26556 = ~a25206 & ~i380;
assign a26558 = a25330 & i376;
assign a26560 = ~a25330 & ~i376;
assign a26562 = a25454 & i374;
assign a26564 = ~a25454 & ~i374;
assign a26566 = ~a25578 & ~i372;
assign a26568 = ~a25702 & ~a24672;
assign a26570 = ~a26568 & ~a26566;
assign a26572 = a25578 & i372;
assign a26574 = ~a26572 & ~a26570;
assign a26576 = ~a26574 & ~a26564;
assign a26578 = ~a26576 & ~a26562;
assign a26580 = ~a26578 & ~a26560;
assign a26582 = ~a26580 & ~a26558;
assign a26584 = ~a26582 & ~a26556;
assign a26586 = ~a26584 & ~a26554;
assign a26588 = ~a26586 & ~a26552;
assign a26590 = a25082 & ~i378;
assign a26592 = ~a26590 & ~a26588;
assign a26594 = a26592 & ~a24958;
assign a26596 = a26594 & a24832;
assign a26598 = ~a26594 & ~a24832;
assign a26600 = ~a26598 & ~a26596;
assign a26602 = ~a26600 & a11986;
assign a26606 = a22712 & a22696;
assign a26608 = a26606 & a22688;
assign a26610 = ~a26608 & a10854;
assign a26612 = a26608 & ~a10862;
assign a26618 = ~a22654 & a10846;
assign a26620 = a22654 & ~a10862;
assign a26624 = ~a26540 & ~a11998;
assign a26626 = ~a26624 & ~a26542;
assign a26628 = a26626 & ~a11986;
assign a26630 = ~a26592 & a24958;
assign a26632 = ~a26630 & ~a26594;
assign a26634 = a26632 & a11986;
assign a26638 = a26636 & a2548;
assign a26640 = ~a26636 & ~a2548;
assign a26642 = a26538 & ~a12186;
assign a26644 = ~a24710 & ~a24662;
assign a26646 = ~a26644 & ~a24706;
assign a26648 = a26644 & a24706;
assign a26650 = ~a26648 & ~a26646;
assign a26652 = a26650 & ~a26538;
assign a26654 = ~a26652 & ~a26642;
assign a26656 = ~a26654 & ~a11986;
assign a26658 = ~a26590 & ~a26552;
assign a26660 = ~a26658 & a26586;
assign a26662 = a26658 & ~a26586;
assign a26664 = ~a26662 & ~a26660;
assign a26666 = ~a26664 & a11986;
assign a26668 = ~a26666 & ~a26656;
assign a26670 = a26668 & a4404;
assign a26672 = ~a26668 & ~a4404;
assign a26674 = ~a24704 & ~a24700;
assign a26676 = a26674 & ~a26538;
assign a26678 = ~a26676 & a12386;
assign a26680 = a26676 & ~a12386;
assign a26682 = ~a26680 & ~a26678;
assign a26684 = a26682 & ~a11986;
assign a26686 = ~a26556 & ~a26554;
assign a26688 = ~a26686 & a26582;
assign a26690 = a26584 & ~a26554;
assign a26692 = ~a26690 & ~a26688;
assign a26694 = ~a26692 & a11986;
assign a26696 = ~a26694 & ~a26684;
assign a26698 = a26696 & a2566;
assign a26700 = ~a26696 & ~a2566;
assign a26702 = ~a24696 & ~a24692;
assign a26704 = a26702 & ~a26538;
assign a26706 = ~a26704 & a12586;
assign a26708 = a26704 & ~a12586;
assign a26710 = ~a26708 & ~a26706;
assign a26712 = a26710 & ~a11986;
assign a26714 = ~a26560 & ~a26558;
assign a26716 = ~a26714 & a26578;
assign a26718 = a26580 & ~a26558;
assign a26720 = ~a26718 & ~a26716;
assign a26722 = ~a26720 & a11986;
assign a26724 = ~a26722 & ~a26712;
assign a26726 = a26724 & a4428;
assign a26728 = ~a26724 & ~a4428;
assign a26730 = ~a24688 & ~a24684;
assign a26732 = a26730 & ~a26538;
assign a26734 = ~a26732 & a12786;
assign a26736 = a26732 & ~a12786;
assign a26738 = ~a26736 & ~a26734;
assign a26740 = a26738 & ~a11986;
assign a26742 = ~a26564 & ~a26562;
assign a26744 = ~a26742 & a26574;
assign a26746 = a26576 & ~a26562;
assign a26748 = ~a26746 & ~a26744;
assign a26750 = ~a26748 & a11986;
assign a26752 = ~a26750 & ~a26740;
assign a26754 = a26752 & a4464;
assign a26756 = ~a26752 & ~a4464;
assign a26758 = ~a24680 & ~a24676;
assign a26760 = a26758 & ~a26538;
assign a26762 = ~a26760 & a12986;
assign a26764 = a26760 & ~a12986;
assign a26766 = ~a26764 & ~a26762;
assign a26768 = a26766 & ~a11986;
assign a26770 = ~a26572 & ~a26566;
assign a26772 = ~a26770 & a26568;
assign a26774 = a26770 & ~a26568;
assign a26776 = ~a26774 & ~a26772;
assign a26778 = ~a26776 & a11986;
assign a26780 = ~a26778 & ~a26768;
assign a26782 = a26780 & a4500;
assign a26784 = ~a26780 & ~a4500;
assign a26786 = ~a26538 & ~a24672;
assign a26788 = ~a26786 & a13158;
assign a26790 = ~a26538 & a24674;
assign a26792 = ~a26790 & ~a26788;
assign a26794 = a26792 & ~a11986;
assign a26796 = a25702 & a24672;
assign a26798 = ~a26796 & ~a26568;
assign a26800 = a26798 & a11986;
assign a26802 = ~a26800 & ~a26794;
assign a26804 = ~a26802 & ~a4536;
assign a26806 = ~a26804 & ~a26784;
assign a26808 = ~a26806 & ~a26782;
assign a26810 = ~a26808 & ~a26756;
assign a26812 = ~a26810 & ~a26754;
assign a26814 = ~a26812 & ~a26728;
assign a26816 = ~a26814 & ~a26726;
assign a26818 = ~a26816 & ~a26700;
assign a26820 = ~a26818 & ~a26698;
assign a26822 = ~a26820 & ~a26672;
assign a26824 = ~a26822 & ~a26670;
assign a26826 = ~a26824 & ~a26640;
assign a26828 = ~a26826 & ~a26638;
assign a26830 = ~a26604 & ~a2268;
assign a26832 = a26604 & a2268;
assign a26834 = ~a26832 & ~a26830;
assign a26836 = a26834 & ~a26828;
assign a26838 = ~a26834 & a26828;
assign a26840 = ~a26838 & ~a26836;
assign a26842 = ~a26636 & a26010;
assign a26844 = a26636 & ~a26010;
assign a26846 = ~a26668 & a26080;
assign a26848 = a26668 & ~a26080;
assign a26850 = ~a26696 & a26150;
assign a26852 = a26696 & ~a26150;
assign a26854 = ~a26724 & a26220;
assign a26856 = a26724 & ~a26220;
assign a26858 = ~a26752 & a26290;
assign a26860 = a26752 & ~a26290;
assign a26862 = ~a26780 & a26360;
assign a26864 = a26780 & ~a26360;
assign a26866 = a26802 & ~a26430;
assign a26868 = ~a26866 & ~a26864;
assign a26870 = ~a26868 & ~a26862;
assign a26872 = ~a26870 & ~a26860;
assign a26874 = ~a26872 & ~a26858;
assign a26876 = ~a26874 & ~a26856;
assign a26878 = ~a26876 & ~a26854;
assign a26880 = ~a26878 & ~a26852;
assign a26882 = ~a26880 & ~a26850;
assign a26884 = ~a26882 & ~a26848;
assign a26886 = ~a26884 & ~a26846;
assign a26888 = ~a26886 & ~a26844;
assign a26890 = ~a26888 & ~a26842;
assign a26892 = ~a26604 & a24832;
assign a26894 = a26604 & ~a24832;
assign a26896 = ~a26894 & ~a26892;
assign a26898 = ~a26636 & a24958;
assign a26900 = a26636 & ~a24958;
assign a26902 = ~a26668 & a25082;
assign a26904 = a26668 & ~a25082;
assign a26906 = ~a26696 & a25206;
assign a26908 = a26696 & ~a25206;
assign a26910 = ~a26724 & a25330;
assign a26912 = a26724 & ~a25330;
assign a26914 = ~a26752 & a25454;
assign a26916 = a26752 & ~a25454;
assign a26918 = ~a26780 & a25578;
assign a26920 = a26780 & ~a25578;
assign a26922 = a26802 & ~a25702;
assign a26924 = ~a26922 & ~a26920;
assign a26926 = ~a26924 & ~a26918;
assign a26928 = ~a26926 & ~a26916;
assign a26930 = ~a26928 & ~a26914;
assign a26932 = ~a26930 & ~a26912;
assign a26934 = ~a26932 & ~a26910;
assign a26936 = ~a26934 & ~a26908;
assign a26938 = ~a26936 & ~a26906;
assign a26940 = ~a26938 & ~a26904;
assign a26942 = ~a26940 & ~a26902;
assign a26944 = ~a26942 & ~a26900;
assign a26946 = ~a26944 & ~a26898;
assign a26948 = ~a26946 & a26896;
assign a26950 = a26948 & a26890;
assign a26952 = ~a26604 & a25936;
assign a26954 = a26604 & ~a25936;
assign a26956 = ~a26954 & ~a26952;
assign a26958 = a26956 & a26890;
assign a26960 = ~a26958 & ~a26948;
assign a26962 = ~a26960 & ~a26466;
assign a26964 = ~a26962 & ~a26950;
assign a26966 = ~a26964 & a26840;
assign a26968 = ~a26966 & ~a25928;
assign a26970 = a26968 & ~a11986;
assign a26972 = ~a8862 & ~a6592;
assign a26974 = a8862 & a6592;
assign a26976 = ~a26974 & ~a26972;
assign a26978 = ~a8866 & ~a6476;
assign a26980 = a8866 & a6476;
assign a26982 = ~a26980 & ~a26978;
assign a26984 = a26982 & a26976;
assign a26986 = ~a8860 & ~a6548;
assign a26988 = a8860 & a6548;
assign a26990 = ~a26988 & ~a26986;
assign a26992 = ~a10706 & ~a6512;
assign a26994 = a10706 & a6512;
assign a26996 = ~a26994 & ~a26992;
assign a26998 = a26996 & a26990;
assign a27000 = a26998 & a26984;
assign a27002 = ~a10706 & ~a6522;
assign a27004 = ~a27002 & a27000;
assign a27006 = a8862 & a6608;
assign a27008 = ~a27006 & a27004;
assign a27010 = a10706 & a6522;
assign a27012 = ~a8866 & ~a6494;
assign a27014 = ~a27012 & ~a27010;
assign a27016 = a27014 & a27008;
assign a27018 = a8860 & a6566;
assign a27020 = ~a8862 & ~a6608;
assign a27022 = ~a27020 & ~a27018;
assign a27024 = a8866 & a6494;
assign a27026 = ~a8860 & ~a6566;
assign a27028 = ~a27026 & ~a27024;
assign a27030 = a27028 & a27022;
assign a27032 = a27030 & a27016;
assign a27034 = ~a27032 & a26970;
assign a27036 = a27034 & a25766;
assign a27038 = a27036 & i400;
assign a27040 = a27034 & ~a25766;
assign a27042 = a27040 & i398;
assign a27044 = ~a27042 & ~a27038;
assign a27046 = a27044 & a8866;
assign a27048 = a27042 & ~a25828;
assign a27050 = ~a27048 & ~a27046;
assign a27052 = ~a27050 & ~a24508;
assign a27054 = a24508 & ~a6476;
assign a27056 = ~a27054 & ~a27052;
assign a27058 = ~a27056 & ~l494;
assign a27062 = ~a13508 & a8874;
assign a27064 = ~a24490 & ~a24444;
assign a27066 = ~a27064 & a24486;
assign a27068 = a27064 & ~a24486;
assign a27070 = ~a27068 & ~a27066;
assign a27072 = ~a27070 & a13508;
assign a27074 = ~a27072 & ~a27062;
assign a27076 = ~a27074 & a24518;
assign a27078 = ~a24568 & ~a24522;
assign a27080 = ~a27078 & a24564;
assign a27082 = a27078 & ~a24564;
assign a27084 = ~a27082 & ~a27080;
assign a27086 = ~a27084 & ~a24518;
assign a27088 = ~a27086 & ~a27076;
assign a27090 = ~a27088 & ~l1494;
assign a27092 = ~a24636 & ~a24590;
assign a27094 = ~a27092 & a24632;
assign a27096 = a27092 & ~a24632;
assign a27098 = ~a27096 & ~a27094;
assign a27100 = ~a27098 & l1494;
assign a27102 = ~a27100 & ~a27090;
assign a27104 = ~a27102 & a13494;
assign a27106 = ~a13494 & a11486;
assign a27110 = ~a13508 & a10044;
assign a27112 = ~a24484 & ~a24446;
assign a27114 = ~a27112 & a24480;
assign a27116 = a27112 & ~a24480;
assign a27118 = ~a27116 & ~a27114;
assign a27120 = ~a27118 & a13508;
assign a27122 = ~a27120 & ~a27110;
assign a27124 = ~a27122 & a24518;
assign a27126 = ~a24562 & ~a24524;
assign a27128 = ~a27126 & a24558;
assign a27130 = a27126 & ~a24558;
assign a27132 = ~a27130 & ~a27128;
assign a27134 = ~a27132 & ~a24518;
assign a27136 = ~a27134 & ~a27124;
assign a27138 = ~a27136 & ~l1494;
assign a27140 = ~a24630 & ~a24592;
assign a27142 = ~a27140 & a24626;
assign a27144 = a27140 & ~a24626;
assign a27146 = ~a27144 & ~a27142;
assign a27148 = ~a27146 & l1494;
assign a27150 = ~a27148 & ~a27138;
assign a27152 = ~a27150 & a13494;
assign a27154 = ~a13494 & a11478;
assign a27158 = ~a13508 & a10074;
assign a27160 = ~a24478 & ~a24448;
assign a27162 = ~a27160 & a24474;
assign a27164 = a27160 & ~a24474;
assign a27166 = ~a27164 & ~a27162;
assign a27168 = ~a27166 & a13508;
assign a27170 = ~a27168 & ~a27158;
assign a27172 = ~a27170 & a24518;
assign a27174 = ~a24556 & ~a24526;
assign a27176 = ~a27174 & a24552;
assign a27178 = a27174 & ~a24552;
assign a27180 = ~a27178 & ~a27176;
assign a27182 = ~a27180 & ~a24518;
assign a27184 = ~a27182 & ~a27172;
assign a27186 = ~a27184 & ~l1494;
assign a27188 = ~a24624 & ~a24594;
assign a27190 = ~a27188 & a24620;
assign a27192 = a27188 & ~a24620;
assign a27194 = ~a27192 & ~a27190;
assign a27196 = ~a27194 & l1494;
assign a27198 = ~a27196 & ~a27186;
assign a27200 = ~a27198 & a13494;
assign a27202 = ~a13494 & a11472;
assign a27206 = ~a13508 & a10100;
assign a27208 = ~a24472 & ~a24450;
assign a27210 = ~a27208 & a24468;
assign a27212 = a27208 & ~a24468;
assign a27214 = ~a27212 & ~a27210;
assign a27216 = ~a27214 & a13508;
assign a27218 = ~a27216 & ~a27206;
assign a27220 = ~a27218 & a24518;
assign a27222 = ~a24550 & ~a24528;
assign a27224 = ~a27222 & a24546;
assign a27226 = a27222 & ~a24546;
assign a27228 = ~a27226 & ~a27224;
assign a27230 = ~a27228 & ~a24518;
assign a27232 = ~a27230 & ~a27220;
assign a27234 = ~a27232 & ~l1494;
assign a27236 = ~a24618 & ~a24596;
assign a27238 = ~a27236 & a24614;
assign a27240 = a27236 & ~a24614;
assign a27242 = ~a27240 & ~a27238;
assign a27244 = ~a27242 & l1494;
assign a27246 = ~a27244 & ~a27234;
assign a27248 = ~a27246 & a13494;
assign a27250 = ~a13494 & a11462;
assign a27254 = ~a13508 & a10126;
assign a27256 = ~a24466 & ~a24452;
assign a27258 = ~a27256 & a24462;
assign a27260 = a27256 & ~a24462;
assign a27262 = ~a27260 & ~a27258;
assign a27264 = ~a27262 & a13508;
assign a27266 = ~a27264 & ~a27254;
assign a27268 = ~a27266 & a24518;
assign a27270 = ~a24544 & ~a24530;
assign a27272 = ~a27270 & a24540;
assign a27274 = a27270 & ~a24540;
assign a27276 = ~a27274 & ~a27272;
assign a27278 = ~a27276 & ~a24518;
assign a27280 = ~a27278 & ~a27268;
assign a27282 = ~a27280 & ~l1494;
assign a27284 = ~a24612 & ~a24598;
assign a27286 = ~a27284 & a24608;
assign a27288 = a27284 & ~a24608;
assign a27290 = ~a27288 & ~a27286;
assign a27292 = ~a27290 & l1494;
assign a27294 = ~a27292 & ~a27282;
assign a27296 = ~a27294 & a13494;
assign a27298 = ~a13494 & a11452;
assign a27302 = ~a13508 & a10152;
assign a27304 = ~a24460 & ~a24454;
assign a27306 = ~a27304 & a24456;
assign a27308 = a27304 & ~a24456;
assign a27310 = ~a27308 & ~a27306;
assign a27312 = ~a27310 & a13508;
assign a27314 = ~a27312 & ~a27302;
assign a27316 = ~a27314 & a24518;
assign a27318 = ~a24538 & ~a24532;
assign a27320 = ~a27318 & a24534;
assign a27322 = ~a24538 & a24536;
assign a27324 = ~a27322 & ~a27320;
assign a27326 = ~a27324 & ~a24518;
assign a27328 = ~a27326 & ~a27316;
assign a27330 = ~a27328 & ~l1494;
assign a27332 = ~a24606 & ~a24600;
assign a27334 = ~a27332 & a24602;
assign a27336 = ~a24606 & a24604;
assign a27338 = ~a27336 & ~a27334;
assign a27340 = ~a27338 & l1494;
assign a27342 = ~a27340 & ~a27330;
assign a27344 = ~a27342 & a13494;
assign a27346 = ~a13494 & a11442;
assign a27350 = a24258 & a13508;
assign a27352 = ~a27350 & a10178;
assign a27354 = a27350 & ~a10178;
assign a27356 = ~a27354 & ~a27352;
assign a27358 = ~a27356 & a24518;
assign a27360 = ~a24258 & ~a11432;
assign a27362 = ~a27360 & ~a24518;
assign a27364 = a27362 & ~a24534;
assign a27366 = ~a27364 & ~a27358;
assign a27368 = ~a27366 & ~l1494;
assign a27370 = ~a24258 & ~a15350;
assign a27372 = ~a27370 & l1494;
assign a27374 = a27372 & ~a24602;
assign a27376 = ~a27374 & ~a27368;
assign a27378 = ~a27376 & a13494;
assign a27380 = ~a13494 & a11432;
assign a27384 = ~a27042 & a8862;
assign a27386 = a27042 & a25798;
assign a27388 = ~a27386 & ~a27384;
assign a27390 = ~a27388 & ~a24508;
assign a27392 = a24508 & ~a6592;
assign a27394 = ~a27392 & ~a27390;
assign a27396 = ~a27394 & ~l494;
assign a27400 = ~a27042 & a8860;
assign a27402 = a27042 & ~a25778;
assign a27404 = ~a27402 & ~a27400;
assign a27406 = ~a27404 & ~a24508;
assign a27408 = a24508 & ~a6548;
assign a27410 = ~a27408 & ~a27406;
assign a27412 = ~a27410 & ~l494;
assign a27416 = a27044 & a10706;
assign a27418 = a27042 & ~a10706;
assign a27420 = ~a27418 & ~a27416;
assign a27422 = ~a27420 & ~a24508;
assign a27424 = a24508 & ~a6512;
assign a27426 = ~a27424 & ~a27422;
assign a27428 = ~a27426 & ~l494;
assign a27432 = l1686 & l1560;
assign a27434 = ~a27432 & ~a5538;
assign a27436 = l1686 & ~l1562;
assign a27438 = l1686 & ~l1564;
assign a27440 = ~a27438 & ~a27436;
assign a27442 = a27440 & ~a27434;
assign a27444 = ~a27442 & a8068;
assign a27446 = ~a27444 & ~l494;
assign a27448 = a22686 & i440;
assign a27450 = ~a27448 & ~a10802;
assign a27456 = ~a26608 & a10790;
assign a27458 = a26608 & ~a10798;
assign a27462 = ~a22654 & a10760;
assign a27464 = a22654 & ~a10798;
assign a27468 = ~a26608 & a10940;
assign a27470 = a26608 & ~a10948;
assign a27474 = ~a22654 & a10932;
assign a27476 = a22654 & ~a10948;
assign a27480 = ~a26608 & a10898;
assign a27482 = a26608 & ~a10906;
assign a27486 = ~a22654 & a10890;
assign a27488 = a22654 & ~a10906;
assign a27492 = l1686 & ~l1490;
assign a27494 = a11986 & ~a6934;
assign a27496 = ~a27494 & ~l494;
assign a27500 = ~a16548 & ~a16544;
assign a27502 = a27500 & ~a16570;
assign a27504 = a27502 & ~a16554;
assign a27506 = ~a27504 & ~a5542;
assign a27508 = ~a11630 & a8860;
assign a27510 = a11750 & ~a10706;
assign a27512 = ~a27510 & ~a27508;
assign a27514 = a8862 & l1090;
assign a27516 = ~a11750 & a10706;
assign a27518 = ~a27516 & ~a27514;
assign a27520 = a27518 & a27512;
assign a27522 = a11624 & l1058;
assign a27524 = a11630 & ~a8860;
assign a27526 = ~a27524 & ~a27522;
assign a27528 = a8866 & l1082;
assign a27530 = a11622 & l1010;
assign a27532 = ~a27530 & ~a27528;
assign a27534 = a27532 & a27526;
assign a27536 = a27534 & a27520;
assign a27538 = ~a19362 & a11114;
assign a27540 = a25758 & ~a8866;
assign a27542 = ~a25758 & i366;
assign a27544 = a25758 & ~a10706;
assign a27546 = ~a27544 & ~a27542;
assign a27548 = ~a27546 & a27540;
assign a27550 = ~a25758 & i364;
assign a27552 = a25758 & ~a8860;
assign a27554 = ~a27552 & ~a27550;
assign a27556 = ~a27554 & a27548;
assign a27558 = ~a25758 & i362;
assign a27560 = a25758 & ~a8862;
assign a27562 = ~a27560 & ~a27558;
assign a27564 = ~a27562 & a27556;
assign a27566 = a27564 & a27538;
assign a27568 = ~a27566 & a11842;
assign a27570 = ~a27568 & ~a1690;
assign a27574 = a27572 & ~a11750;
assign a27576 = a27546 & a27540;
assign a27578 = a27576 & ~a27554;
assign a27580 = a27578 & ~a27562;
assign a27582 = a27580 & a27538;
assign a27584 = ~a27582 & a11850;
assign a27586 = ~a27584 & ~a1690;
assign a27590 = a27588 & a11750;
assign a27592 = ~a27590 & ~a27574;
assign a27594 = a11730 & ~l1686;
assign a27596 = l1686 & l1558;
assign a27598 = ~a27596 & ~a27594;
assign a27600 = a13508 & ~a11842;
assign a27602 = ~a27600 & a27598;
assign a27604 = a14070 & a14058;
assign a27606 = a13522 & a13068;
assign a27608 = ~a27606 & ~a14076;
assign a27610 = a27608 & a14084;
assign a27612 = a27610 & a27604;
assign a27614 = ~a14074 & ~a14072;
assign a27616 = a27614 & a14064;
assign a27618 = ~a14100 & ~a14078;
assign a27620 = a27618 & a14108;
assign a27622 = a27620 & a27616;
assign a27624 = a27622 & a27612;
assign a27626 = ~a27624 & a13508;
assign a27628 = ~a27626 & ~a27602;
assign a27632 = a27630 & ~a11750;
assign a27634 = a13508 & ~a11850;
assign a27636 = ~a27634 & ~l1556;
assign a27638 = a14738 & a14726;
assign a27640 = a13522 & a13078;
assign a27642 = ~a27640 & ~a14744;
assign a27644 = a27642 & a14752;
assign a27646 = a27644 & a27638;
assign a27648 = ~a14742 & ~a14740;
assign a27650 = a27648 & a14732;
assign a27652 = ~a14768 & ~a14746;
assign a27654 = a27652 & a14776;
assign a27656 = a27654 & a27650;
assign a27658 = a27656 & a27646;
assign a27660 = ~a27658 & a13508;
assign a27662 = ~a27660 & ~a27636;
assign a27666 = a27664 & a11750;
assign a27668 = ~a27666 & ~a27632;
assign a27670 = a27668 & ~a27592;
assign a27672 = ~a27670 & ~a11630;
assign a27674 = a27554 & a27548;
assign a27676 = a27674 & ~a27562;
assign a27678 = a27676 & a27538;
assign a27680 = ~a27678 & ~l1104;
assign a27682 = ~a27680 & ~a1690;
assign a27686 = a27684 & ~a11750;
assign a27688 = a27576 & a27554;
assign a27690 = a27688 & ~a27562;
assign a27692 = a27690 & a27538;
assign a27694 = ~a27692 & ~l1102;
assign a27696 = ~a27694 & ~a1690;
assign a27700 = a27698 & a11750;
assign a27702 = ~a27700 & ~a27686;
assign a27704 = a13508 & l1104;
assign a27706 = ~a27704 & ~l1554;
assign a27708 = a14574 & a14562;
assign a27710 = a13522 & a13086;
assign a27712 = ~a27710 & ~a14580;
assign a27714 = a27712 & a14588;
assign a27716 = a27714 & a27708;
assign a27718 = ~a14578 & ~a14576;
assign a27720 = a27718 & a14568;
assign a27722 = ~a14604 & ~a14582;
assign a27724 = a27722 & a14612;
assign a27726 = a27724 & a27720;
assign a27728 = a27726 & a27716;
assign a27730 = ~a27728 & a13508;
assign a27732 = ~a27730 & ~a27706;
assign a27736 = a27734 & ~a11750;
assign a27738 = a13508 & l1102;
assign a27740 = ~a27738 & ~l1552;
assign a27742 = a14904 & a14892;
assign a27744 = a13522 & a13090;
assign a27746 = ~a27744 & ~a14910;
assign a27748 = a27746 & a14918;
assign a27750 = a27748 & a27742;
assign a27752 = ~a14908 & ~a14906;
assign a27754 = a27752 & a14898;
assign a27756 = ~a14934 & ~a14912;
assign a27758 = a27756 & a14942;
assign a27760 = a27758 & a27754;
assign a27762 = a27760 & a27750;
assign a27764 = ~a27762 & a13508;
assign a27766 = ~a27764 & ~a27740;
assign a27770 = a27768 & a11750;
assign a27772 = ~a27770 & ~a27736;
assign a27774 = a27772 & ~a27702;
assign a27776 = ~a27774 & a11630;
assign a27778 = ~a27776 & ~a27672;
assign a27780 = ~a27778 & ~a11624;
assign a27782 = a27562 & a27556;
assign a27784 = a27782 & a27538;
assign a27786 = ~a27784 & ~l1100;
assign a27788 = ~a27786 & ~a1690;
assign a27792 = a27790 & ~a11750;
assign a27794 = a27578 & a27562;
assign a27796 = a27794 & a27538;
assign a27798 = ~a27796 & ~l1098;
assign a27800 = ~a27798 & ~a1690;
assign a27804 = a27802 & a11750;
assign a27806 = ~a27804 & ~a27792;
assign a27808 = a13508 & l1100;
assign a27810 = ~a27808 & ~l1550;
assign a27812 = a15234 & a15222;
assign a27814 = a13522 & a13102;
assign a27816 = ~a27814 & ~a15240;
assign a27818 = a27816 & a15248;
assign a27820 = a27818 & a27812;
assign a27822 = ~a15238 & ~a15236;
assign a27824 = a27822 & a15228;
assign a27826 = ~a15264 & ~a15242;
assign a27828 = a27826 & a15272;
assign a27830 = a27828 & a27824;
assign a27832 = a27830 & a27820;
assign a27834 = ~a27832 & a13508;
assign a27836 = ~a27834 & ~a27810;
assign a27840 = a27838 & ~a11750;
assign a27842 = a13508 & l1098;
assign a27844 = ~a27842 & ~l1548;
assign a27846 = a13900 & a13888;
assign a27848 = a13522 & a13106;
assign a27850 = ~a27848 & ~a13906;
assign a27852 = a27850 & a13914;
assign a27854 = a27852 & a27846;
assign a27856 = ~a13904 & ~a13902;
assign a27858 = a27856 & a13894;
assign a27860 = ~a13930 & ~a13908;
assign a27862 = a27860 & a13938;
assign a27864 = a27862 & a27858;
assign a27866 = a27864 & a27854;
assign a27868 = ~a27866 & a13508;
assign a27870 = ~a27868 & ~a27844;
assign a27874 = a27872 & a11750;
assign a27876 = ~a27874 & ~a27840;
assign a27878 = a27876 & ~a27806;
assign a27880 = ~a27878 & ~a11630;
assign a27882 = a27674 & a27562;
assign a27884 = a27882 & a27538;
assign a27886 = ~a27884 & ~l1096;
assign a27888 = ~a27886 & ~a1690;
assign a27892 = a27890 & ~a11750;
assign a27894 = a27688 & a27562;
assign a27896 = a27894 & a27538;
assign a27898 = ~a27896 & ~l1094;
assign a27900 = ~a27898 & ~a1690;
assign a27904 = a27902 & a11750;
assign a27906 = ~a27904 & ~a27892;
assign a27908 = a13508 & l1096;
assign a27910 = ~a27908 & ~l1546;
assign a27912 = a15070 & a15058;
assign a27914 = a13522 & a13114;
assign a27916 = ~a27914 & ~a15076;
assign a27918 = a27916 & a15084;
assign a27920 = a27918 & a27912;
assign a27922 = ~a15074 & ~a15072;
assign a27924 = a27922 & a15064;
assign a27926 = ~a15100 & ~a15078;
assign a27928 = a27926 & a15108;
assign a27930 = a27928 & a27924;
assign a27932 = a27930 & a27920;
assign a27934 = ~a27932 & a13508;
assign a27936 = ~a27934 & ~a27910;
assign a27940 = a27938 & ~a11750;
assign a27942 = a13508 & l1094;
assign a27944 = ~a27942 & ~l1544;
assign a27946 = a13734 & a13722;
assign a27948 = a13522 & a13118;
assign a27950 = ~a27948 & ~a13740;
assign a27952 = a27950 & a13748;
assign a27954 = a27952 & a27946;
assign a27956 = ~a13738 & ~a13736;
assign a27958 = a27956 & a13728;
assign a27960 = ~a13764 & ~a13742;
assign a27962 = a27960 & a13772;
assign a27964 = a27962 & a27958;
assign a27966 = a27964 & a27954;
assign a27968 = ~a27966 & a13508;
assign a27970 = ~a27968 & ~a27944;
assign a27974 = a27972 & a11750;
assign a27976 = ~a27974 & ~a27940;
assign a27978 = a27976 & ~a27906;
assign a27980 = ~a27978 & a11630;
assign a27982 = ~a27980 & ~a27880;
assign a27984 = ~a27982 & a11624;
assign a27986 = ~a27984 & ~a27780;
assign a27988 = ~a27986 & ~a11622;
assign a27990 = ~a27562 & a27552;
assign a27992 = a27990 & a8866;
assign a27994 = a27992 & a27546;
assign a27996 = a27994 & a27538;
assign a27998 = ~a27996 & ~l1086;
assign a28000 = ~a27998 & ~l494;
assign a28002 = a28000 & ~a1690;
assign a28006 = ~a14406 & ~a14404;
assign a28008 = a28006 & ~a14402;
assign a28010 = a28008 & ~a14400;
assign a28012 = a28010 & ~a14398;
assign a28014 = a28012 & ~a14396;
assign a28016 = a28014 & ~a14394;
assign a28018 = a28016 & ~a14392;
assign a28020 = a28018 & ~a14390;
assign a28022 = a28020 & ~a14388;
assign a28024 = a28022 & ~a14386;
assign a28026 = a13522 & a13138;
assign a28028 = ~a28026 & a28024;
assign a28030 = a28028 & a14440;
assign a28032 = a28030 & a14412;
assign a28034 = a28032 & a14458;
assign a28036 = ~a28034 & ~l1542;
assign a28038 = a28036 & a28004;
assign a28040 = ~a28038 & a11750;
assign a28042 = a13508 & l1088;
assign a28044 = ~a28042 & ~l1540;
assign a28046 = a14236 & a14224;
assign a28048 = a13522 & a13134;
assign a28050 = ~a28048 & ~a14242;
assign a28052 = a28050 & a14250;
assign a28054 = a28052 & a28046;
assign a28056 = ~a14240 & ~a14238;
assign a28058 = a28056 & a14230;
assign a28060 = ~a14266 & ~a14244;
assign a28062 = a28060 & a14274;
assign a28064 = a28062 & a28058;
assign a28066 = a28064 & a28054;
assign a28068 = ~a28066 & a13508;
assign a28070 = ~a28068 & ~a28044;
assign a28074 = a27992 & ~a27546;
assign a28076 = a28074 & a27538;
assign a28078 = ~a28076 & ~l1088;
assign a28080 = ~a28078 & ~a1690;
assign a28084 = a28082 & ~a28072;
assign a28086 = ~a28084 & ~a11750;
assign a28088 = ~a28086 & ~a28040;
assign a28090 = ~a28088 & a11622;
assign a28092 = ~a28090 & ~a27988;
assign a28094 = ~a28092 & ~a27536;
assign a28096 = a28094 & a27506;
assign a28098 = a11750 & ~a5542;
assign a28100 = ~a11750 & ~a5548;
assign a28102 = ~a28100 & ~a28098;
assign a28104 = a11750 & ~a11630;
assign a28106 = ~a11750 & a11630;
assign a28108 = ~a28106 & ~a28104;
assign a28110 = a28108 & ~a28102;
assign a28112 = a28104 & ~a5556;
assign a28114 = a28106 & ~a5572;
assign a28116 = ~a28114 & ~a28112;
assign a28118 = a28116 & ~a28110;
assign a28120 = a11750 & a11630;
assign a28122 = ~a28120 & ~a11624;
assign a28124 = a28120 & a11624;
assign a28126 = ~a28124 & ~a28122;
assign a28128 = ~a28126 & ~a28118;
assign a28130 = a11750 & l576;
assign a28132 = ~a11750 & l578;
assign a28134 = ~a28132 & ~a28130;
assign a28136 = ~a28134 & a28108;
assign a28138 = a28104 & l580;
assign a28140 = a28106 & l582;
assign a28142 = ~a28140 & ~a28138;
assign a28144 = a28142 & ~a28136;
assign a28146 = ~a28144 & a28126;
assign a28148 = ~a28146 & ~a28128;
assign a28150 = a28124 & ~a11622;
assign a28152 = ~a28124 & a11622;
assign a28154 = ~a28152 & ~a28150;
assign a28156 = a28154 & ~a28148;
assign a28158 = a11750 & l586;
assign a28160 = ~a11750 & l584;
assign a28162 = ~a28160 & ~a28158;
assign a28164 = ~a28162 & ~a28154;
assign a28166 = ~a28164 & ~a28156;
assign a28168 = a16548 & a11750;
assign a28170 = ~a16548 & ~a11750;
assign a28172 = ~a28170 & ~a28168;
assign a28174 = a28108 & a16544;
assign a28176 = ~a28174 & a28172;
assign a28178 = ~a28126 & a16554;
assign a28180 = ~a28178 & a28176;
assign a28182 = a28154 & a16570;
assign a28184 = ~a28182 & a28180;
assign a28186 = ~a28108 & ~a16544;
assign a28188 = a28126 & ~a16554;
assign a28190 = ~a28188 & ~a28186;
assign a28192 = ~a28154 & ~a16570;
assign a28194 = ~a28192 & a28190;
assign a28196 = a28194 & a28184;
assign a28198 = ~a28196 & ~a28166;
assign a28200 = a28104 & a11830;
assign a28202 = ~a28200 & a28198;
assign a28204 = a28202 & a28094;
assign a28206 = ~a28204 & ~a28096;
assign a28208 = a28206 & a11622;
assign a28210 = a28204 & ~a28154;
assign a28212 = ~a28210 & ~a28208;
assign a28214 = ~a28212 & ~a6950;
assign a28216 = ~a16334 & a6950;
assign a28218 = ~a28216 & ~a28214;
assign a28220 = ~a28218 & ~a1690;
assign a28222 = ~a28220 & ~a6478;
assign a28224 = ~a28222 & ~l494;
assign a28226 = l1686 & ~l1538;
assign a28228 = a28226 & l494;
assign a28232 = a28206 & a11750;
assign a28234 = a28204 & ~a11750;
assign a28236 = ~a28234 & ~a28232;
assign a28238 = ~a28236 & ~a6950;
assign a28240 = ~a16340 & a6950;
assign a28242 = ~a28240 & ~a28238;
assign a28244 = ~a28242 & ~a1690;
assign a28246 = ~a28244 & ~a6514;
assign a28248 = ~a28246 & ~l494;
assign a28250 = l1686 & ~l1532;
assign a28252 = a28250 & l494;
assign a28256 = a28206 & a11624;
assign a28258 = a28204 & a28126;
assign a28260 = ~a28258 & ~a28256;
assign a28262 = ~a28260 & ~a6950;
assign a28264 = ~a16326 & a6950;
assign a28266 = ~a28264 & ~a28262;
assign a28268 = ~a28266 & ~a1690;
assign a28270 = ~a28268 & ~a6594;
assign a28272 = ~a28270 & ~l494;
assign a28274 = l1686 & ~l1534;
assign a28276 = a28274 & l494;
assign a28280 = a28206 & a11630;
assign a28282 = a28204 & ~a28108;
assign a28284 = ~a28282 & ~a28280;
assign a28286 = ~a28284 & ~a6950;
assign a28288 = ~a16320 & a6950;
assign a28290 = ~a28288 & ~a28286;
assign a28292 = ~a28290 & ~a1690;
assign a28294 = ~a28292 & ~a6550;
assign a28296 = ~a28294 & ~l494;
assign a28298 = l1686 & ~l1536;
assign a28300 = a28298 & l494;
assign a28304 = ~a27994 & a13316;
assign a28306 = ~a25758 & i414;
assign a28308 = a25758 & ~a13332;
assign a28310 = ~a28308 & ~a28306;
assign a28312 = a28310 & a27994;
assign a28316 = ~a28074 & a13312;
assign a28318 = a28310 & a28074;
assign a28322 = ~a27894 & a13296;
assign a28324 = a28310 & a27894;
assign a28328 = ~a27882 & a13292;
assign a28330 = a28310 & a27882;
assign a28334 = ~a27794 & a13284;
assign a28336 = a28310 & a27794;
assign a28340 = ~a27782 & a13280;
assign a28342 = a28310 & a27782;
assign a28346 = ~a27690 & a13268;
assign a28348 = a28310 & a27690;
assign a28352 = ~a27676 & a13264;
assign a28354 = a28310 & a27676;
assign a28358 = ~a27580 & a13256;
assign a28360 = a28310 & a27580;
assign a28364 = ~a27564 & a13252;
assign a28366 = a28310 & a27564;
assign a28370 = ~a27994 & a13138;
assign a28372 = ~a25758 & i412;
assign a28374 = a25758 & a13158;
assign a28376 = ~a28374 & ~a28372;
assign a28378 = a28376 & a27994;
assign a28382 = ~a28074 & a13134;
assign a28384 = a28376 & a28074;
assign a28388 = ~a27894 & a13118;
assign a28390 = a28376 & a27894;
assign a28394 = ~a27882 & a13114;
assign a28396 = a28376 & a27882;
assign a28400 = ~a27794 & a13106;
assign a28402 = a28376 & a27794;
assign a28406 = ~a27782 & a13102;
assign a28408 = a28376 & a27782;
assign a28412 = ~a27690 & a13090;
assign a28414 = a28376 & a27690;
assign a28418 = ~a27676 & a13086;
assign a28420 = a28376 & a27676;
assign a28424 = ~a27580 & a13078;
assign a28426 = a28376 & a27580;
assign a28430 = ~a27564 & a13068;
assign a28432 = a28376 & a27564;
assign a28436 = ~a27994 & a12966;
assign a28438 = ~a25758 & i410;
assign a28440 = a25758 & a12986;
assign a28442 = ~a28440 & ~a28438;
assign a28444 = a28442 & a27994;
assign a28448 = ~a28074 & a12962;
assign a28450 = a28442 & a28074;
assign a28454 = ~a27894 & a12946;
assign a28456 = a28442 & a27894;
assign a28460 = ~a27882 & a12942;
assign a28462 = a28442 & a27882;
assign a28466 = ~a27794 & a12934;
assign a28468 = a28442 & a27794;
assign a28472 = ~a27782 & a12930;
assign a28474 = a28442 & a27782;
assign a28478 = ~a27690 & a12918;
assign a28480 = a28442 & a27690;
assign a28484 = ~a27676 & a12914;
assign a28486 = a28442 & a27676;
assign a28490 = ~a27580 & a12906;
assign a28492 = a28442 & a27580;
assign a28496 = ~a27564 & a12896;
assign a28498 = a28442 & a27564;
assign a28502 = ~a27994 & a12766;
assign a28504 = ~a25758 & i408;
assign a28506 = a25758 & a12786;
assign a28508 = ~a28506 & ~a28504;
assign a28510 = a28508 & a27994;
assign a28514 = ~a28074 & a12762;
assign a28516 = a28508 & a28074;
assign a28520 = ~a27894 & a12746;
assign a28522 = a28508 & a27894;
assign a28526 = ~a27882 & a12742;
assign a28528 = a28508 & a27882;
assign a28532 = ~a27794 & a12734;
assign a28534 = a28508 & a27794;
assign a28538 = ~a27782 & a12730;
assign a28540 = a28508 & a27782;
assign a28544 = ~a27690 & a12718;
assign a28546 = a28508 & a27690;
assign a28550 = ~a27676 & a12714;
assign a28552 = a28508 & a27676;
assign a28556 = ~a27580 & a12706;
assign a28558 = a28508 & a27580;
assign a28562 = ~a27564 & a12696;
assign a28564 = a28508 & a27564;
assign a28568 = ~a27994 & a12566;
assign a28570 = ~a25758 & i406;
assign a28572 = a25758 & a12586;
assign a28574 = ~a28572 & ~a28570;
assign a28576 = a28574 & a27994;
assign a28580 = ~a28074 & a12562;
assign a28582 = a28574 & a28074;
assign a28586 = ~a27894 & a12546;
assign a28588 = a28574 & a27894;
assign a28592 = ~a27882 & a12542;
assign a28594 = a28574 & a27882;
assign a28598 = ~a27794 & a12534;
assign a28600 = a28574 & a27794;
assign a28604 = ~a27782 & a12530;
assign a28606 = a28574 & a27782;
assign a28610 = ~a27690 & a12518;
assign a28612 = a28574 & a27690;
assign a28616 = ~a27676 & a12514;
assign a28618 = a28574 & a27676;
assign a28622 = ~a27580 & a12506;
assign a28624 = a28574 & a27580;
assign a28628 = ~a27564 & a12496;
assign a28630 = a28574 & a27564;
assign a28634 = ~a27994 & a12366;
assign a28636 = ~a25758 & i404;
assign a28638 = a25758 & a12386;
assign a28640 = ~a28638 & ~a28636;
assign a28642 = a28640 & a27994;
assign a28646 = ~a28074 & a12362;
assign a28648 = a28640 & a28074;
assign a28652 = ~a27894 & a12346;
assign a28654 = a28640 & a27894;
assign a28658 = ~a27882 & a12342;
assign a28660 = a28640 & a27882;
assign a28664 = ~a27794 & a12334;
assign a28666 = a28640 & a27794;
assign a28670 = ~a27782 & a12330;
assign a28672 = a28640 & a27782;
assign a28676 = ~a27690 & a12318;
assign a28678 = a28640 & a27690;
assign a28682 = ~a27676 & a12314;
assign a28684 = a28640 & a27676;
assign a28688 = ~a27580 & a12306;
assign a28690 = a28640 & a27580;
assign a28694 = ~a27564 & a12296;
assign a28696 = a28640 & a27564;
assign a28700 = ~a27994 & a12166;
assign a28702 = ~a25758 & i402;
assign a28704 = a25758 & a12186;
assign a28706 = ~a28704 & ~a28702;
assign a28708 = a28706 & a27994;
assign a28712 = ~a28074 & a12162;
assign a28714 = a28706 & a28074;
assign a28718 = ~a27894 & a12146;
assign a28720 = a28706 & a27894;
assign a28724 = ~a27882 & a12142;
assign a28726 = a28706 & a27882;
assign a28730 = ~a27794 & a12134;
assign a28732 = a28706 & a27794;
assign a28736 = ~a27782 & a12130;
assign a28738 = a28706 & a27782;
assign a28742 = ~a27690 & a12118;
assign a28744 = a28706 & a27690;
assign a28748 = ~a27676 & a12114;
assign a28750 = a28706 & a27676;
assign a28754 = ~a27580 & a12106;
assign a28756 = a28706 & a27580;
assign a28760 = ~a27564 & a12096;
assign a28762 = a28706 & a27564;
assign a28766 = ~a27994 & a11970;
assign a28768 = ~a25758 & i368;
assign a28770 = a25758 & ~a11998;
assign a28772 = ~a28770 & ~a28768;
assign a28774 = a28772 & a27994;
assign a28778 = ~a28074 & a11966;
assign a28780 = a28772 & a28074;
assign a28784 = ~a27894 & a11950;
assign a28786 = a28772 & a27894;
assign a28790 = ~a27882 & a11946;
assign a28792 = a28772 & a27882;
assign a28796 = ~a27794 & a11938;
assign a28798 = a28772 & a27794;
assign a28802 = ~a27782 & a11934;
assign a28804 = a28772 & a27782;
assign a28808 = ~a27690 & a11922;
assign a28810 = a28772 & a27690;
assign a28814 = ~a27676 & a11918;
assign a28816 = a28772 & a27676;
assign a28820 = ~a27580 & a11910;
assign a28822 = a28772 & a27580;
assign a28826 = ~a27564 & a11906;
assign a28828 = a28772 & a27564;
assign a28832 = a13494 & a11426;
assign a28836 = a13708 & ~a6934;
assign a28838 = ~a28836 & ~a16342;
assign a28840 = a28838 & ~a1690;
assign a28842 = ~a28840 & ~a6514;
assign a28844 = ~a16652 & a1690;
assign a28846 = a28844 & ~a17864;
assign a28848 = a13710 & ~a6934;
assign a28850 = ~a28848 & ~a17478;
assign a28852 = a28850 & ~a1690;
assign a28854 = ~a28852 & ~a28846;
assign a28856 = a13696 & ~a6934;
assign a28858 = ~a28856 & ~a16938;
assign a28860 = ~a28858 & ~a1690;
assign a28862 = ~a17198 & ~a16650;
assign a28864 = ~a28862 & a28844;
assign a28868 = a13702 & ~a6934;
assign a28870 = ~a28868 & ~a16664;
assign a28872 = ~a28870 & ~a1690;
assign a28874 = ~a16926 & ~a16648;
assign a28876 = ~a28874 & a28844;
assign a28880 = ~a27492 & ~a24508;
assign a28884 = ~a22654 & a15350;
assign a28886 = a22654 & a10178;
assign a28890 = ~a22654 & a15384;
assign a28892 = a22654 & a10152;
assign a28896 = ~a22654 & a15488;
assign a28898 = a22654 & a10126;
assign a28902 = ~a22654 & a15592;
assign a28904 = a22654 & a10100;
assign a28908 = ~a22654 & a15696;
assign a28910 = a22654 & a10074;
assign a28914 = ~a22654 & a15794;
assign a28916 = a22654 & a10044;
assign a28920 = ~a22654 & a15892;
assign a28922 = a22654 & a8874;
assign a28926 = ~a8850 & ~l1686;
assign a28928 = l1686 & l1502;
assign a28930 = ~a28928 & ~a28926;
assign a28932 = ~a28930 & a25742;
assign a28934 = a28932 & ~l664;
assign a28936 = ~a25752 & ~i396;
assign a28940 = ~i394 & i392;
assign a28944 = ~a27414 & ~a8860;
assign a28946 = a27398 & a8862;
assign a28948 = ~a28946 & ~a28944;
assign a28950 = ~a27398 & ~a8862;
assign a28952 = a27414 & a8860;
assign a28954 = ~a28952 & ~a28950;
assign a28956 = a28954 & a28948;
assign a28958 = a27430 & a10706;
assign a28960 = a27060 & a8866;
assign a28962 = ~a28960 & ~a28958;
assign a28964 = a28962 & a28956;
assign a28966 = ~a27430 & ~a10706;
assign a28968 = ~a27060 & ~a8866;
assign a28970 = ~a28968 & ~a28966;
assign a28974 = ~a16548 & l586;
assign a28976 = a16548 & l584;
assign a28978 = ~a28976 & ~a28974;
assign a28980 = ~a28978 & a16570;
assign a28982 = ~a28980 & ~a5580;
assign a28984 = ~a16548 & ~a5542;
assign a28986 = a16548 & ~a5548;
assign a28988 = ~a28986 & ~a28984;
assign a28990 = ~a28988 & ~a16544;
assign a28992 = ~a16548 & ~a5556;
assign a28994 = a16548 & ~a5572;
assign a28996 = ~a28994 & ~a28992;
assign a28998 = ~a28996 & a16544;
assign a29000 = ~a28998 & ~a28990;
assign a29002 = ~a29000 & ~a16554;
assign a29004 = ~a16548 & l576;
assign a29006 = a16548 & l578;
assign a29008 = ~a29006 & ~a29004;
assign a29010 = ~a29008 & ~a16544;
assign a29012 = ~a16548 & l580;
assign a29014 = a16548 & l582;
assign a29016 = ~a29014 & ~a29012;
assign a29018 = ~a29016 & a16544;
assign a29020 = ~a29018 & ~a29010;
assign a29022 = ~a29020 & a16554;
assign a29024 = ~a29022 & ~a29002;
assign a29026 = ~a29024 & ~a16570;
assign a29028 = ~a29026 & a28982;
assign a29030 = ~a29028 & a16570;
assign a29032 = a16548 & a16544;
assign a29034 = a29032 & a16554;
assign a29036 = a29034 & ~a16570;
assign a29038 = ~a29034 & a16570;
assign a29040 = ~a29038 & ~a29036;
assign a29042 = a16548 & l1508;
assign a29044 = a29042 & a16570;
assign a29046 = a29044 & ~a16554;
assign a29048 = ~a29046 & a29028;
assign a29050 = a29048 & ~a29040;
assign a29052 = ~a29050 & ~a29030;
assign a29054 = ~a29052 & ~l664;
assign a29056 = a28226 & l664;
assign a29060 = a29048 & a16548;
assign a29062 = ~a29060 & ~a16544;
assign a29064 = a29048 & a29032;
assign a29066 = ~a29064 & ~a29062;
assign a29068 = a29066 & ~l664;
assign a29070 = a28298 & l664;
assign a29074 = ~a29064 & a16554;
assign a29076 = a29064 & ~a16554;
assign a29078 = ~a29076 & ~a29074;
assign a29080 = ~a29078 & ~l664;
assign a29082 = a28274 & l664;
assign a29086 = ~a29028 & a16548;
assign a29088 = a29048 & ~a16548;
assign a29090 = ~a29088 & ~a29086;
assign a29092 = ~a29090 & ~l664;
assign a29094 = a28250 & l664;
assign a29098 = a28250 & ~a6682;
assign a29100 = a6682 & ~a5124;
assign a29104 = a28274 & ~a6682;
assign a29106 = a6682 & ~a6604;
assign a29110 = a28298 & ~a6682;
assign a29112 = a6682 & ~a6562;
assign a29116 = a28226 & ~a6682;
assign a29118 = a6682 & ~a6490;
assign a29124 = ~a15296 & a11416;
assign a29126 = a29124 & a6934;
assign a29128 = ~a29126 & a27434;
assign a29130 = ~a29128 & ~l494;
assign a29134 = a6666 & i468;
assign a29136 = a29134 & ~l1686;
assign a29138 = l1686 & l1568;
assign a29140 = ~a29138 & ~a29136;
assign a29142 = a21812 & a20890;
assign a29146 = a6666 & i470;
assign a29148 = a29146 & ~l1686;
assign a29150 = l1686 & l1570;
assign a29152 = ~a29150 & ~a29148;
assign a29156 = a20890 & i472;
assign a29158 = a29156 & a6674;
assign a29162 = a19386 & ~a6950;
assign a29164 = ~a19494 & a6950;
assign a29166 = ~a29164 & ~a29162;
assign a29168 = ~a29166 & ~a6906;
assign a29172 = a19382 & ~a6950;
assign a29174 = ~a19484 & a6950;
assign a29176 = ~a29174 & ~a29172;
assign a29178 = ~a29176 & ~a6906;
assign a29182 = a19378 & ~a6950;
assign a29184 = ~a19474 & a6950;
assign a29186 = ~a29184 & ~a29182;
assign a29188 = ~a29186 & ~a6906;
assign a29192 = a19376 & ~a6950;
assign a29194 = ~a19510 & a6950;
assign a29196 = ~a29194 & ~a29192;
assign a29198 = ~a29196 & ~a6906;
assign a29202 = a19374 & ~a6950;
assign a29204 = ~a19518 & a6950;
assign a29206 = ~a29204 & ~a29202;
assign a29208 = ~a29206 & ~a6906;
assign a29212 = a19372 & ~a6950;
assign a29214 = ~a19526 & a6950;
assign a29216 = ~a29214 & ~a29212;
assign a29218 = ~a29216 & ~a6906;
assign a29222 = a19370 & ~a6950;
assign a29224 = ~a19534 & a6950;
assign a29226 = ~a29224 & ~a29222;
assign a29228 = ~a29226 & ~a6906;
assign a29232 = a19864 & ~a6950;
assign a29234 = ~a19886 & a6950;
assign a29236 = ~a29234 & ~a29232;
assign a29238 = ~a29236 & ~a6906;
assign a29242 = l1686 & ~l1602;
assign a29244 = l1686 & ~l1612;
assign a29246 = ~a6604 & l1604;
assign a29250 = l1686 & ~l1610;
assign a29252 = ~a6490 & l1604;
assign a29256 = a29254 & a29248;
assign a29258 = l1686 & ~l1608;
assign a29260 = ~a6562 & l1604;
assign a29264 = ~a29262 & a29256;
assign a29266 = l1686 & ~l1606;
assign a29268 = ~a5124 & l1604;
assign a29272 = ~a29270 & a29264;
assign a29274 = a29272 & a17976;
assign a29276 = a29262 & a29248;
assign a29278 = a29276 & ~a29254;
assign a29280 = a29278 & ~a29270;
assign a29282 = a29280 & a17992;
assign a29284 = ~a29282 & ~a29274;
assign a29286 = a29254 & ~a29248;
assign a29288 = a29286 & a29262;
assign a29290 = a29288 & a29270;
assign a29292 = a29290 & a17926;
assign a29294 = a29286 & ~a29262;
assign a29296 = a29294 & a29270;
assign a29298 = a29296 & a17956;
assign a29300 = ~a29298 & ~a29292;
assign a29302 = a29300 & a29284;
assign a29304 = a29262 & a29256;
assign a29306 = a29304 & ~a29270;
assign a29308 = a29306 & a18004;
assign a29310 = a29278 & a29270;
assign a29312 = a29310 & a17934;
assign a29314 = ~a29312 & ~a29308;
assign a29316 = a29314 & a29302;
assign a29318 = a29270 & a29264;
assign a29320 = a29318 & a18012;
assign a29322 = a29294 & ~a29270;
assign a29324 = a29322 & a17944;
assign a29326 = ~a29324 & ~a29320;
assign a29328 = a29304 & a29270;
assign a29330 = a29328 & a17962;
assign a29332 = a29288 & ~a29270;
assign a29334 = a29332 & a17986;
assign a29336 = ~a29334 & ~a29330;
assign a29338 = a29336 & a29326;
assign a29342 = l1686 & ~l1644;
assign a29344 = ~a29248 & ~a19224;
assign a29346 = a29248 & a19224;
assign a29348 = ~a29346 & ~a29344;
assign a29350 = ~a29254 & ~a19218;
assign a29352 = a29254 & a19218;
assign a29354 = ~a29352 & ~a29350;
assign a29356 = a29354 & a29348;
assign a29358 = a29270 & a19232;
assign a29360 = ~a29270 & ~a19232;
assign a29362 = ~a29360 & ~a29358;
assign a29364 = a29262 & a19222;
assign a29366 = ~a29364 & a29362;
assign a29368 = ~a29262 & ~a19222;
assign a29370 = ~a29368 & a29366;
assign a29372 = a29370 & a29356;
assign a29374 = ~a29372 & l1614;
assign a29376 = ~a27436 & ~l664;
assign a29378 = a29376 & a29374;
assign a29380 = a29378 & a29270;
assign a29382 = ~a29380 & ~a29342;
assign a29384 = ~a29374 & ~l1496;
assign a29386 = a29384 & a29376;
assign a29388 = a29386 & ~a29270;
assign a29392 = l1686 & ~l1640;
assign a29394 = ~a29270 & a29262;
assign a29396 = a29394 & a29254;
assign a29398 = a29270 & ~a29262;
assign a29400 = ~a29398 & ~a29396;
assign a29402 = ~a29400 & a29378;
assign a29404 = ~a29402 & ~a29392;
assign a29406 = a29386 & ~a29262;
assign a29410 = l1686 & ~l1632;
assign a29412 = a29270 & ~a29254;
assign a29414 = ~a29270 & ~a29262;
assign a29416 = a29414 & ~a29248;
assign a29418 = ~a29416 & ~a29412;
assign a29420 = ~a29418 & a29378;
assign a29422 = ~a29420 & ~a29410;
assign a29424 = a29386 & ~a29254;
assign a29428 = l1686 & ~l1616;
assign a29430 = ~a29414 & a29248;
assign a29432 = ~a29430 & ~a29416;
assign a29434 = a29432 & a29378;
assign a29436 = ~a29434 & ~a29428;
assign a29438 = a29386 & ~a29248;
assign a29442 = a29272 & l910;
assign a29444 = a29280 & ~a18104;
assign a29446 = ~a29444 & ~a29442;
assign a29448 = a29290 & l912;
assign a29450 = a29294 & a18144;
assign a29452 = a29450 & a29270;
assign a29454 = ~a29452 & ~a29448;
assign a29456 = a29454 & a29446;
assign a29458 = a29306 & l904;
assign a29460 = a29278 & ~a18136;
assign a29462 = a29460 & a29270;
assign a29464 = ~a29462 & ~a29458;
assign a29466 = a29464 & a29456;
assign a29468 = a29264 & l916;
assign a29470 = a29468 & a29270;
assign a29472 = a29322 & l906;
assign a29474 = ~a29472 & ~a29470;
assign a29476 = a29328 & ~a18126;
assign a29478 = a29332 & l902;
assign a29480 = ~a29478 & ~a29476;
assign a29482 = a29480 & a29474;
assign a29484 = a29482 & a29466;
assign a29486 = ~a29484 & a29374;
assign a29488 = ~a29468 & ~a29460;
assign a29490 = ~a29488 & ~a29270;
assign a29492 = a29290 & l910;
assign a29494 = a29296 & l902;
assign a29496 = ~a29494 & ~a29492;
assign a29498 = a29496 & ~a29490;
assign a29500 = a29306 & ~a18126;
assign a29502 = a29310 & l906;
assign a29504 = ~a29502 & ~a29500;
assign a29506 = a29504 & a29498;
assign a29508 = a29318 & l904;
assign a29510 = a29450 & ~a29270;
assign a29512 = ~a29510 & ~a29508;
assign a29514 = a29328 & ~a18104;
assign a29516 = a29332 & l912;
assign a29518 = ~a29516 & ~a29514;
assign a29520 = a29518 & a29512;
assign a29522 = a29520 & a29506;
assign a29524 = ~a29522 & ~a29374;
assign a29526 = ~a29524 & ~a29486;
assign a29528 = a29328 & a18246;
assign a29530 = a29280 & a18212;
assign a29532 = ~a29530 & ~a29528;
assign a29534 = a29278 & a18218;
assign a29536 = a29294 & a18204;
assign a29538 = ~a29536 & ~a29534;
assign a29540 = ~a29538 & a29270;
assign a29542 = ~a29540 & a29532;
assign a29544 = a29290 & a18224;
assign a29546 = a29332 & a18232;
assign a29548 = ~a29546 & ~a29544;
assign a29550 = a29548 & a29542;
assign a29552 = a29322 & a18200;
assign a29554 = a29264 & a18252;
assign a29556 = a29554 & a29270;
assign a29558 = ~a29556 & ~a29552;
assign a29560 = a29256 & a18256;
assign a29562 = a29560 & a29394;
assign a29564 = a29272 & a18236;
assign a29566 = ~a29564 & ~a29562;
assign a29568 = a29566 & a29558;
assign a29570 = a29568 & a29550;
assign a29572 = ~a29570 & a29374;
assign a29574 = ~a29554 & ~a29534;
assign a29576 = ~a29574 & ~a29270;
assign a29578 = a29254 & a18236;
assign a29580 = a29262 & ~a29248;
assign a29582 = a29580 & a29270;
assign a29584 = a29582 & a29578;
assign a29586 = ~a29584 & ~a29576;
assign a29588 = a29536 & ~a29270;
assign a29590 = a29276 & a18212;
assign a29592 = a29270 & a29254;
assign a29594 = a29592 & a29590;
assign a29596 = a29560 & a29398;
assign a29598 = ~a29596 & ~a29594;
assign a29600 = a29598 & ~a29588;
assign a29602 = a29600 & a29586;
assign a29604 = a29332 & a18224;
assign a29606 = a29306 & a18246;
assign a29608 = ~a29606 & ~a29604;
assign a29610 = a29296 & a18232;
assign a29612 = a29310 & a18200;
assign a29614 = ~a29612 & ~a29610;
assign a29616 = a29614 & a29608;
assign a29618 = a29616 & a29602;
assign a29620 = ~a29618 & ~a29374;
assign a29622 = ~a29620 & ~a29572;
assign a29624 = ~a29622 & a22006;
assign a29626 = ~a29624 & ~a29526;
assign a29628 = a29622 & ~a22006;
assign a29630 = ~a29628 & a29626;
assign a29632 = a29328 & a18366;
assign a29634 = a29280 & a18328;
assign a29636 = ~a29634 & ~a29632;
assign a29638 = a29278 & a18334;
assign a29640 = a29294 & a18320;
assign a29642 = ~a29640 & ~a29638;
assign a29644 = ~a29642 & a29270;
assign a29646 = ~a29644 & a29636;
assign a29648 = a29290 & a18340;
assign a29650 = a29332 & a18348;
assign a29652 = ~a29650 & ~a29648;
assign a29654 = a29652 & a29646;
assign a29656 = a29322 & a18316;
assign a29658 = a29264 & a18372;
assign a29660 = a29658 & a29270;
assign a29662 = ~a29660 & ~a29656;
assign a29664 = a29256 & a18376;
assign a29666 = a29664 & a29394;
assign a29668 = a29272 & a18352;
assign a29670 = ~a29668 & ~a29666;
assign a29672 = a29670 & a29662;
assign a29674 = a29672 & a29654;
assign a29676 = ~a29674 & a29374;
assign a29678 = ~a29658 & ~a29638;
assign a29680 = ~a29678 & ~a29270;
assign a29682 = a29254 & a18352;
assign a29684 = a29682 & a29582;
assign a29686 = ~a29684 & ~a29680;
assign a29688 = a29640 & ~a29270;
assign a29690 = a29276 & a18328;
assign a29692 = a29690 & a29592;
assign a29694 = a29664 & a29398;
assign a29696 = ~a29694 & ~a29692;
assign a29698 = a29696 & ~a29688;
assign a29700 = a29698 & a29686;
assign a29702 = a29332 & a18340;
assign a29704 = a29306 & a18366;
assign a29706 = ~a29704 & ~a29702;
assign a29708 = a29296 & a18348;
assign a29710 = a29310 & a18316;
assign a29712 = ~a29710 & ~a29708;
assign a29714 = a29712 & a29706;
assign a29716 = a29714 & a29700;
assign a29718 = ~a29716 & ~a29374;
assign a29720 = ~a29718 & ~a29676;
assign a29722 = ~a29720 & a21872;
assign a29724 = ~a29722 & a29630;
assign a29726 = a29720 & ~a21872;
assign a29728 = ~a29726 & a29724;
assign a29730 = a29328 & a19100;
assign a29732 = a29280 & a19062;
assign a29734 = ~a29732 & ~a29730;
assign a29736 = a29278 & a19068;
assign a29738 = a29294 & a19052;
assign a29740 = ~a29738 & ~a29736;
assign a29742 = ~a29740 & a29270;
assign a29744 = ~a29742 & a29734;
assign a29746 = a29290 & a19074;
assign a29748 = a29332 & a19082;
assign a29750 = ~a29748 & ~a29746;
assign a29752 = a29750 & a29744;
assign a29754 = a29322 & a19048;
assign a29756 = a29264 & a19106;
assign a29758 = a29756 & a29270;
assign a29760 = ~a29758 & ~a29754;
assign a29762 = a29256 & a19110;
assign a29764 = a29762 & a29394;
assign a29766 = a29272 & a19086;
assign a29768 = ~a29766 & ~a29764;
assign a29770 = a29768 & a29760;
assign a29772 = a29770 & a29752;
assign a29774 = ~a29772 & a29374;
assign a29776 = ~a29756 & ~a29736;
assign a29778 = ~a29776 & ~a29270;
assign a29780 = a29254 & a19086;
assign a29782 = a29780 & a29582;
assign a29784 = ~a29782 & ~a29778;
assign a29786 = a29738 & ~a29270;
assign a29788 = a29276 & a19062;
assign a29790 = a29788 & a29592;
assign a29792 = a29762 & a29398;
assign a29794 = ~a29792 & ~a29790;
assign a29796 = a29794 & ~a29786;
assign a29798 = a29796 & a29784;
assign a29800 = a29332 & a19074;
assign a29802 = a29306 & a19100;
assign a29804 = ~a29802 & ~a29800;
assign a29806 = a29296 & a19082;
assign a29808 = a29310 & a19048;
assign a29810 = ~a29808 & ~a29806;
assign a29812 = a29810 & a29804;
assign a29814 = a29812 & a29798;
assign a29816 = ~a29814 & ~a29374;
assign a29818 = ~a29816 & ~a29774;
assign a29820 = ~a29818 & a21888;
assign a29822 = ~a29820 & a29728;
assign a29824 = a29818 & ~a21888;
assign a29826 = ~a29824 & a29822;
assign a29828 = a29328 & a18976;
assign a29830 = a29280 & a18938;
assign a29832 = ~a29830 & ~a29828;
assign a29834 = a29278 & a18944;
assign a29836 = a29294 & a18928;
assign a29838 = ~a29836 & ~a29834;
assign a29840 = ~a29838 & a29270;
assign a29842 = ~a29840 & a29832;
assign a29844 = a29290 & a18950;
assign a29846 = a29332 & a18958;
assign a29848 = ~a29846 & ~a29844;
assign a29850 = a29848 & a29842;
assign a29852 = a29322 & a18924;
assign a29854 = a29264 & a18982;
assign a29856 = a29854 & a29270;
assign a29858 = ~a29856 & ~a29852;
assign a29860 = a29256 & a18986;
assign a29862 = a29860 & a29394;
assign a29864 = a29272 & a18962;
assign a29866 = ~a29864 & ~a29862;
assign a29868 = a29866 & a29858;
assign a29870 = a29868 & a29850;
assign a29872 = ~a29870 & a29374;
assign a29874 = ~a29854 & ~a29834;
assign a29876 = ~a29874 & ~a29270;
assign a29878 = a29254 & a18962;
assign a29880 = a29878 & a29582;
assign a29882 = ~a29880 & ~a29876;
assign a29884 = a29836 & ~a29270;
assign a29886 = a29276 & a18938;
assign a29888 = a29886 & a29592;
assign a29890 = a29860 & a29398;
assign a29892 = ~a29890 & ~a29888;
assign a29894 = a29892 & ~a29884;
assign a29896 = a29894 & a29882;
assign a29898 = a29332 & a18950;
assign a29900 = a29306 & a18976;
assign a29902 = ~a29900 & ~a29898;
assign a29904 = a29296 & a18958;
assign a29906 = a29310 & a18924;
assign a29908 = ~a29906 & ~a29904;
assign a29910 = a29908 & a29902;
assign a29912 = a29910 & a29896;
assign a29914 = ~a29912 & ~a29374;
assign a29916 = ~a29914 & ~a29872;
assign a29918 = ~a29916 & a21904;
assign a29920 = ~a29918 & a29826;
assign a29922 = a29916 & ~a21904;
assign a29924 = ~a29922 & a29920;
assign a29926 = a29328 & a18852;
assign a29928 = a29280 & a18814;
assign a29930 = ~a29928 & ~a29926;
assign a29932 = a29278 & a18820;
assign a29934 = a29294 & a18804;
assign a29936 = ~a29934 & ~a29932;
assign a29938 = ~a29936 & a29270;
assign a29940 = ~a29938 & a29930;
assign a29942 = a29290 & a18826;
assign a29944 = a29332 & a18834;
assign a29946 = ~a29944 & ~a29942;
assign a29948 = a29946 & a29940;
assign a29950 = a29322 & a18800;
assign a29952 = a29264 & a18858;
assign a29954 = a29952 & a29270;
assign a29956 = ~a29954 & ~a29950;
assign a29958 = a29256 & a18862;
assign a29960 = a29958 & a29394;
assign a29962 = a29272 & a18838;
assign a29964 = ~a29962 & ~a29960;
assign a29966 = a29964 & a29956;
assign a29968 = a29966 & a29948;
assign a29970 = ~a29968 & a29374;
assign a29972 = ~a29952 & ~a29932;
assign a29974 = ~a29972 & ~a29270;
assign a29976 = a29254 & a18838;
assign a29978 = a29976 & a29582;
assign a29980 = ~a29978 & ~a29974;
assign a29982 = a29934 & ~a29270;
assign a29984 = a29276 & a18814;
assign a29986 = a29984 & a29592;
assign a29988 = a29958 & a29398;
assign a29990 = ~a29988 & ~a29986;
assign a29992 = a29990 & ~a29982;
assign a29994 = a29992 & a29980;
assign a29996 = a29332 & a18826;
assign a29998 = a29306 & a18852;
assign a30000 = ~a29998 & ~a29996;
assign a30002 = a29296 & a18834;
assign a30004 = a29310 & a18800;
assign a30006 = ~a30004 & ~a30002;
assign a30008 = a30006 & a30000;
assign a30010 = a30008 & a29994;
assign a30012 = ~a30010 & ~a29374;
assign a30014 = ~a30012 & ~a29970;
assign a30016 = ~a30014 & a21920;
assign a30018 = ~a30016 & a29924;
assign a30020 = a30014 & ~a21920;
assign a30022 = ~a30020 & a30018;
assign a30024 = a29328 & a18728;
assign a30026 = a29280 & a18690;
assign a30028 = ~a30026 & ~a30024;
assign a30030 = a29278 & a18696;
assign a30032 = a29294 & a18680;
assign a30034 = ~a30032 & ~a30030;
assign a30036 = ~a30034 & a29270;
assign a30038 = ~a30036 & a30028;
assign a30040 = a29290 & a18702;
assign a30042 = a29332 & a18710;
assign a30044 = ~a30042 & ~a30040;
assign a30046 = a30044 & a30038;
assign a30048 = a29322 & a18676;
assign a30050 = a29264 & a18734;
assign a30052 = a30050 & a29270;
assign a30054 = ~a30052 & ~a30048;
assign a30056 = a29256 & a18738;
assign a30058 = a30056 & a29394;
assign a30060 = a29272 & a18714;
assign a30062 = ~a30060 & ~a30058;
assign a30064 = a30062 & a30054;
assign a30066 = a30064 & a30046;
assign a30068 = ~a30066 & a29374;
assign a30070 = ~a30050 & ~a30030;
assign a30072 = ~a30070 & ~a29270;
assign a30074 = a29254 & a18714;
assign a30076 = a30074 & a29582;
assign a30078 = ~a30076 & ~a30072;
assign a30080 = a30032 & ~a29270;
assign a30082 = a29276 & a18690;
assign a30084 = a30082 & a29592;
assign a30086 = a30056 & a29398;
assign a30088 = ~a30086 & ~a30084;
assign a30090 = a30088 & ~a30080;
assign a30092 = a30090 & a30078;
assign a30094 = a29332 & a18702;
assign a30096 = a29306 & a18728;
assign a30098 = ~a30096 & ~a30094;
assign a30100 = a29296 & a18710;
assign a30102 = a29310 & a18676;
assign a30104 = ~a30102 & ~a30100;
assign a30106 = a30104 & a30098;
assign a30108 = a30106 & a30092;
assign a30110 = ~a30108 & ~a29374;
assign a30112 = ~a30110 & ~a30068;
assign a30114 = ~a30112 & a21936;
assign a30116 = ~a30114 & a30022;
assign a30118 = a30112 & ~a21936;
assign a30120 = ~a30118 & a30116;
assign a30122 = a29328 & a18604;
assign a30124 = a29280 & a18566;
assign a30126 = ~a30124 & ~a30122;
assign a30128 = a29278 & a18572;
assign a30130 = a29294 & a18556;
assign a30132 = ~a30130 & ~a30128;
assign a30134 = ~a30132 & a29270;
assign a30136 = ~a30134 & a30126;
assign a30138 = a29290 & a18578;
assign a30140 = a29332 & a18586;
assign a30142 = ~a30140 & ~a30138;
assign a30144 = a30142 & a30136;
assign a30146 = a29322 & a18552;
assign a30148 = a29264 & a18610;
assign a30150 = a30148 & a29270;
assign a30152 = ~a30150 & ~a30146;
assign a30154 = a29256 & a18614;
assign a30156 = a30154 & a29394;
assign a30158 = a29272 & a18590;
assign a30160 = ~a30158 & ~a30156;
assign a30162 = a30160 & a30152;
assign a30164 = a30162 & a30144;
assign a30166 = ~a30164 & a29374;
assign a30168 = ~a30148 & ~a30128;
assign a30170 = ~a30168 & ~a29270;
assign a30172 = a29254 & a18590;
assign a30174 = a30172 & a29582;
assign a30176 = ~a30174 & ~a30170;
assign a30178 = a30130 & ~a29270;
assign a30180 = a29276 & a18566;
assign a30182 = a30180 & a29592;
assign a30184 = a30154 & a29398;
assign a30186 = ~a30184 & ~a30182;
assign a30188 = a30186 & ~a30178;
assign a30190 = a30188 & a30176;
assign a30192 = a29332 & a18578;
assign a30194 = a29306 & a18604;
assign a30196 = ~a30194 & ~a30192;
assign a30198 = a29296 & a18586;
assign a30200 = a29310 & a18552;
assign a30202 = ~a30200 & ~a30198;
assign a30204 = a30202 & a30196;
assign a30206 = a30204 & a30190;
assign a30208 = ~a30206 & ~a29374;
assign a30210 = ~a30208 & ~a30166;
assign a30212 = ~a30210 & a21952;
assign a30214 = ~a30212 & a30120;
assign a30216 = a30210 & ~a21952;
assign a30218 = ~a30216 & a30214;
assign a30220 = a29328 & a18486;
assign a30222 = a29280 & a18448;
assign a30224 = ~a30222 & ~a30220;
assign a30226 = a29278 & a18454;
assign a30228 = a29294 & a18438;
assign a30230 = ~a30228 & ~a30226;
assign a30232 = ~a30230 & a29270;
assign a30234 = ~a30232 & a30224;
assign a30236 = a29290 & a18460;
assign a30238 = a29332 & a18468;
assign a30240 = ~a30238 & ~a30236;
assign a30242 = a30240 & a30234;
assign a30244 = a29322 & a18434;
assign a30246 = a29264 & a18492;
assign a30248 = a30246 & a29270;
assign a30250 = ~a30248 & ~a30244;
assign a30252 = a29256 & a18496;
assign a30254 = a30252 & a29394;
assign a30256 = a29272 & a18472;
assign a30258 = ~a30256 & ~a30254;
assign a30260 = a30258 & a30250;
assign a30262 = a30260 & a30242;
assign a30264 = ~a30262 & a29374;
assign a30266 = ~a30246 & ~a30226;
assign a30268 = ~a30266 & ~a29270;
assign a30270 = a29254 & a18472;
assign a30272 = a30270 & a29582;
assign a30274 = ~a30272 & ~a30268;
assign a30276 = a30228 & ~a29270;
assign a30278 = a29276 & a18448;
assign a30280 = a30278 & a29592;
assign a30282 = a30252 & a29398;
assign a30284 = ~a30282 & ~a30280;
assign a30286 = a30284 & ~a30276;
assign a30288 = a30286 & a30274;
assign a30290 = a29332 & a18460;
assign a30292 = a29306 & a18486;
assign a30294 = ~a30292 & ~a30290;
assign a30296 = a29296 & a18468;
assign a30298 = a29310 & a18434;
assign a30300 = ~a30298 & ~a30296;
assign a30302 = a30300 & a30294;
assign a30304 = a30302 & a30288;
assign a30306 = ~a30304 & ~a29374;
assign a30308 = ~a30306 & ~a30264;
assign a30310 = ~a30308 & a21968;
assign a30312 = ~a30310 & a30218;
assign a30314 = a30308 & ~a21968;
assign a30316 = ~a30314 & a30312;
assign a30320 = l1686 & ~l1624;
assign a30322 = a30320 & l988;
assign a30324 = ~l988 & l962;
assign a30326 = l1686 & ~l1618;
assign a30328 = l1686 & ~l1620;
assign a30330 = l1686 & ~l1622;
assign a30332 = a30330 & a30328;
assign a30334 = ~a30332 & ~a30326;
assign a30336 = a30332 & a30326;
assign a30338 = ~a30336 & ~a30334;
assign a30340 = a30338 & a30324;
assign a30342 = ~a30340 & ~a30322;
assign a30344 = ~l988 & ~l494;
assign a30346 = a30344 & ~a27452;
assign a30348 = a30346 & ~l962;
assign a30350 = a30348 & a30326;
assign a30354 = l1686 & ~l1630;
assign a30356 = l1686 & ~l1628;
assign a30358 = l1686 & ~l1626;
assign a30360 = a22640 & a15334;
assign a30362 = ~a30360 & a30320;
assign a30364 = a30360 & a30326;
assign a30368 = l1686 & ~l1636;
assign a30370 = a30368 & l988;
assign a30372 = l1686 & ~l1634;
assign a30374 = a30372 & l1622;
assign a30376 = ~a30374 & ~a30336;
assign a30378 = ~a30376 & a30324;
assign a30380 = ~a30378 & ~a30370;
assign a30382 = a30372 & a30348;
assign a30386 = l1686 & ~l1638;
assign a30388 = a30368 & ~a30360;
assign a30390 = a30372 & a30360;
assign a30394 = l1686 & ~l1642;
assign a30396 = a30394 & l988;
assign a30398 = a30330 & l1634;
assign a30400 = ~a30398 & ~a30328;
assign a30402 = ~a30400 & ~a30332;
assign a30404 = a30402 & a30324;
assign a30406 = ~a30404 & ~a30396;
assign a30408 = a30348 & a30328;
assign a30412 = a30394 & ~a30360;
assign a30414 = a30360 & a30328;
assign a30418 = l1686 & ~l1646;
assign a30420 = a30418 & l988;
assign a30422 = ~a30330 & a30324;
assign a30424 = ~a30422 & ~a30420;
assign a30426 = a30348 & a30330;
assign a30430 = a30418 & ~a30360;
assign a30432 = a30360 & a30330;
assign a30436 = a19222 & a6696;
assign a30438 = a19218 & a6708;
assign a30440 = ~a30438 & ~a30436;
assign a30442 = ~a19222 & ~a6696;
assign a30444 = ~a19224 & ~a6690;
assign a30446 = ~a30444 & ~a30442;
assign a30448 = a30446 & a30440;
assign a30450 = ~a19232 & ~a6702;
assign a30452 = a19232 & a6702;
assign a30454 = ~a30452 & ~a30450;
assign a30456 = a19224 & a6690;
assign a30458 = ~a30456 & a30454;
assign a30460 = ~a19218 & ~a6708;
assign a30462 = ~a30460 & a30458;
assign a30464 = a30462 & a30448;
assign a30466 = ~a30464 & l1660;
assign a30470 = a30468 & ~l1658;
assign a30472 = a30470 & ~a6690;
assign a30474 = ~a17946 & ~a17936;
assign a30476 = ~a6702 & ~a6690;
assign a30478 = ~a30476 & a30474;
assign a30480 = ~a30478 & l1658;
assign a30484 = a30470 & ~a6708;
assign a30486 = ~a17994 & ~a17968;
assign a30488 = ~a30486 & l1658;
assign a30492 = a30470 & ~a6702;
assign a30494 = a6702 & l1658;
assign a30498 = a30470 & ~a6696;
assign a30500 = ~a17978 & ~a17936;
assign a30502 = a30500 & ~a17930;
assign a30504 = ~a30502 & l1658;
assign a30508 = ~a6708 & a6690;
assign a30510 = a30508 & a18144;
assign a30512 = a30510 & ~a6702;
assign a30514 = ~a18104 & a6690;
assign a30516 = a30514 & a18016;
assign a30518 = ~a30516 & ~a30512;
assign a30520 = a17930 & l904;
assign a30522 = a17938 & l902;
assign a30524 = ~a30522 & ~a30520;
assign a30526 = a30524 & a30518;
assign a30528 = ~a18136 & a6690;
assign a30530 = a30528 & a18008;
assign a30532 = a6708 & l916;
assign a30534 = a30532 & ~a6702;
assign a30536 = a30534 & a17928;
assign a30538 = ~a30536 & ~a30530;
assign a30540 = a6708 & ~a6690;
assign a30542 = a30540 & l912;
assign a30544 = a30542 & ~a6696;
assign a30546 = a30544 & ~a6702;
assign a30548 = ~a30546 & a30538;
assign a30550 = a30548 & a30526;
assign a30552 = a6708 & l910;
assign a30554 = a30552 & ~a6690;
assign a30556 = a30554 & a18014;
assign a30558 = a6708 & a6690;
assign a30560 = a30558 & ~a18126;
assign a30562 = a30560 & ~a6702;
assign a30564 = a30562 & ~a6696;
assign a30566 = ~a30564 & ~a30556;
assign a30568 = a17968 & l906;
assign a30570 = ~a30568 & a30566;
assign a30572 = a30570 & a30550;
assign a30574 = ~a30572 & l1658;
assign a30576 = a30508 & l906;
assign a30578 = a30576 & a6702;
assign a30580 = a17930 & l910;
assign a30582 = ~a30580 & ~a30578;
assign a30584 = a30562 & a6696;
assign a30586 = ~a30584 & a30582;
assign a30588 = a30542 & a18006;
assign a30590 = a30540 & l902;
assign a30592 = a30590 & ~a6696;
assign a30594 = a30592 & a6702;
assign a30596 = ~a30594 & ~a30588;
assign a30598 = a30596 & a30586;
assign a30600 = ~a18104 & a17968;
assign a30602 = ~a6696 & a6690;
assign a30604 = a30602 & a30534;
assign a30606 = a30558 & l904;
assign a30608 = a30606 & a18014;
assign a30610 = ~a30608 & ~a30604;
assign a30612 = a30610 & ~a30600;
assign a30614 = a30528 & ~a6708;
assign a30616 = a18144 & a17948;
assign a30618 = ~a30616 & ~a30614;
assign a30620 = ~a30618 & ~a6702;
assign a30622 = ~a30620 & a30612;
assign a30624 = a30622 & a30598;
assign a30626 = ~a30624 & ~a30468;
assign a30628 = ~a30626 & ~a30574;
assign a30630 = a30510 & a6702;
assign a30632 = a17930 & l916;
assign a30634 = ~a30632 & ~a30630;
assign a30636 = ~a18136 & a17968;
assign a30638 = ~a30636 & a30634;
assign a30640 = a30554 & a18006;
assign a30642 = a30544 & a6702;
assign a30644 = ~a30642 & ~a30640;
assign a30646 = a30644 & a30638;
assign a30648 = a30606 & ~a6702;
assign a30650 = a30648 & ~a6696;
assign a30652 = a30560 & a18014;
assign a30654 = a30514 & ~a6702;
assign a30656 = a30654 & a17964;
assign a30658 = ~a30656 & ~a30652;
assign a30660 = a30658 & ~a30650;
assign a30662 = ~a30592 & ~a30576;
assign a30664 = ~a30662 & ~a6702;
assign a30666 = ~a30664 & a30660;
assign a30668 = a30666 & a30646;
assign a30670 = ~a30668 & a30470;
assign a30672 = ~a30670 & a30628;
assign a30674 = ~a30672 & ~l494;
assign a30676 = a30508 & a18204;
assign a30678 = a30676 & ~a6702;
assign a30680 = a18212 & a6690;
assign a30682 = a30680 & a18016;
assign a30684 = ~a30682 & ~a30678;
assign a30686 = a18256 & a17930;
assign a30688 = a18232 & a17938;
assign a30690 = ~a30688 & ~a30686;
assign a30692 = a30690 & a30684;
assign a30694 = a18218 & a6690;
assign a30696 = a30694 & a18008;
assign a30698 = a18252 & a6708;
assign a30700 = a30698 & ~a6702;
assign a30702 = a30700 & a17928;
assign a30704 = ~a30702 & ~a30696;
assign a30706 = a30540 & a18224;
assign a30708 = a30706 & ~a6696;
assign a30710 = a30708 & ~a6702;
assign a30712 = ~a30710 & a30704;
assign a30714 = a30712 & a30692;
assign a30716 = a18236 & a6708;
assign a30718 = a30716 & ~a6690;
assign a30720 = a30718 & a18014;
assign a30722 = a30558 & a18246;
assign a30724 = a30722 & ~a6702;
assign a30726 = a30724 & ~a6696;
assign a30728 = ~a30726 & ~a30720;
assign a30730 = a18200 & a17968;
assign a30732 = ~a30730 & a30728;
assign a30734 = a30732 & a30714;
assign a30736 = ~a30734 & l1658;
assign a30738 = a18200 & a17996;
assign a30740 = a18252 & a17930;
assign a30742 = ~a30740 & ~a30738;
assign a30744 = a30540 & a18232;
assign a30746 = a30744 & ~a6696;
assign a30748 = a30746 & ~a6702;
assign a30750 = ~a30748 & a30742;
assign a30752 = a30718 & a18006;
assign a30754 = a30676 & a6702;
assign a30756 = ~a30754 & ~a30752;
assign a30758 = a30558 & a18256;
assign a30760 = a30758 & ~a6702;
assign a30762 = a30760 & ~a6696;
assign a30764 = ~a30762 & a30756;
assign a30766 = a30764 & a30750;
assign a30768 = a30722 & a18014;
assign a30770 = a30680 & ~a6702;
assign a30772 = a30770 & a17964;
assign a30774 = ~a30772 & ~a30768;
assign a30776 = a30708 & a6702;
assign a30778 = ~a30776 & a30774;
assign a30780 = a18218 & a17968;
assign a30782 = ~a30780 & a30778;
assign a30784 = a30782 & a30766;
assign a30786 = ~a30784 & a30470;
assign a30788 = ~a30786 & ~a30736;
assign a30790 = a18200 & a17938;
assign a30792 = a18236 & a17930;
assign a30794 = ~a30792 & ~a30790;
assign a30796 = a30724 & a6696;
assign a30798 = ~a30796 & a30794;
assign a30800 = a30706 & a18006;
assign a30802 = a30746 & a6702;
assign a30804 = ~a30802 & ~a30800;
assign a30806 = a30804 & a30798;
assign a30808 = a18212 & a17968;
assign a30810 = a30700 & a30602;
assign a30812 = a30758 & a18014;
assign a30814 = ~a30812 & ~a30810;
assign a30816 = a30814 & ~a30808;
assign a30818 = a30694 & ~a6708;
assign a30820 = a18204 & a17948;
assign a30822 = ~a30820 & ~a30818;
assign a30824 = ~a30822 & ~a6702;
assign a30826 = ~a30824 & a30816;
assign a30828 = a30826 & a30806;
assign a30830 = ~a30828 & ~a30468;
assign a30832 = ~a30830 & a30788;
assign a30834 = ~a30832 & a16304;
assign a30836 = a30832 & ~a16304;
assign a30838 = ~a30836 & ~a30834;
assign a30840 = a30508 & a18320;
assign a30842 = a30840 & ~a6702;
assign a30844 = a18328 & a6690;
assign a30846 = a30844 & a18016;
assign a30848 = ~a30846 & ~a30842;
assign a30850 = a18376 & a17930;
assign a30852 = a18348 & a17938;
assign a30854 = ~a30852 & ~a30850;
assign a30856 = a30854 & a30848;
assign a30858 = a18334 & a6690;
assign a30860 = a30858 & a18008;
assign a30862 = a18372 & a6708;
assign a30864 = a30862 & ~a6702;
assign a30866 = a30864 & a17928;
assign a30868 = ~a30866 & ~a30860;
assign a30870 = a30540 & a18340;
assign a30872 = a30870 & ~a6696;
assign a30874 = a30872 & ~a6702;
assign a30876 = ~a30874 & a30868;
assign a30878 = a30876 & a30856;
assign a30880 = a18352 & a6708;
assign a30882 = a30880 & ~a6690;
assign a30884 = a30882 & a18014;
assign a30886 = a30558 & a18366;
assign a30888 = a30886 & ~a6702;
assign a30890 = a30888 & ~a6696;
assign a30892 = ~a30890 & ~a30884;
assign a30894 = a18316 & a17968;
assign a30896 = ~a30894 & a30892;
assign a30898 = a30896 & a30878;
assign a30900 = ~a30898 & l1658;
assign a30902 = a30840 & a6702;
assign a30904 = a18372 & a17930;
assign a30906 = ~a30904 & ~a30902;
assign a30908 = a18334 & a17968;
assign a30910 = ~a30908 & a30906;
assign a30912 = a30882 & a18006;
assign a30914 = a30872 & a6702;
assign a30916 = ~a30914 & ~a30912;
assign a30918 = a30916 & a30910;
assign a30920 = a30558 & a18376;
assign a30922 = a30920 & ~a6702;
assign a30924 = a30922 & ~a6696;
assign a30926 = a30886 & a18014;
assign a30928 = a30844 & ~a6702;
assign a30930 = a30928 & a17964;
assign a30932 = ~a30930 & ~a30926;
assign a30934 = a30932 & ~a30924;
assign a30936 = a30508 & a18316;
assign a30938 = a30540 & a18348;
assign a30940 = a30938 & ~a6696;
assign a30942 = ~a30940 & ~a30936;
assign a30944 = ~a30942 & ~a6702;
assign a30946 = ~a30944 & a30934;
assign a30948 = a30946 & a30918;
assign a30950 = ~a30948 & a30470;
assign a30952 = ~a30950 & ~a30900;
assign a30954 = a30936 & a6702;
assign a30956 = a18352 & a17930;
assign a30958 = ~a30956 & ~a30954;
assign a30960 = a30888 & a6696;
assign a30962 = ~a30960 & a30958;
assign a30964 = a30870 & a18006;
assign a30966 = a30940 & a6702;
assign a30968 = ~a30966 & ~a30964;
assign a30970 = a30968 & a30962;
assign a30972 = a18328 & a17968;
assign a30974 = a30864 & a30602;
assign a30976 = a30920 & a18014;
assign a30978 = ~a30976 & ~a30974;
assign a30980 = a30978 & ~a30972;
assign a30982 = a30858 & ~a6708;
assign a30984 = a18320 & a17948;
assign a30986 = ~a30984 & ~a30982;
assign a30988 = ~a30986 & ~a6702;
assign a30990 = ~a30988 & a30980;
assign a30992 = a30990 & a30970;
assign a30994 = ~a30992 & ~a30468;
assign a30996 = ~a30994 & a30952;
assign a30998 = ~a30996 & a16298;
assign a31000 = ~a30998 & ~a30838;
assign a31002 = a30508 & a18438;
assign a31004 = a31002 & ~a6702;
assign a31006 = a18448 & a6690;
assign a31008 = a31006 & a18016;
assign a31010 = ~a31008 & ~a31004;
assign a31012 = a18496 & a17930;
assign a31014 = a18468 & a17938;
assign a31016 = ~a31014 & ~a31012;
assign a31018 = a31016 & a31010;
assign a31020 = a18454 & a6690;
assign a31022 = a31020 & a18008;
assign a31024 = a18492 & a6708;
assign a31026 = a31024 & ~a6702;
assign a31028 = a31026 & a17928;
assign a31030 = ~a31028 & ~a31022;
assign a31032 = a30540 & a18460;
assign a31034 = a31032 & ~a6696;
assign a31036 = a31034 & ~a6702;
assign a31038 = ~a31036 & a31030;
assign a31040 = a31038 & a31018;
assign a31042 = a18472 & a6708;
assign a31044 = a31042 & ~a6690;
assign a31046 = a31044 & a18014;
assign a31048 = a30558 & a18486;
assign a31050 = a31048 & ~a6702;
assign a31052 = a31050 & ~a6696;
assign a31054 = ~a31052 & ~a31046;
assign a31056 = a18434 & a17968;
assign a31058 = ~a31056 & a31054;
assign a31060 = a31058 & a31040;
assign a31062 = ~a31060 & l1658;
assign a31064 = a18434 & a17996;
assign a31066 = a18492 & a17930;
assign a31068 = ~a31066 & ~a31064;
assign a31070 = a30540 & a18468;
assign a31072 = a31070 & ~a6696;
assign a31074 = a31072 & ~a6702;
assign a31076 = ~a31074 & a31068;
assign a31078 = a31044 & a18006;
assign a31080 = a31002 & a6702;
assign a31082 = ~a31080 & ~a31078;
assign a31084 = a30558 & a18496;
assign a31086 = a31084 & ~a6702;
assign a31088 = a31086 & ~a6696;
assign a31090 = ~a31088 & a31082;
assign a31092 = a31090 & a31076;
assign a31094 = a31048 & a18014;
assign a31096 = a31006 & ~a6702;
assign a31098 = a31096 & a17964;
assign a31100 = ~a31098 & ~a31094;
assign a31102 = a31034 & a6702;
assign a31104 = ~a31102 & a31100;
assign a31106 = a18454 & a17968;
assign a31108 = ~a31106 & a31104;
assign a31110 = a31108 & a31092;
assign a31112 = ~a31110 & a30470;
assign a31114 = ~a31112 & ~a31062;
assign a31116 = a18434 & a17938;
assign a31118 = a18472 & a17930;
assign a31120 = ~a31118 & ~a31116;
assign a31122 = a31050 & a6696;
assign a31124 = ~a31122 & a31120;
assign a31126 = a31032 & a18006;
assign a31128 = a31072 & a6702;
assign a31130 = ~a31128 & ~a31126;
assign a31132 = a31130 & a31124;
assign a31134 = a18448 & a17968;
assign a31136 = a31026 & a30602;
assign a31138 = a31084 & a18014;
assign a31140 = ~a31138 & ~a31136;
assign a31142 = a31140 & ~a31134;
assign a31144 = a31020 & ~a6708;
assign a31146 = a18438 & a17948;
assign a31148 = ~a31146 & ~a31144;
assign a31150 = ~a31148 & ~a6702;
assign a31152 = ~a31150 & a31142;
assign a31154 = a31152 & a31132;
assign a31156 = ~a31154 & ~a30468;
assign a31158 = ~a31156 & a31114;
assign a31160 = a31158 & ~a16310;
assign a31162 = a30508 & a18556;
assign a31164 = a31162 & ~a6702;
assign a31166 = a18566 & a6690;
assign a31168 = a31166 & a18016;
assign a31170 = ~a31168 & ~a31164;
assign a31172 = a18614 & a17930;
assign a31174 = a18586 & a17938;
assign a31176 = ~a31174 & ~a31172;
assign a31178 = a31176 & a31170;
assign a31180 = a18572 & a6690;
assign a31182 = a31180 & a18008;
assign a31184 = a18610 & a6708;
assign a31186 = a31184 & ~a6702;
assign a31188 = a31186 & a17928;
assign a31190 = ~a31188 & ~a31182;
assign a31192 = a30540 & a18578;
assign a31194 = a31192 & ~a6696;
assign a31196 = a31194 & ~a6702;
assign a31198 = ~a31196 & a31190;
assign a31200 = a31198 & a31178;
assign a31202 = a18590 & a6708;
assign a31204 = a31202 & ~a6690;
assign a31206 = a31204 & a18014;
assign a31208 = a30558 & a18604;
assign a31210 = a31208 & ~a6702;
assign a31212 = a31210 & ~a6696;
assign a31214 = ~a31212 & ~a31206;
assign a31216 = a18552 & a17968;
assign a31218 = ~a31216 & a31214;
assign a31220 = a31218 & a31200;
assign a31222 = ~a31220 & l1658;
assign a31224 = a18552 & a17996;
assign a31226 = a18610 & a17930;
assign a31228 = ~a31226 & ~a31224;
assign a31230 = a30540 & a18586;
assign a31232 = a31230 & ~a6696;
assign a31234 = a31232 & ~a6702;
assign a31236 = ~a31234 & a31228;
assign a31238 = a31204 & a18006;
assign a31240 = a31162 & a6702;
assign a31242 = ~a31240 & ~a31238;
assign a31244 = a30558 & a18614;
assign a31246 = a31244 & ~a6702;
assign a31248 = a31246 & ~a6696;
assign a31250 = ~a31248 & a31242;
assign a31252 = a31250 & a31236;
assign a31254 = a31208 & a18014;
assign a31256 = a31166 & ~a6702;
assign a31258 = a31256 & a17964;
assign a31260 = ~a31258 & ~a31254;
assign a31262 = a31194 & a6702;
assign a31264 = ~a31262 & a31260;
assign a31266 = a18572 & a17968;
assign a31268 = ~a31266 & a31264;
assign a31270 = a31268 & a31252;
assign a31272 = ~a31270 & a30470;
assign a31274 = ~a31272 & ~a31222;
assign a31276 = a18552 & a17938;
assign a31278 = a18590 & a17930;
assign a31280 = ~a31278 & ~a31276;
assign a31282 = a31210 & a6696;
assign a31284 = ~a31282 & a31280;
assign a31286 = a31192 & a18006;
assign a31288 = a31232 & a6702;
assign a31290 = ~a31288 & ~a31286;
assign a31292 = a31290 & a31284;
assign a31294 = a18566 & a17968;
assign a31296 = a31186 & a30602;
assign a31298 = a31244 & a18014;
assign a31300 = ~a31298 & ~a31296;
assign a31302 = a31300 & ~a31294;
assign a31304 = a31180 & ~a6708;
assign a31306 = a18556 & a17948;
assign a31308 = ~a31306 & ~a31304;
assign a31310 = ~a31308 & ~a6702;
assign a31312 = ~a31310 & a31302;
assign a31314 = a31312 & a31292;
assign a31316 = ~a31314 & ~a30468;
assign a31318 = ~a31316 & a31274;
assign a31320 = a31318 & ~a16268;
assign a31322 = ~a31320 & ~a31160;
assign a31324 = ~a31318 & a16268;
assign a31326 = ~a31324 & ~a31322;
assign a31328 = a30508 & a18680;
assign a31330 = a31328 & ~a6702;
assign a31332 = a18690 & a6690;
assign a31334 = a31332 & a18016;
assign a31336 = ~a31334 & ~a31330;
assign a31338 = a18738 & a17930;
assign a31340 = a18710 & a17938;
assign a31342 = ~a31340 & ~a31338;
assign a31344 = a31342 & a31336;
assign a31346 = a18696 & a6690;
assign a31348 = a31346 & a18008;
assign a31350 = a18734 & a6708;
assign a31352 = a31350 & ~a6702;
assign a31354 = a31352 & a17928;
assign a31356 = ~a31354 & ~a31348;
assign a31358 = a30540 & a18702;
assign a31360 = a31358 & ~a6696;
assign a31362 = a31360 & ~a6702;
assign a31364 = ~a31362 & a31356;
assign a31366 = a31364 & a31344;
assign a31368 = a18714 & a6708;
assign a31370 = a31368 & ~a6690;
assign a31372 = a31370 & a18014;
assign a31374 = a30558 & a18728;
assign a31376 = a31374 & ~a6702;
assign a31378 = a31376 & ~a6696;
assign a31380 = ~a31378 & ~a31372;
assign a31382 = a18676 & a17968;
assign a31384 = ~a31382 & a31380;
assign a31386 = a31384 & a31366;
assign a31388 = ~a31386 & l1658;
assign a31390 = a31328 & a6702;
assign a31392 = a18734 & a17930;
assign a31394 = ~a31392 & ~a31390;
assign a31396 = a18696 & a17968;
assign a31398 = ~a31396 & a31394;
assign a31400 = a31370 & a18006;
assign a31402 = a31360 & a6702;
assign a31404 = ~a31402 & ~a31400;
assign a31406 = a31404 & a31398;
assign a31408 = a30558 & a18738;
assign a31410 = a31408 & ~a6702;
assign a31412 = a31410 & ~a6696;
assign a31414 = a31374 & a18014;
assign a31416 = a31332 & ~a6702;
assign a31418 = a31416 & a17964;
assign a31420 = ~a31418 & ~a31414;
assign a31422 = a31420 & ~a31412;
assign a31424 = a30508 & a18676;
assign a31426 = a30540 & a18710;
assign a31428 = a31426 & ~a6696;
assign a31430 = ~a31428 & ~a31424;
assign a31432 = ~a31430 & ~a6702;
assign a31434 = ~a31432 & a31422;
assign a31436 = a31434 & a31406;
assign a31438 = ~a31436 & a30470;
assign a31440 = ~a31438 & ~a31388;
assign a31442 = a31424 & a6702;
assign a31444 = a18714 & a17930;
assign a31446 = ~a31444 & ~a31442;
assign a31448 = a31376 & a6696;
assign a31450 = ~a31448 & a31446;
assign a31452 = a31358 & a18006;
assign a31454 = a31428 & a6702;
assign a31456 = ~a31454 & ~a31452;
assign a31458 = a31456 & a31450;
assign a31460 = a18690 & a17968;
assign a31462 = a31352 & a30602;
assign a31464 = a31408 & a18014;
assign a31466 = ~a31464 & ~a31462;
assign a31468 = a31466 & ~a31460;
assign a31470 = a31346 & ~a6708;
assign a31472 = a18680 & a17948;
assign a31474 = ~a31472 & ~a31470;
assign a31476 = ~a31474 & ~a6702;
assign a31478 = ~a31476 & a31468;
assign a31480 = a31478 & a31458;
assign a31482 = ~a31480 & ~a30468;
assign a31484 = ~a31482 & a31440;
assign a31486 = a31484 & ~a16274;
assign a31488 = ~a31486 & ~a31326;
assign a31490 = ~a31484 & a16274;
assign a31492 = ~a31490 & ~a31488;
assign a31494 = a30508 & a18804;
assign a31496 = a31494 & ~a6702;
assign a31498 = a18814 & a6690;
assign a31500 = a31498 & a18016;
assign a31502 = ~a31500 & ~a31496;
assign a31504 = a18862 & a17930;
assign a31506 = a18834 & a17938;
assign a31508 = ~a31506 & ~a31504;
assign a31510 = a31508 & a31502;
assign a31512 = a18820 & a6690;
assign a31514 = a31512 & a18008;
assign a31516 = a18858 & a6708;
assign a31518 = a31516 & ~a6702;
assign a31520 = a31518 & a17928;
assign a31522 = ~a31520 & ~a31514;
assign a31524 = a30540 & a18826;
assign a31526 = a31524 & ~a6696;
assign a31528 = a31526 & ~a6702;
assign a31530 = ~a31528 & a31522;
assign a31532 = a31530 & a31510;
assign a31534 = a18838 & a6708;
assign a31536 = a31534 & ~a6690;
assign a31538 = a31536 & a18014;
assign a31540 = a30558 & a18852;
assign a31542 = a31540 & ~a6702;
assign a31544 = a31542 & ~a6696;
assign a31546 = ~a31544 & ~a31538;
assign a31548 = a18800 & a17968;
assign a31550 = ~a31548 & a31546;
assign a31552 = a31550 & a31532;
assign a31554 = ~a31552 & l1658;
assign a31556 = a31494 & a6702;
assign a31558 = a18858 & a17930;
assign a31560 = ~a31558 & ~a31556;
assign a31562 = a18820 & a17968;
assign a31564 = ~a31562 & a31560;
assign a31566 = a31536 & a18006;
assign a31568 = a31526 & a6702;
assign a31570 = ~a31568 & ~a31566;
assign a31572 = a31570 & a31564;
assign a31574 = a30558 & a18862;
assign a31576 = a31574 & ~a6702;
assign a31578 = a31576 & ~a6696;
assign a31580 = a31540 & a18014;
assign a31582 = a31498 & ~a6702;
assign a31584 = a31582 & a17964;
assign a31586 = ~a31584 & ~a31580;
assign a31588 = a31586 & ~a31578;
assign a31590 = a30508 & a18800;
assign a31592 = a30540 & a18834;
assign a31594 = a31592 & ~a6696;
assign a31596 = ~a31594 & ~a31590;
assign a31598 = ~a31596 & ~a6702;
assign a31600 = ~a31598 & a31588;
assign a31602 = a31600 & a31572;
assign a31604 = ~a31602 & a30470;
assign a31606 = ~a31604 & ~a31554;
assign a31608 = a31590 & a6702;
assign a31610 = a18838 & a17930;
assign a31612 = ~a31610 & ~a31608;
assign a31614 = a31542 & a6696;
assign a31616 = ~a31614 & a31612;
assign a31618 = a31524 & a18006;
assign a31620 = a31594 & a6702;
assign a31622 = ~a31620 & ~a31618;
assign a31624 = a31622 & a31616;
assign a31626 = a18814 & a17968;
assign a31628 = a31518 & a30602;
assign a31630 = a31574 & a18014;
assign a31632 = ~a31630 & ~a31628;
assign a31634 = a31632 & ~a31626;
assign a31636 = a31512 & ~a6708;
assign a31638 = a18804 & a17948;
assign a31640 = ~a31638 & ~a31636;
assign a31642 = ~a31640 & ~a6702;
assign a31644 = ~a31642 & a31634;
assign a31646 = a31644 & a31624;
assign a31648 = ~a31646 & ~a30468;
assign a31650 = ~a31648 & a31606;
assign a31652 = a31650 & ~a16280;
assign a31654 = ~a31652 & ~a31492;
assign a31656 = ~a31650 & a16280;
assign a31658 = ~a31656 & ~a31654;
assign a31660 = a30508 & a18928;
assign a31662 = a31660 & ~a6702;
assign a31664 = a18938 & a6690;
assign a31666 = a31664 & a18016;
assign a31668 = ~a31666 & ~a31662;
assign a31670 = a18986 & a17930;
assign a31672 = a18958 & a17938;
assign a31674 = ~a31672 & ~a31670;
assign a31676 = a31674 & a31668;
assign a31678 = a18944 & a6690;
assign a31680 = a31678 & a18008;
assign a31682 = a18982 & a6708;
assign a31684 = a31682 & ~a6702;
assign a31686 = a31684 & a17928;
assign a31688 = ~a31686 & ~a31680;
assign a31690 = a30540 & a18950;
assign a31692 = a31690 & ~a6696;
assign a31694 = a31692 & ~a6702;
assign a31696 = ~a31694 & a31688;
assign a31698 = a31696 & a31676;
assign a31700 = a18962 & a6708;
assign a31702 = a31700 & ~a6690;
assign a31704 = a31702 & a18014;
assign a31706 = a30558 & a18976;
assign a31708 = a31706 & ~a6702;
assign a31710 = a31708 & ~a6696;
assign a31712 = ~a31710 & ~a31704;
assign a31714 = a18924 & a17968;
assign a31716 = ~a31714 & a31712;
assign a31718 = a31716 & a31698;
assign a31720 = ~a31718 & l1658;
assign a31722 = a31660 & a6702;
assign a31724 = a18982 & a17930;
assign a31726 = ~a31724 & ~a31722;
assign a31728 = a18944 & a17968;
assign a31730 = ~a31728 & a31726;
assign a31732 = a31702 & a18006;
assign a31734 = a31692 & a6702;
assign a31736 = ~a31734 & ~a31732;
assign a31738 = a31736 & a31730;
assign a31740 = a30558 & a18986;
assign a31742 = a31740 & ~a6702;
assign a31744 = a31742 & ~a6696;
assign a31746 = a31706 & a18014;
assign a31748 = a31664 & ~a6702;
assign a31750 = a31748 & a17964;
assign a31752 = ~a31750 & ~a31746;
assign a31754 = a31752 & ~a31744;
assign a31756 = a30508 & a18924;
assign a31758 = a30540 & a18958;
assign a31760 = a31758 & ~a6696;
assign a31762 = ~a31760 & ~a31756;
assign a31764 = ~a31762 & ~a6702;
assign a31766 = ~a31764 & a31754;
assign a31768 = a31766 & a31738;
assign a31770 = ~a31768 & a30470;
assign a31772 = ~a31770 & ~a31720;
assign a31774 = a31756 & a6702;
assign a31776 = a18962 & a17930;
assign a31778 = ~a31776 & ~a31774;
assign a31780 = a31708 & a6696;
assign a31782 = ~a31780 & a31778;
assign a31784 = a31690 & a18006;
assign a31786 = a31760 & a6702;
assign a31788 = ~a31786 & ~a31784;
assign a31790 = a31788 & a31782;
assign a31792 = a18938 & a17968;
assign a31794 = a31684 & a30602;
assign a31796 = a31740 & a18014;
assign a31798 = ~a31796 & ~a31794;
assign a31800 = a31798 & ~a31792;
assign a31802 = a31678 & ~a6708;
assign a31804 = a18928 & a17948;
assign a31806 = ~a31804 & ~a31802;
assign a31808 = ~a31806 & ~a6702;
assign a31810 = ~a31808 & a31800;
assign a31812 = a31810 & a31790;
assign a31814 = ~a31812 & ~a30468;
assign a31816 = ~a31814 & a31772;
assign a31818 = a31816 & ~a16286;
assign a31820 = ~a31818 & ~a31658;
assign a31822 = ~a31816 & a16286;
assign a31824 = ~a31822 & ~a31820;
assign a31826 = a30508 & a19052;
assign a31828 = a31826 & ~a6702;
assign a31830 = a19062 & a6690;
assign a31832 = a31830 & a18016;
assign a31834 = ~a31832 & ~a31828;
assign a31836 = a19110 & a17930;
assign a31838 = a19082 & a17938;
assign a31840 = ~a31838 & ~a31836;
assign a31842 = a31840 & a31834;
assign a31844 = a19068 & a6690;
assign a31846 = a31844 & a18008;
assign a31848 = a19106 & a6708;
assign a31850 = a31848 & ~a6702;
assign a31852 = a31850 & a17928;
assign a31854 = ~a31852 & ~a31846;
assign a31856 = a30540 & a19074;
assign a31858 = a31856 & ~a6696;
assign a31860 = a31858 & ~a6702;
assign a31862 = ~a31860 & a31854;
assign a31864 = a31862 & a31842;
assign a31866 = a19086 & a6708;
assign a31868 = a31866 & ~a6690;
assign a31870 = a31868 & a18014;
assign a31872 = a30558 & a19100;
assign a31874 = a31872 & ~a6702;
assign a31876 = a31874 & ~a6696;
assign a31878 = ~a31876 & ~a31870;
assign a31880 = a19048 & a17968;
assign a31882 = ~a31880 & a31878;
assign a31884 = a31882 & a31864;
assign a31886 = ~a31884 & l1658;
assign a31888 = a31826 & a6702;
assign a31890 = a19106 & a17930;
assign a31892 = ~a31890 & ~a31888;
assign a31894 = a19068 & a17968;
assign a31896 = ~a31894 & a31892;
assign a31898 = a31868 & a18006;
assign a31900 = a31858 & a6702;
assign a31902 = ~a31900 & ~a31898;
assign a31904 = a31902 & a31896;
assign a31906 = a30558 & a19110;
assign a31908 = a31906 & ~a6702;
assign a31910 = a31908 & ~a6696;
assign a31912 = a31872 & a18014;
assign a31914 = a31830 & ~a6702;
assign a31916 = a31914 & a17964;
assign a31918 = ~a31916 & ~a31912;
assign a31920 = a31918 & ~a31910;
assign a31922 = a30508 & a19048;
assign a31924 = a30540 & a19082;
assign a31926 = a31924 & ~a6696;
assign a31928 = ~a31926 & ~a31922;
assign a31930 = ~a31928 & ~a6702;
assign a31932 = ~a31930 & a31920;
assign a31934 = a31932 & a31904;
assign a31936 = ~a31934 & a30470;
assign a31938 = ~a31936 & ~a31886;
assign a31940 = a31922 & a6702;
assign a31942 = a19086 & a17930;
assign a31944 = ~a31942 & ~a31940;
assign a31946 = a31874 & a6696;
assign a31948 = ~a31946 & a31944;
assign a31950 = a31856 & a18006;
assign a31952 = a31926 & a6702;
assign a31954 = ~a31952 & ~a31950;
assign a31956 = a31954 & a31948;
assign a31958 = a19062 & a17968;
assign a31960 = a31850 & a30602;
assign a31962 = a31906 & a18014;
assign a31964 = ~a31962 & ~a31960;
assign a31966 = a31964 & ~a31958;
assign a31968 = a31844 & ~a6708;
assign a31970 = a19052 & a17948;
assign a31972 = ~a31970 & ~a31968;
assign a31974 = ~a31972 & ~a6702;
assign a31976 = ~a31974 & a31966;
assign a31978 = a31976 & a31956;
assign a31980 = ~a31978 & ~a30468;
assign a31982 = ~a31980 & a31938;
assign a31984 = a31982 & ~a16292;
assign a31986 = ~a31984 & ~a31824;
assign a31988 = ~a31982 & a16292;
assign a31990 = ~a31988 & ~a31986;
assign a31992 = a30996 & ~a16298;
assign a31994 = ~a31992 & ~a31990;
assign a31996 = ~a31994 & a31000;
assign a31998 = ~a31992 & a30838;
assign a32000 = ~a31158 & a16310;
assign a32002 = ~a32000 & ~a31324;
assign a32004 = ~a32002 & ~a31320;
assign a32006 = ~a32004 & ~a31490;
assign a32008 = ~a32006 & ~a31486;
assign a32010 = ~a32008 & ~a31656;
assign a32012 = ~a32010 & ~a31652;
assign a32014 = ~a32012 & ~a31822;
assign a32016 = ~a32014 & ~a31818;
assign a32018 = ~a32016 & ~a31988;
assign a32020 = ~a32018 & ~a31984;
assign a32022 = ~a32020 & ~a30998;
assign a32024 = ~a32022 & a31998;
assign a32026 = ~a32024 & ~a31996;
assign a32030 = a30602 & a6702;
assign a32032 = a32030 & a30532;
assign a32034 = a30590 & a18006;
assign a32036 = ~a32034 & ~a32032;
assign a32038 = ~a18126 & a17968;
assign a32040 = ~a32038 & a32036;
assign a32042 = a30552 & a17980;
assign a32044 = a17930 & l912;
assign a32046 = ~a32044 & ~a32042;
assign a32048 = a30648 & a6696;
assign a32050 = ~a32048 & a32046;
assign a32052 = a32050 & a32040;
assign a32054 = ~a30618 & a6702;
assign a32056 = a30654 & ~a6708;
assign a32058 = ~a32056 & ~a32054;
assign a32060 = a17950 & l906;
assign a32062 = ~a32060 & a32058;
assign a32064 = a32062 & a32052;
assign a32066 = ~a32064 & ~a30468;
assign a32068 = ~a30624 & a30470;
assign a32070 = ~a32068 & ~a32066;
assign a32072 = ~a30668 & l1658;
assign a32074 = ~a32072 & a32070;
assign a32076 = ~a30784 & l1658;
assign a32078 = a30770 & ~a6708;
assign a32080 = a18224 & a17930;
assign a32082 = ~a32080 & ~a32078;
assign a32084 = a18200 & a17950;
assign a32086 = ~a32084 & a32082;
assign a32088 = a30744 & a18006;
assign a32090 = a30818 & a6702;
assign a32092 = ~a32090 & ~a32088;
assign a32094 = a18246 & a17968;
assign a32096 = ~a32094 & a32092;
assign a32098 = a32096 & a32086;
assign a32100 = a30716 & a17980;
assign a32102 = a32030 & a30698;
assign a32104 = ~a32102 & ~a32100;
assign a32106 = a30820 & a6702;
assign a32108 = ~a32106 & a32104;
assign a32110 = a30760 & a6696;
assign a32112 = ~a32110 & a32108;
assign a32114 = a32112 & a32098;
assign a32116 = ~a32114 & ~a30468;
assign a32118 = ~a32116 & ~a32076;
assign a32120 = ~a30828 & a30470;
assign a32122 = ~a32120 & a32118;
assign a32124 = ~a32122 & a16304;
assign a32126 = a32122 & ~a16304;
assign a32128 = ~a32126 & ~a32124;
assign a32130 = ~a30948 & l1658;
assign a32132 = a30928 & ~a6708;
assign a32134 = a18340 & a17930;
assign a32136 = ~a32134 & ~a32132;
assign a32138 = a18316 & a17950;
assign a32140 = ~a32138 & a32136;
assign a32142 = a30938 & a18006;
assign a32144 = a30982 & a6702;
assign a32146 = ~a32144 & ~a32142;
assign a32148 = a18366 & a17968;
assign a32150 = ~a32148 & a32146;
assign a32152 = a32150 & a32140;
assign a32154 = a30880 & a17980;
assign a32156 = a32030 & a30862;
assign a32158 = ~a32156 & ~a32154;
assign a32160 = a30984 & a6702;
assign a32162 = ~a32160 & a32158;
assign a32164 = a30922 & a6696;
assign a32166 = ~a32164 & a32162;
assign a32168 = a32166 & a32152;
assign a32170 = ~a32168 & ~a30468;
assign a32172 = ~a32170 & ~a32130;
assign a32174 = ~a30992 & a30470;
assign a32176 = ~a32174 & a32172;
assign a32178 = a32176 & ~a16298;
assign a32180 = ~a32178 & a32128;
assign a32182 = ~a31110 & l1658;
assign a32184 = a31096 & ~a6708;
assign a32186 = a18460 & a17930;
assign a32188 = ~a32186 & ~a32184;
assign a32190 = a18434 & a17950;
assign a32192 = ~a32190 & a32188;
assign a32194 = a31070 & a18006;
assign a32196 = a31144 & a6702;
assign a32198 = ~a32196 & ~a32194;
assign a32200 = a18486 & a17968;
assign a32202 = ~a32200 & a32198;
assign a32204 = a32202 & a32192;
assign a32206 = a31042 & a17980;
assign a32208 = a32030 & a31024;
assign a32210 = ~a32208 & ~a32206;
assign a32212 = a31146 & a6702;
assign a32214 = ~a32212 & a32210;
assign a32216 = a31086 & a6696;
assign a32218 = ~a32216 & a32214;
assign a32220 = a32218 & a32204;
assign a32222 = ~a32220 & ~a30468;
assign a32224 = ~a32222 & ~a32182;
assign a32226 = ~a31154 & a30470;
assign a32228 = ~a32226 & a32224;
assign a32230 = ~a32228 & a16310;
assign a32232 = ~a31270 & l1658;
assign a32234 = a31256 & ~a6708;
assign a32236 = a18578 & a17930;
assign a32238 = ~a32236 & ~a32234;
assign a32240 = a18552 & a17950;
assign a32242 = ~a32240 & a32238;
assign a32244 = a31230 & a18006;
assign a32246 = a31304 & a6702;
assign a32248 = ~a32246 & ~a32244;
assign a32250 = a18604 & a17968;
assign a32252 = ~a32250 & a32248;
assign a32254 = a32252 & a32242;
assign a32256 = a31202 & a17980;
assign a32258 = a32030 & a31184;
assign a32260 = ~a32258 & ~a32256;
assign a32262 = a31306 & a6702;
assign a32264 = ~a32262 & a32260;
assign a32266 = a31246 & a6696;
assign a32268 = ~a32266 & a32264;
assign a32270 = a32268 & a32254;
assign a32272 = ~a32270 & ~a30468;
assign a32274 = ~a32272 & ~a32232;
assign a32276 = ~a31314 & a30470;
assign a32278 = ~a32276 & a32274;
assign a32280 = ~a32278 & a16268;
assign a32282 = ~a32280 & ~a32230;
assign a32284 = a32278 & ~a16268;
assign a32286 = ~a32284 & ~a32282;
assign a32288 = ~a31436 & l1658;
assign a32290 = a31416 & ~a6708;
assign a32292 = a18702 & a17930;
assign a32294 = ~a32292 & ~a32290;
assign a32296 = a18676 & a17950;
assign a32298 = ~a32296 & a32294;
assign a32300 = a31426 & a18006;
assign a32302 = a31470 & a6702;
assign a32304 = ~a32302 & ~a32300;
assign a32306 = a18728 & a17968;
assign a32308 = ~a32306 & a32304;
assign a32310 = a32308 & a32298;
assign a32312 = a31368 & a17980;
assign a32314 = a32030 & a31350;
assign a32316 = ~a32314 & ~a32312;
assign a32318 = a31472 & a6702;
assign a32320 = ~a32318 & a32316;
assign a32322 = a31410 & a6696;
assign a32324 = ~a32322 & a32320;
assign a32326 = a32324 & a32310;
assign a32328 = ~a32326 & ~a30468;
assign a32330 = ~a32328 & ~a32288;
assign a32332 = ~a31480 & a30470;
assign a32334 = ~a32332 & a32330;
assign a32336 = ~a32334 & a16274;
assign a32338 = ~a32336 & ~a32286;
assign a32340 = a32334 & ~a16274;
assign a32342 = ~a32340 & ~a32338;
assign a32344 = ~a31602 & l1658;
assign a32346 = a31582 & ~a6708;
assign a32348 = a18826 & a17930;
assign a32350 = ~a32348 & ~a32346;
assign a32352 = a18800 & a17950;
assign a32354 = ~a32352 & a32350;
assign a32356 = a31592 & a18006;
assign a32358 = a31636 & a6702;
assign a32360 = ~a32358 & ~a32356;
assign a32362 = a18852 & a17968;
assign a32364 = ~a32362 & a32360;
assign a32366 = a32364 & a32354;
assign a32368 = a31534 & a17980;
assign a32370 = a32030 & a31516;
assign a32372 = ~a32370 & ~a32368;
assign a32374 = a31638 & a6702;
assign a32376 = ~a32374 & a32372;
assign a32378 = a31576 & a6696;
assign a32380 = ~a32378 & a32376;
assign a32382 = a32380 & a32366;
assign a32384 = ~a32382 & ~a30468;
assign a32386 = ~a32384 & ~a32344;
assign a32388 = ~a31646 & a30470;
assign a32390 = ~a32388 & a32386;
assign a32392 = ~a32390 & a16280;
assign a32394 = ~a32392 & ~a32342;
assign a32396 = a32390 & ~a16280;
assign a32398 = ~a32396 & ~a32394;
assign a32400 = ~a31768 & l1658;
assign a32402 = a31748 & ~a6708;
assign a32404 = a18950 & a17930;
assign a32406 = ~a32404 & ~a32402;
assign a32408 = a18924 & a17950;
assign a32410 = ~a32408 & a32406;
assign a32412 = a31758 & a18006;
assign a32414 = a31802 & a6702;
assign a32416 = ~a32414 & ~a32412;
assign a32418 = a18976 & a17968;
assign a32420 = ~a32418 & a32416;
assign a32422 = a32420 & a32410;
assign a32424 = a31700 & a17980;
assign a32426 = a32030 & a31682;
assign a32428 = ~a32426 & ~a32424;
assign a32430 = a31804 & a6702;
assign a32432 = ~a32430 & a32428;
assign a32434 = a31742 & a6696;
assign a32436 = ~a32434 & a32432;
assign a32438 = a32436 & a32422;
assign a32440 = ~a32438 & ~a30468;
assign a32442 = ~a32440 & ~a32400;
assign a32444 = ~a31812 & a30470;
assign a32446 = ~a32444 & a32442;
assign a32448 = ~a32446 & a16286;
assign a32450 = ~a32448 & ~a32398;
assign a32452 = a32446 & ~a16286;
assign a32454 = ~a32452 & ~a32450;
assign a32456 = ~a31934 & l1658;
assign a32458 = a31914 & ~a6708;
assign a32460 = a19074 & a17930;
assign a32462 = ~a32460 & ~a32458;
assign a32464 = a19048 & a17950;
assign a32466 = ~a32464 & a32462;
assign a32468 = a31924 & a18006;
assign a32470 = a31968 & a6702;
assign a32472 = ~a32470 & ~a32468;
assign a32474 = a19100 & a17968;
assign a32476 = ~a32474 & a32472;
assign a32478 = a32476 & a32466;
assign a32480 = a31866 & a17980;
assign a32482 = a32030 & a31848;
assign a32484 = ~a32482 & ~a32480;
assign a32486 = a31970 & a6702;
assign a32488 = ~a32486 & a32484;
assign a32490 = a31908 & a6696;
assign a32492 = ~a32490 & a32488;
assign a32494 = a32492 & a32478;
assign a32496 = ~a32494 & ~a30468;
assign a32498 = ~a32496 & ~a32456;
assign a32500 = ~a31978 & a30470;
assign a32502 = ~a32500 & a32498;
assign a32504 = ~a32502 & a16292;
assign a32506 = ~a32504 & ~a32454;
assign a32508 = a32502 & ~a16292;
assign a32510 = ~a32508 & ~a32506;
assign a32512 = ~a32176 & a16298;
assign a32514 = ~a32512 & ~a32510;
assign a32516 = ~a32514 & a32180;
assign a32518 = ~a32516 & ~a32074;
assign a32520 = ~a32512 & ~a32128;
assign a32522 = a32228 & ~a16310;
assign a32524 = ~a32522 & ~a32284;
assign a32526 = ~a32524 & ~a32280;
assign a32528 = ~a32526 & ~a32340;
assign a32530 = ~a32528 & ~a32336;
assign a32532 = ~a32530 & ~a32396;
assign a32534 = ~a32532 & ~a32392;
assign a32536 = ~a32534 & ~a32452;
assign a32538 = ~a32536 & ~a32448;
assign a32540 = ~a32538 & ~a32508;
assign a32542 = ~a32540 & ~a32504;
assign a32544 = ~a32542 & ~a32178;
assign a32546 = ~a32544 & a32520;
assign a32550 = l1686 & ~l1664;
assign a32552 = l1686 & ~l1668;
assign a32554 = l1686 & ~l1672;
assign a32556 = l1686 & ~l1676;
assign a32558 = a11700 & ~l1686;
assign a32560 = l1686 & l1682;
assign a32562 = ~a32560 & ~a32558;
assign p0 = ~a6640;

assert property (~p0);

endmodule
