module m6s19 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70;

output p0;

wire na560,a564,a570,a572,a578,a584,a590,a592,a596,a602,a604,na610,na1008,nl478,na1046,
a606,na1048,na1056,na1102,a1104,a1124,a1122,na1128,a1130,a1154,z0,na1164,na1172,na550,a1176,
a1180,a1182,a1184,a1186,a1188,a1190,a1192,a1194,a1196,a1198,z1,z2,z3,na1226,na1228,
na1236,na1330,na1334,a1336,na1346,na1354,a1836,na1844,na1850,na1856,na1862,na1868,na1874,na1880,na1812,
na1830,na1716,na1624,na1532,na1444,z4,na1908,na1910,na1918,na1922,a1924,na1934,na1942,z5,na1970,
na1972,na1980,na1984,a1986,na1996,na2004,z6,na2032,na2034,na2042,na2046,a2048,na2058,na2066,z7,
na2094,na2096,na2104,na2108,a2110,na2120,na2128,z8,na2156,na2158,na2166,na2170,a2172,na2182,na2190,
z9,na2218,na2220,na2228,na2232,a2234,na2244,na2252,a2254,na2432,a2484,z10,na2490,na2496,na2502,
na2508,na2514,na2520,na2526,na2532,na2538,na2544,na2550,na2556,na2562,na2568,na2574,na2580,na2586,na2592,
na2598,na2604,na2610,na2616,na2622,na2628,na2408,na2402,na2394,na2382,na2374,na2364,na2356,na2644,na2656,
na2668,na2680,na2692,na2704,na2716,na2726,a2728,a2712,na2732,a2700,na2736,a2688,na2740,a2676,na2744,
a2664,na2748,a2652,na2752,a2640,na2756,na2762,na2768,na2774,na2780,na2786,na2792,na2798,na2804,na2814,
na2824,na2834,na2844,na2854,na2864,na2874,na2884,na2890,na2896,na2902,na2908,na2914,na2920,na2926,na2932,
a2936,na2940,na2944,na2946,c1,a488,a490,a492,a494,a496,a498,a500,a502,a504,a506,
a508,a510,a512,a514,a516,a518,a520,a522,a524,a526,a528,a530,a532,a534,a536,
a538,a540,a542,a544,a546,a548,a550,a552,a554,a556,a558,a560,a562,a566,a568,
a574,a576,a580,a582,a586,a588,a594,a598,a600,a608,a610,a612,a614,a616,a618,
a620,a622,a624,a626,a628,a630,a632,a634,a636,a638,a640,a642,a644,a646,a648,
a650,a652,a654,a656,a658,a660,a662,a664,a666,a668,a670,a672,a674,a676,a678,
a680,a682,a684,a686,a688,a690,a692,a694,a696,a698,a700,a702,a704,a706,a708,
a710,a712,a714,a716,a718,a720,a722,a724,a726,a728,a730,a732,a734,a736,a738,
a740,a742,a744,a746,a748,a750,a752,a754,a756,a758,a760,a762,a764,a766,a768,
a770,a772,a774,a776,a778,a780,a782,a784,a786,a788,a790,a792,a794,a796,a798,
a800,a802,a804,a806,a808,a810,a812,a814,a816,a818,a820,a822,a824,a826,a828,
a830,a832,a834,a836,a838,a840,a842,a844,a846,a848,a850,a852,a854,a856,a858,
a860,a862,a864,a866,a868,a870,a872,a874,a876,a878,a880,a882,a884,a886,a888,
a890,a892,a894,a896,a898,a900,a902,a904,a906,a908,a910,a912,a914,a916,a918,
a920,a922,a924,a926,a928,a930,a932,a934,a936,a938,a940,a942,a944,a946,a948,
a950,a952,a954,a956,a958,a960,a962,a964,a966,a968,a970,a972,a974,a976,a978,
a980,a982,a984,a986,a988,a990,a992,a994,a996,a998,a1000,a1002,a1004,a1006,a1008,
a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,a1038,
a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,a1062,a1064,a1066,a1068,
a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,a1092,a1094,a1096,a1098,
a1100,a1102,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1126,a1128,a1132,a1134,a1136,
a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,a1156,a1158,a1160,a1162,a1164,a1166,a1168,
a1170,a1172,a1174,a1178,a1200,a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,a1218,a1220,
a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,a1248,a1250,
a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,a1268,a1270,a1272,a1274,a1276,a1278,a1280,
a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,a1310,
a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,a1334,a1338,a1340,a1342,
a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,a1368,a1370,a1372,
a1374,a1376,a1378,a1380,a1382,a1384,a1386,a1388,a1390,a1392,a1394,a1396,a1398,a1400,a1402,
a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1426,a1428,a1430,a1432,
a1434,a1436,a1438,a1440,a1442,a1444,a1446,a1448,a1450,a1452,a1454,a1456,a1458,a1460,a1462,
a1464,a1466,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1482,a1484,a1486,a1488,a1490,a1492,
a1494,a1496,a1498,a1500,a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,a1518,a1520,a1522,
a1524,a1526,a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,a1548,a1550,a1552,
a1554,a1556,a1558,a1560,a1562,a1564,a1566,a1568,a1570,a1572,a1574,a1576,a1578,a1580,a1582,
a1584,a1586,a1588,a1590,a1592,a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,a1610,a1612,
a1614,a1616,a1618,a1620,a1622,a1624,a1626,a1628,a1630,a1632,a1634,a1636,a1638,a1640,a1642,
a1644,a1646,a1648,a1650,a1652,a1654,a1656,a1658,a1660,a1662,a1664,a1666,a1668,a1670,a1672,
a1674,a1676,a1678,a1680,a1682,a1684,a1686,a1688,a1690,a1692,a1694,a1696,a1698,a1700,a1702,
a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,a1732,
a1734,a1736,a1738,a1740,a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,a1758,a1760,a1762,
a1764,a1766,a1768,a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,a1790,a1792,
a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,a1822,
a1824,a1826,a1828,a1830,a1832,a1834,a1838,a1840,a1842,a1844,a1846,a1848,a1850,a1852,a1854,
a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,a1882,a1884,
a1886,a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,a1910,a1912,a1914,
a1916,a1918,a1920,a1922,a1926,a1928,a1930,a1932,a1934,a1936,a1938,a1940,a1942,a1944,a1946,
a1948,a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,a1972,a1974,a1976,
a1978,a1980,a1982,a1984,a1988,a1990,a1992,a1994,a1996,a1998,a2000,a2002,a2004,a2006,a2008,
a2010,a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,a2030,a2032,a2034,a2036,a2038,
a2040,a2042,a2044,a2046,a2050,a2052,a2054,a2056,a2058,a2060,a2062,a2064,a2066,a2068,a2070,
a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,a2090,a2092,a2094,a2096,a2098,a2100,
a2102,a2104,a2106,a2108,a2112,a2114,a2116,a2118,a2120,a2122,a2124,a2126,a2128,a2130,a2132,
a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,a2152,a2154,a2156,a2158,a2160,a2162,
a2164,a2166,a2168,a2170,a2174,a2176,a2178,a2180,a2182,a2184,a2186,a2188,a2190,a2192,a2194,
a2196,a2198,a2200,a2202,a2204,a2206,a2208,a2210,a2212,a2214,a2216,a2218,a2220,a2222,a2224,
a2226,a2228,a2230,a2232,a2236,a2238,a2240,a2242,a2244,a2246,a2248,a2250,a2252,a2256,a2258,
a2260,a2262,a2264,a2266,a2268,a2270,a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,
a2290,a2292,a2294,a2296,a2298,a2300,a2302,a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,
a2320,a2322,a2324,a2326,a2328,a2330,a2332,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,
a2350,a2352,a2354,a2356,a2358,a2360,a2362,a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,
a2380,a2382,a2384,a2386,a2388,a2390,a2392,a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,
a2410,a2412,a2414,a2416,a2418,a2420,a2422,a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,
a2440,a2442,a2444,a2446,a2448,a2450,a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,
a2470,a2472,a2474,a2476,a2478,a2480,a2482,a2486,a2488,a2490,a2492,a2494,a2496,a2498,a2500,
a2502,a2504,a2506,a2508,a2510,a2512,a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2528,a2530,
a2532,a2534,a2536,a2538,a2540,a2542,a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,
a2562,a2564,a2566,a2568,a2570,a2572,a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,
a2592,a2594,a2596,a2598,a2600,a2602,a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,
a2622,a2624,a2626,a2628,a2630,a2632,a2634,a2636,a2638,a2642,a2644,a2646,a2648,a2650,a2654,
a2656,a2658,a2660,a2662,a2666,a2668,a2670,a2672,a2674,a2678,a2680,a2682,a2684,a2686,a2690,
a2692,a2694,a2696,a2698,a2702,a2704,a2706,a2708,a2710,a2714,a2716,a2718,a2720,a2722,a2724,
a2726,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,a2752,a2754,a2756,
a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,a2782,a2784,a2786,
a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,a2810,a2812,a2814,a2816,
a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,a2840,a2842,a2844,a2846,
a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,a2870,a2872,a2874,a2876,
a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,a2900,a2902,a2904,a2906,
a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2930,a2932,a2934,a2938,
a2940,a2942,a2944,a2946,p0;

reg l72,l74,l76,l78,l80,l82,l84,l86,l88,l90,l92,l94,l96,l98,l100,
l102,l104,l106,l108,l110,l112,l114,l116,l118,l120,l122,l124,l126,l128,l130,
l132,l134,l136,l138,l140,l142,l144,l146,l148,l150,l152,l154,l156,l158,l160,
l162,l164,l166,l168,l170,l172,l174,l176,l178,l180,l182,l184,l186,l188,l190,
l192,l194,l196,l198,l200,l202,l204,l206,l208,l210,l212,l214,l216,l218,l220,
l222,l224,l226,l228,l230,l232,l234,l236,l238,l240,l242,l244,l246,l248,l250,
l252,l254,l256,l258,l260,l262,l264,l266,l268,l270,l272,l274,l276,l278,l280,
l282,l284,l286,l288,l290,l292,l294,l296,l298,l300,l302,l304,l306,l308,l310,
l312,l314,l316,l318,l320,l322,l324,l326,l328,l330,l332,l334,l336,l338,l340,
l342,l344,l346,l348,l350,l352,l354,l356,l358,l360,l362,l364,l366,l368,l370,
l372,l374,l376,l378,l380,l382,l384,l386,l388,l390,l392,l394,l396,l398,l400,
l402,l404,l406,l408,l410,l412,l414,l416,l418,l420,l422,l424,l426,l428,l430,
l432,l434,l436,l438,l440,l442,l444,l446,l448,l450,l452,l454,l456,l458,l460,
l462,l464,l466,l468,l470,l472,l474,l476,l478,l480,l482,l484,l486;

initial
begin
   l72 = 0;
   l74 = 0;
   l76 = 0;
   l78 = 0;
   l80 = 0;
   l82 = 0;
   l84 = 0;
   l86 = 0;
   l88 = 0;
   l90 = 0;
   l92 = 0;
   l94 = 0;
   l96 = 0;
   l98 = 0;
   l100 = 0;
   l102 = 0;
   l104 = 0;
   l106 = 0;
   l108 = 0;
   l110 = 0;
   l112 = 0;
   l114 = 0;
   l116 = 0;
   l118 = 0;
   l120 = 0;
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
   l392 = 0;
   l394 = 0;
   l396 = 0;
   l398 = 0;
   l400 = 0;
   l402 = 0;
   l404 = 0;
   l406 = 0;
   l408 = 0;
   l410 = 0;
   l412 = 0;
   l414 = 0;
   l416 = 0;
   l418 = 0;
   l420 = 0;
   l422 = 0;
   l424 = 0;
   l426 = 0;
   l428 = 0;
   l430 = 0;
   l432 = 0;
   l434 = 0;
   l436 = 0;
   l438 = 0;
   l440 = 0;
   l442 = 0;
   l444 = 0;
   l446 = 0;
   l448 = 0;
   l450 = 0;
   l452 = 0;
   l454 = 0;
   l456 = 0;
   l458 = 0;
   l460 = 0;
   l462 = 0;
   l464 = 0;
   l466 = 0;
   l468 = 0;
   l470 = 0;
   l472 = 0;
   l474 = 0;
   l476 = 0;
   l478 = 0;
   l480 = 0;
   l482 = 0;
   l484 = 0;
   l486 = 0;
end

always @(posedge na560)
   l72 <= na560;

always @(posedge a564)
   l74 <= a564;

always @(posedge a570)
   l76 <= a570;

always @(posedge a572)
   l78 <= a572;

always @(posedge a578)
   l80 <= a578;

always @(posedge a584)
   l82 <= a584;

always @(posedge a590)
   l84 <= a590;

always @(posedge a592)
   l86 <= a592;

always @(posedge a596)
   l88 <= a596;

always @(posedge a602)
   l90 <= a602;

always @(posedge a604)
   l92 <= a604;

always @(posedge na610)
   l94 <= na610;

always @(posedge na1008)
   l96 <= na1008;

always @(posedge nl478)
   l98 <= nl478;

always @(posedge na1046)
   l100 <= na1046;

always @(posedge a606)
   l102 <= a606;

always @(posedge na1048)
   l104 <= na1048;

always @(posedge na1056)
   l106 <= na1056;

always @(posedge na1102)
   l108 <= na1102;

always @(posedge a1104)
   l110 <= a1104;

always @(posedge a1124)
   l112 <= a1124;

always @(posedge a1122)
   l114 <= a1122;

always @(posedge na1128)
   l116 <= na1128;

always @(posedge a1130)
   l118 <= a1130;

always @(posedge l122)
   l120 <= l122;

always @(posedge a1154)
   l122 <= a1154;

always @(posedge z0)
   l124 <= z0;

always @(posedge na1164)
   l126 <= na1164;

always @(posedge na1172)
   l128 <= na1172;

always @(posedge na550)
   l130 <= na550;

always @(posedge a1176)
   l132 <= a1176;

always @(posedge a1180)
   l134 <= a1180;

always @(posedge a1182)
   l136 <= a1182;

always @(posedge a1184)
   l138 <= a1184;

always @(posedge a1186)
   l140 <= a1186;

always @(posedge a1188)
   l142 <= a1188;

always @(posedge a1190)
   l144 <= a1190;

always @(posedge a1192)
   l146 <= a1192;

always @(posedge a1194)
   l148 <= a1194;

always @(posedge a1196)
   l150 <= a1196;

always @(posedge a1198)
   l152 <= a1198;

always @(posedge z1)
   l154 <= z1;

always @(posedge z2)
   l156 <= z2;

always @(posedge l162)
   l158 <= l162;

always @(posedge z3)
   l160 <= z3;

always @(posedge na1226)
   l162 <= na1226;

always @(posedge na1228)
   l164 <= na1228;

always @(posedge na1236)
   l166 <= na1236;

always @(posedge na1330)
   l168 <= na1330;

always @(posedge na1334)
   l170 <= na1334;

always @(posedge a1336)
   l172 <= a1336;

always @(posedge na1346)
   l174 <= na1346;

always @(posedge na1354)
   l176 <= na1354;

always @(posedge a1836)
   l178 <= a1836;

always @(posedge na1844)
   l180 <= na1844;

always @(posedge na1850)
   l182 <= na1850;

always @(posedge na1856)
   l184 <= na1856;

always @(posedge na1862)
   l186 <= na1862;

always @(posedge na1868)
   l188 <= na1868;

always @(posedge na1874)
   l190 <= na1874;

always @(posedge na1880)
   l192 <= na1880;

always @(posedge na1812)
   l194 <= na1812;

always @(posedge na1830)
   l196 <= na1830;

always @(posedge na1716)
   l198 <= na1716;

always @(posedge na1624)
   l200 <= na1624;

always @(posedge na1532)
   l202 <= na1532;

always @(posedge na1444)
   l204 <= na1444;

always @(posedge l210)
   l206 <= l210;

always @(posedge z4)
   l208 <= z4;

always @(posedge na1908)
   l210 <= na1908;

always @(posedge na1910)
   l212 <= na1910;

always @(posedge na1918)
   l214 <= na1918;

always @(posedge na1922)
   l216 <= na1922;

always @(posedge a1924)
   l218 <= a1924;

always @(posedge na1934)
   l220 <= na1934;

always @(posedge na1942)
   l222 <= na1942;

always @(posedge l228)
   l224 <= l228;

always @(posedge z5)
   l226 <= z5;

always @(posedge na1970)
   l228 <= na1970;

always @(posedge na1972)
   l230 <= na1972;

always @(posedge na1980)
   l232 <= na1980;

always @(posedge na1984)
   l234 <= na1984;

always @(posedge a1986)
   l236 <= a1986;

always @(posedge na1996)
   l238 <= na1996;

always @(posedge na2004)
   l240 <= na2004;

always @(posedge l246)
   l242 <= l246;

always @(posedge z6)
   l244 <= z6;

always @(posedge na2032)
   l246 <= na2032;

always @(posedge na2034)
   l248 <= na2034;

always @(posedge na2042)
   l250 <= na2042;

always @(posedge na2046)
   l252 <= na2046;

always @(posedge a2048)
   l254 <= a2048;

always @(posedge na2058)
   l256 <= na2058;

always @(posedge na2066)
   l258 <= na2066;

always @(posedge l264)
   l260 <= l264;

always @(posedge z7)
   l262 <= z7;

always @(posedge na2094)
   l264 <= na2094;

always @(posedge na2096)
   l266 <= na2096;

always @(posedge na2104)
   l268 <= na2104;

always @(posedge na2108)
   l270 <= na2108;

always @(posedge a2110)
   l272 <= a2110;

always @(posedge na2120)
   l274 <= na2120;

always @(posedge na2128)
   l276 <= na2128;

always @(posedge l282)
   l278 <= l282;

always @(posedge z8)
   l280 <= z8;

always @(posedge na2156)
   l282 <= na2156;

always @(posedge na2158)
   l284 <= na2158;

always @(posedge na2166)
   l286 <= na2166;

always @(posedge na2170)
   l288 <= na2170;

always @(posedge a2172)
   l290 <= a2172;

always @(posedge na2182)
   l292 <= na2182;

always @(posedge na2190)
   l294 <= na2190;

always @(posedge l300)
   l296 <= l300;

always @(posedge z9)
   l298 <= z9;

always @(posedge na2218)
   l300 <= na2218;

always @(posedge na2220)
   l302 <= na2220;

always @(posedge na2228)
   l304 <= na2228;

always @(posedge na2232)
   l306 <= na2232;

always @(posedge a2234)
   l308 <= a2234;

always @(posedge na2244)
   l310 <= na2244;

always @(posedge na2252)
   l312 <= na2252;

always @(posedge a2254)
   l314 <= a2254;

always @(posedge na2432)
   l316 <= na2432;

always @(posedge a2484)
   l318 <= a2484;

always @(posedge z10)
   l320 <= z10;

always @(posedge na2490)
   l322 <= na2490;

always @(posedge na2496)
   l324 <= na2496;

always @(posedge na2502)
   l326 <= na2502;

always @(posedge na2508)
   l328 <= na2508;

always @(posedge na2514)
   l330 <= na2514;

always @(posedge na2520)
   l332 <= na2520;

always @(posedge na2526)
   l334 <= na2526;

always @(posedge na2532)
   l336 <= na2532;

always @(posedge na2538)
   l338 <= na2538;

always @(posedge na2544)
   l340 <= na2544;

always @(posedge na2550)
   l342 <= na2550;

always @(posedge na2556)
   l344 <= na2556;

always @(posedge na2562)
   l346 <= na2562;

always @(posedge na2568)
   l348 <= na2568;

always @(posedge na2574)
   l350 <= na2574;

always @(posedge na2580)
   l352 <= na2580;

always @(posedge na2586)
   l354 <= na2586;

always @(posedge na2592)
   l356 <= na2592;

always @(posedge na2598)
   l358 <= na2598;

always @(posedge na2604)
   l360 <= na2604;

always @(posedge na2610)
   l362 <= na2610;

always @(posedge na2616)
   l364 <= na2616;

always @(posedge na2622)
   l366 <= na2622;

always @(posedge na2628)
   l368 <= na2628;

always @(posedge na2408)
   l370 <= na2408;

always @(posedge na2402)
   l372 <= na2402;

always @(posedge na2394)
   l374 <= na2394;

always @(posedge na2382)
   l376 <= na2382;

always @(posedge na2374)
   l378 <= na2374;

always @(posedge na2364)
   l380 <= na2364;

always @(posedge na2356)
   l382 <= na2356;

always @(posedge na2644)
   l384 <= na2644;

always @(posedge na2656)
   l386 <= na2656;

always @(posedge na2668)
   l388 <= na2668;

always @(posedge na2680)
   l390 <= na2680;

always @(posedge na2692)
   l392 <= na2692;

always @(posedge na2704)
   l394 <= na2704;

always @(posedge na2716)
   l396 <= na2716;

always @(posedge na2726)
   l398 <= na2726;

always @(posedge a2728)
   l400 <= a2728;

always @(posedge a2712)
   l402 <= a2712;

always @(posedge na2732)
   l404 <= na2732;

always @(posedge a2700)
   l406 <= a2700;

always @(posedge na2736)
   l408 <= na2736;

always @(posedge a2688)
   l410 <= a2688;

always @(posedge na2740)
   l412 <= na2740;

always @(posedge a2676)
   l414 <= a2676;

always @(posedge na2744)
   l416 <= na2744;

always @(posedge a2664)
   l418 <= a2664;

always @(posedge na2748)
   l420 <= na2748;

always @(posedge a2652)
   l422 <= a2652;

always @(posedge na2752)
   l424 <= na2752;

always @(posedge a2640)
   l426 <= a2640;

always @(posedge na2756)
   l428 <= na2756;

always @(posedge na2762)
   l430 <= na2762;

always @(posedge na2768)
   l432 <= na2768;

always @(posedge na2774)
   l434 <= na2774;

always @(posedge na2780)
   l436 <= na2780;

always @(posedge na2786)
   l438 <= na2786;

always @(posedge na2792)
   l440 <= na2792;

always @(posedge na2798)
   l442 <= na2798;

always @(posedge na2804)
   l444 <= na2804;

always @(posedge na2814)
   l446 <= na2814;

always @(posedge na2824)
   l448 <= na2824;

always @(posedge na2834)
   l450 <= na2834;

always @(posedge na2844)
   l452 <= na2844;

always @(posedge na2854)
   l454 <= na2854;

always @(posedge na2864)
   l456 <= na2864;

always @(posedge na2874)
   l458 <= na2874;

always @(posedge na2884)
   l460 <= na2884;

always @(posedge na2890)
   l462 <= na2890;

always @(posedge na2896)
   l464 <= na2896;

always @(posedge na2902)
   l466 <= na2902;

always @(posedge na2908)
   l468 <= na2908;

always @(posedge na2914)
   l470 <= na2914;

always @(posedge na2920)
   l472 <= na2920;

always @(posedge na2926)
   l474 <= na2926;

always @(posedge na2932)
   l476 <= na2932;

always @(posedge a2936)
   l478 <= a2936;

always @(posedge na2940)
   l480 <= na2940;

always @(posedge na2944)
   l482 <= na2944;

always @(posedge na2946)
   l484 <= na2946;

always @(posedge c1)
   l486 <= c1;


assign na560 = ~a560;
assign a564 = a562 & a512;
assign a570 = a568 & ~a566;
assign a572 = a562 & a526;
assign a578 = a576 & a562;
assign a584 = a582 & a562;
assign a590 = a588 & a562;
assign a592 = a562 & ~l86;
assign a596 = a594 & ~a536;
assign a602 = a600 & ~a598;
assign a604 = a562 & ~a508;
assign na610 = ~a610;
assign na1008 = ~a1008;
assign nl478 = ~l478;
assign na1046 = ~a1046;
assign a606 = a550 & l100;
assign na1048 = ~a1048;
assign na1056 = ~a1056;
assign na1102 = ~a1102;
assign a1104 = a1086 & l314;
assign a1124 = ~a1122 & a1106;
assign a1122 = ~a1120 & ~a612;
assign na1128 = ~a1128;
assign a1130 = a1038 & l116;
assign a1154 = a1152 & ~a1150;
assign z0 = l120;
assign na1164 = ~a1164;
assign na1172 = ~a1172;
assign na550 = ~a550;
assign a1176 = a1174 & a1132;
assign a1180 = a1178 & ~i6;
assign a1182 = a1178 & i6;
assign a1184 = l298 & l296;
assign a1186 = l280 & l278;
assign a1188 = l262 & l260;
assign a1190 = l244 & l242;
assign a1192 = l226 & l224;
assign a1194 = l208 & l206;
assign a1196 = l160 & l158;
assign a1198 = l156 & l154;
assign z1 = l100;
assign z2 = l154;
assign z3 = l158;
assign na1226 = ~a1226;
assign na1228 = ~a1228;
assign na1236 = ~a1236;
assign na1330 = ~a1330;
assign na1334 = ~a1334;
assign a1336 = a1218 & l170;
assign na1346 = ~a1346;
assign na1354 = ~a1354;
assign a1836 = ~a1834 & ~a1820;
assign na1844 = ~a1844;
assign na1850 = ~a1850;
assign na1856 = ~a1856;
assign na1862 = ~a1862;
assign na1868 = ~a1868;
assign na1874 = ~a1874;
assign na1880 = ~a1880;
assign na1812 = ~a1812;
assign na1830 = ~a1830;
assign na1716 = ~a1716;
assign na1624 = ~a1624;
assign na1532 = ~a1532;
assign na1444 = ~a1444;
assign z4 = l206;
assign na1908 = ~a1908;
assign na1910 = ~a1910;
assign na1918 = ~a1918;
assign na1922 = ~a1922;
assign a1924 = a1900 & l216;
assign na1934 = ~a1934;
assign na1942 = ~a1942;
assign z5 = l224;
assign na1970 = ~a1970;
assign na1972 = ~a1972;
assign na1980 = ~a1980;
assign na1984 = ~a1984;
assign a1986 = a1962 & l234;
assign na1996 = ~a1996;
assign na2004 = ~a2004;
assign z6 = l242;
assign na2032 = ~a2032;
assign na2034 = ~a2034;
assign na2042 = ~a2042;
assign na2046 = ~a2046;
assign a2048 = a2024 & l252;
assign na2058 = ~a2058;
assign na2066 = ~a2066;
assign z7 = l260;
assign na2094 = ~a2094;
assign na2096 = ~a2096;
assign na2104 = ~a2104;
assign na2108 = ~a2108;
assign a2110 = a2086 & l270;
assign na2120 = ~a2120;
assign na2128 = ~a2128;
assign z8 = l278;
assign na2156 = ~a2156;
assign na2158 = ~a2158;
assign na2166 = ~a2166;
assign na2170 = ~a2170;
assign a2172 = a2148 & l288;
assign na2182 = ~a2182;
assign na2190 = ~a2190;
assign z9 = l296;
assign na2218 = ~a2218;
assign na2220 = ~a2220;
assign na2228 = ~a2228;
assign na2232 = ~a2232;
assign a2234 = a2210 & l306;
assign na2244 = ~a2244;
assign na2252 = ~a2252;
assign a2254 = ~a1090 & ~a1086;
assign na2432 = ~a2432;
assign a2484 = ~a2482 & ~a2414;
assign z10 = l114;
assign na2490 = ~a2490;
assign na2496 = ~a2496;
assign na2502 = ~a2502;
assign na2508 = ~a2508;
assign na2514 = ~a2514;
assign na2520 = ~a2520;
assign na2526 = ~a2526;
assign na2532 = ~a2532;
assign na2538 = ~a2538;
assign na2544 = ~a2544;
assign na2550 = ~a2550;
assign na2556 = ~a2556;
assign na2562 = ~a2562;
assign na2568 = ~a2568;
assign na2574 = ~a2574;
assign na2580 = ~a2580;
assign na2586 = ~a2586;
assign na2592 = ~a2592;
assign na2598 = ~a2598;
assign na2604 = ~a2604;
assign na2610 = ~a2610;
assign na2616 = ~a2616;
assign na2622 = ~a2622;
assign na2628 = ~a2628;
assign na2408 = ~a2408;
assign na2402 = ~a2402;
assign na2394 = ~a2394;
assign na2382 = ~a2382;
assign na2374 = ~a2374;
assign na2364 = ~a2364;
assign na2356 = ~a2356;
assign na2644 = ~a2644;
assign na2656 = ~a2656;
assign na2668 = ~a2668;
assign na2680 = ~a2680;
assign na2692 = ~a2692;
assign na2704 = ~a2704;
assign na2716 = ~a2716;
assign na2726 = ~a2726;
assign a2728 = a2472 & l398;
assign a2712 = a2710 & a2708;
assign na2732 = ~a2732;
assign a2700 = a2698 & a2696;
assign na2736 = ~a2736;
assign a2688 = a2686 & a2684;
assign na2740 = ~a2740;
assign a2676 = a2674 & a2672;
assign na2744 = ~a2744;
assign a2664 = a2662 & a2660;
assign na2748 = ~a2748;
assign a2652 = a2650 & a2648;
assign na2752 = ~a2752;
assign a2640 = a2638 & a2636;
assign na2756 = ~a2756;
assign na2762 = ~a2762;
assign na2768 = ~a2768;
assign na2774 = ~a2774;
assign na2780 = ~a2780;
assign na2786 = ~a2786;
assign na2792 = ~a2792;
assign na2798 = ~a2798;
assign na2804 = ~a2804;
assign na2814 = ~a2814;
assign na2824 = ~a2824;
assign na2834 = ~a2834;
assign na2844 = ~a2844;
assign na2854 = ~a2854;
assign na2864 = ~a2864;
assign na2874 = ~a2874;
assign na2884 = ~a2884;
assign na2890 = ~a2890;
assign na2896 = ~a2896;
assign na2902 = ~a2902;
assign na2908 = ~a2908;
assign na2914 = ~a2914;
assign na2920 = ~a2920;
assign na2926 = ~a2926;
assign na2932 = ~a2932;
assign a2936 = ~a2934 & l480;
assign na2940 = ~a2940;
assign na2944 = ~a2944;
assign na2946 = ~a2946;
assign c1 = 1;
assign a488 = l86 & l84;
assign a490 = a488 & l82;
assign a492 = a490 & l80;
assign a494 = a492 & l78;
assign a496 = a494 & l88;
assign a498 = a496 & l90;
assign a500 = a498 & l76;
assign a502 = a500 & l74;
assign a504 = a502 & ~l92;
assign a506 = ~a502 & l92;
assign a508 = ~a506 & ~a504;
assign a510 = ~a500 & ~l74;
assign a512 = ~a510 & ~a502;
assign a514 = ~a488 & l80;
assign a516 = l94 & ~l82;
assign a518 = l82 & ~l80;
assign a520 = ~a518 & ~a516;
assign a522 = a520 & ~a514;
assign a524 = ~a492 & ~l78;
assign a526 = ~a524 & ~a494;
assign a528 = a526 & ~a522;
assign a530 = l90 & ~l76;
assign a532 = ~a530 & ~a528;
assign a534 = ~a496 & l76;
assign a536 = ~a494 & ~l88;
assign a538 = ~a536 & ~a498;
assign a540 = ~a538 & ~a534;
assign a542 = a540 & a532;
assign a544 = a542 & ~a512;
assign a546 = ~l102 & l100;
assign a548 = ~a546 & l96;
assign a550 = l486 & ~l98;
assign a552 = a550 & ~a548;
assign a554 = a552 & ~l96;
assign a556 = a554 & ~a544;
assign a558 = a556 & ~a508;
assign a560 = ~a558 & ~l72;
assign a562 = a552 & l94;
assign a566 = ~a498 & ~l76;
assign a568 = a562 & ~a500;
assign a574 = ~a490 & ~l80;
assign a576 = ~a574 & ~a492;
assign a580 = ~a488 & ~l82;
assign a582 = ~a580 & ~a490;
assign a586 = ~l86 & ~l84;
assign a588 = ~a586 & ~a488;
assign a594 = a562 & ~a496;
assign a598 = ~a496 & ~l90;
assign a600 = a562 & ~a498;
assign a608 = a606 & ~l102;
assign a610 = ~a608 & ~a562;
assign a612 = l486 & ~l112;
assign a614 = l486 & ~l178;
assign a616 = a614 & l114;
assign a618 = ~a616 & a612;
assign a620 = a618 & l96;
assign a622 = l180 & l138;
assign a624 = l182 & l140;
assign a626 = l184 & l142;
assign a628 = l186 & l152;
assign a630 = l188 & l144;
assign a632 = l190 & l148;
assign a634 = ~l190 & l150;
assign a636 = ~a634 & ~a632;
assign a638 = ~a636 & ~l188;
assign a640 = ~a638 & ~a630;
assign a642 = ~a640 & ~l186;
assign a644 = ~a642 & ~a628;
assign a646 = ~a644 & ~l184;
assign a648 = ~a646 & ~a626;
assign a650 = ~a648 & ~l182;
assign a652 = ~a650 & ~a624;
assign a654 = ~a652 & ~l180;
assign a656 = ~a654 & ~a622;
assign a658 = a656 & ~l146;
assign a660 = l180 & l152;
assign a662 = l182 & l144;
assign a664 = l184 & l148;
assign a666 = l186 & l150;
assign a668 = l188 & l138;
assign a670 = l190 & l140;
assign a672 = ~l190 & l142;
assign a674 = ~a672 & ~a670;
assign a676 = ~a674 & ~l188;
assign a678 = ~a676 & ~a668;
assign a680 = ~a678 & ~l186;
assign a682 = ~a680 & ~a666;
assign a684 = ~a682 & ~l184;
assign a686 = ~a684 & ~a664;
assign a688 = ~a686 & ~l182;
assign a690 = ~a688 & ~a662;
assign a692 = ~a690 & ~l180;
assign a694 = ~a692 & ~a660;
assign a696 = l180 & l144;
assign a698 = l182 & l148;
assign a700 = l184 & l150;
assign a702 = l186 & l138;
assign a704 = l188 & l140;
assign a706 = l190 & l142;
assign a708 = ~l190 & l152;
assign a710 = ~a708 & ~a706;
assign a712 = ~a710 & ~l188;
assign a714 = ~a712 & ~a704;
assign a716 = ~a714 & ~l186;
assign a718 = ~a716 & ~a702;
assign a720 = ~a718 & ~l184;
assign a722 = ~a720 & ~a700;
assign a724 = ~a722 & ~l182;
assign a726 = ~a724 & ~a698;
assign a728 = ~a726 & ~l180;
assign a730 = ~a728 & ~a696;
assign a732 = l180 & l150;
assign a734 = l182 & l138;
assign a736 = l184 & l140;
assign a738 = l186 & l142;
assign a740 = l188 & l152;
assign a742 = l190 & l144;
assign a744 = ~l190 & l148;
assign a746 = ~a744 & ~a742;
assign a748 = ~a746 & ~l188;
assign a750 = ~a748 & ~a740;
assign a752 = ~a750 & ~l186;
assign a754 = ~a752 & ~a738;
assign a756 = ~a754 & ~l184;
assign a758 = ~a756 & ~a736;
assign a760 = ~a758 & ~l182;
assign a762 = ~a760 & ~a734;
assign a764 = ~a762 & ~l180;
assign a766 = ~a764 & ~a732;
assign a768 = l180 & l148;
assign a770 = l182 & l150;
assign a772 = l184 & l138;
assign a774 = l186 & l140;
assign a776 = l188 & l142;
assign a778 = l190 & l152;
assign a780 = ~l190 & l144;
assign a782 = ~a780 & ~a778;
assign a784 = ~a782 & ~l188;
assign a786 = ~a784 & ~a776;
assign a788 = ~a786 & ~l186;
assign a790 = ~a788 & ~a774;
assign a792 = ~a790 & ~l184;
assign a794 = ~a792 & ~a772;
assign a796 = ~a794 & ~l182;
assign a798 = ~a796 & ~a770;
assign a800 = ~a798 & ~l180;
assign a802 = ~a800 & ~a768;
assign a804 = a802 & a766;
assign a806 = a804 & a730;
assign a808 = a806 & ~a694;
assign a810 = a808 & a658;
assign a812 = a810 & l180;
assign a814 = l180 & l142;
assign a816 = l182 & l152;
assign a818 = l184 & l144;
assign a820 = l186 & l148;
assign a822 = l188 & l150;
assign a824 = l190 & l138;
assign a826 = ~l190 & l140;
assign a828 = ~a826 & ~a824;
assign a830 = ~a828 & ~l188;
assign a832 = ~a830 & ~a822;
assign a834 = ~a832 & ~l186;
assign a836 = ~a834 & ~a820;
assign a838 = ~a836 & ~l184;
assign a840 = ~a838 & ~a818;
assign a842 = ~a840 & ~l182;
assign a844 = ~a842 & ~a816;
assign a846 = ~a844 & ~l180;
assign a848 = ~a846 & ~a814;
assign a850 = a806 & a694;
assign a852 = a850 & ~a848;
assign a854 = a852 & a658;
assign a856 = a854 & l182;
assign a858 = l180 & l140;
assign a860 = l182 & l142;
assign a862 = l184 & l152;
assign a864 = l186 & l144;
assign a866 = l188 & l148;
assign a868 = l190 & l150;
assign a870 = ~l190 & l138;
assign a872 = ~a870 & ~a868;
assign a874 = ~a872 & ~l188;
assign a876 = ~a874 & ~a866;
assign a878 = ~a876 & ~l186;
assign a880 = ~a878 & ~a864;
assign a882 = ~a880 & ~l184;
assign a884 = ~a882 & ~a862;
assign a886 = ~a884 & ~l182;
assign a888 = ~a886 & ~a860;
assign a890 = ~a888 & ~l180;
assign a892 = ~a890 & ~a858;
assign a894 = a850 & a848;
assign a896 = a894 & ~a892;
assign a898 = a896 & a658;
assign a900 = a898 & l184;
assign a902 = ~a656 & l186;
assign a904 = a902 & ~l146;
assign a906 = ~a766 & a658;
assign a908 = a906 & l188;
assign a910 = ~a802 & a766;
assign a912 = a910 & a658;
assign a914 = a912 & l190;
assign a916 = a804 & ~a730;
assign a918 = a916 & a658;
assign a920 = a918 & ~l190;
assign a922 = ~a920 & ~a914;
assign a924 = ~a922 & ~l188;
assign a926 = ~a924 & ~a908;
assign a928 = ~a926 & ~l186;
assign a930 = ~a928 & ~a904;
assign a932 = ~a930 & ~l184;
assign a934 = ~a932 & ~a900;
assign a936 = ~a934 & ~l182;
assign a938 = ~a936 & ~a856;
assign a940 = ~a938 & ~l180;
assign a942 = ~a940 & ~a812;
assign a944 = ~a614 & l114;
assign a946 = a944 & ~a942;
assign a948 = ~a946 & ~a620;
assign a950 = a656 & l180;
assign a952 = a950 & a808;
assign a954 = a656 & l182;
assign a956 = a954 & a852;
assign a958 = a656 & l184;
assign a960 = a958 & a896;
assign a962 = a656 & l188;
assign a964 = a962 & ~a766;
assign a966 = a656 & l190;
assign a968 = a966 & a910;
assign a970 = a808 & a656;
assign a972 = l486 & ~l192;
assign a974 = a972 & a970;
assign a976 = a916 & a656;
assign a978 = a976 & ~a972;
assign a980 = ~a978 & ~a974;
assign a982 = ~a980 & ~l190;
assign a984 = ~a982 & ~a968;
assign a986 = ~a984 & ~l188;
assign a988 = ~a986 & ~a964;
assign a990 = ~a988 & ~l186;
assign a992 = ~a990 & ~a902;
assign a994 = ~a992 & ~l184;
assign a996 = ~a994 & ~a960;
assign a998 = ~a996 & ~l182;
assign a1000 = ~a998 & ~a956;
assign a1002 = ~a1000 & ~l180;
assign a1004 = ~a1002 & ~a952;
assign a1006 = ~a1004 & a616;
assign a1008 = ~a1006 & a948;
assign a1010 = ~l124 & ~l122;
assign a1012 = a1010 & ~l120;
assign a1014 = a1012 & l126;
assign a1016 = a612 & ~l110;
assign a1018 = a1016 & ~l114;
assign a1020 = a1018 & ~l108;
assign a1022 = a1020 & l96;
assign a1024 = ~a1022 & a1014;
assign a1026 = ~a1024 & ~l118;
assign a1028 = ~l116 & ~l106;
assign a1030 = ~l118 & ~l104;
assign a1032 = ~a1030 & a1028;
assign a1034 = a1022 & l106;
assign a1036 = ~a1034 & ~a1032;
assign a1038 = ~a1022 & ~l106;
assign a1040 = a1038 & l104;
assign a1042 = ~a1040 & ~a1036;
assign a1044 = ~a1042 & l100;
assign a1046 = ~a1044 & a1026;
assign a1048 = ~a1040 & ~l118;
assign a1050 = a1012 & l128;
assign a1052 = a1050 & a1022;
assign a1054 = ~a1052 & l106;
assign a1056 = ~a1054 & ~a1024;
assign a1058 = l198 & l140;
assign a1060 = l194 & l138;
assign a1062 = ~a1060 & ~a1058;
assign a1064 = l202 & l148;
assign a1066 = l152 & l96;
assign a1068 = ~a1066 & ~a1064;
assign a1070 = a1068 & a1062;
assign a1072 = l168 & l150;
assign a1074 = l200 & l142;
assign a1076 = ~a1074 & ~a1072;
assign a1078 = l196 & l146;
assign a1080 = l204 & l144;
assign a1082 = ~a1080 & ~a1078;
assign a1084 = a1082 & a1076;
assign a1086 = a1084 & a1070;
assign a1088 = a1086 & l108;
assign a1090 = ~l314 & ~l108;
assign a1092 = a1090 & ~l320;
assign a1094 = a1092 & a1018;
assign a1096 = a1094 & ~l318;
assign a1098 = a1096 & a1086;
assign a1100 = a1098 & l316;
assign a1102 = ~a1100 & ~a1088;
assign a1106 = ~a1016 & ~l114;
assign a1108 = ~l140 & ~l138;
assign a1110 = ~l144 & ~l142;
assign a1112 = a1110 & a1108;
assign a1114 = ~l148 & ~l146;
assign a1116 = ~l152 & ~l150;
assign a1118 = a1116 & a1114;
assign a1120 = a1118 & a1112;
assign a1126 = ~a1038 & l116;
assign a1128 = ~a1126 & ~a1034;
assign a1132 = i6 & i4;
assign a1134 = a1132 & ~l132;
assign a1136 = l134 & ~i6;
assign a1138 = l136 & i6;
assign a1140 = ~a1138 & ~i4;
assign a1142 = a1140 & ~a1136;
assign a1144 = ~a1142 & ~a1134;
assign a1146 = ~i6 & i4;
assign a1148 = ~a1146 & ~i8;
assign a1150 = a1148 & a1144;
assign a1152 = ~a550 & ~l130;
assign a1156 = a1012 & ~l128;
assign a1158 = a1156 & i2;
assign a1160 = a1050 & ~a1024;
assign a1162 = a1160 & l126;
assign a1164 = ~a1162 & ~a1158;
assign a1166 = ~a1158 & ~a1024;
assign a1168 = a1048 & a1032;
assign a1170 = ~a1168 & a1160;
assign a1172 = ~a1170 & a1166;
assign a1174 = a1152 & ~i8;
assign a1178 = a1174 & ~i4;
assign a1200 = a1012 & l174;
assign a1202 = a1020 & l168;
assign a1204 = ~a1202 & a1200;
assign a1206 = ~a1204 & ~l172;
assign a1208 = ~l170 & ~l166;
assign a1210 = ~l172 & ~l164;
assign a1212 = ~a1210 & a1208;
assign a1214 = a1202 & l166;
assign a1216 = ~a1214 & ~a1212;
assign a1218 = ~a1202 & ~l166;
assign a1220 = a1218 & l164;
assign a1222 = ~a1220 & ~a1216;
assign a1224 = ~a1222 & l162;
assign a1226 = ~a1224 & a1206;
assign a1228 = ~a1220 & ~l172;
assign a1230 = a1012 & l176;
assign a1232 = a1230 & a1202;
assign a1234 = ~a1232 & l166;
assign a1236 = ~a1234 & ~a1204;
assign a1238 = a618 & l168;
assign a1240 = a950 & ~a766;
assign a1242 = a954 & a910;
assign a1244 = a958 & a916;
assign a1246 = a656 & l186;
assign a1248 = a1246 & a808;
assign a1250 = a962 & a852;
assign a1252 = a966 & a896;
assign a1254 = ~a766 & a656;
assign a1256 = a1254 & a972;
assign a1258 = ~a972 & ~a656;
assign a1260 = ~a1258 & ~a1256;
assign a1262 = ~a1260 & ~l190;
assign a1264 = ~a1262 & ~a1252;
assign a1266 = ~a1264 & ~l188;
assign a1268 = ~a1266 & ~a1250;
assign a1270 = ~a1268 & ~l186;
assign a1272 = ~a1270 & ~a1248;
assign a1274 = ~a1272 & ~l184;
assign a1276 = ~a1274 & ~a1244;
assign a1278 = ~a1276 & ~l182;
assign a1280 = ~a1278 & ~a1242;
assign a1282 = ~a1280 & ~l180;
assign a1284 = ~a1282 & ~a1240;
assign a1286 = ~a1284 & a616;
assign a1288 = ~a1286 & ~a1238;
assign a1290 = a906 & l180;
assign a1292 = a912 & l182;
assign a1294 = a918 & l184;
assign a1296 = a810 & l186;
assign a1298 = a854 & l188;
assign a1300 = a898 & l190;
assign a1302 = ~a656 & ~l146;
assign a1304 = a1302 & ~l190;
assign a1306 = ~a1304 & ~a1300;
assign a1308 = ~a1306 & ~l188;
assign a1310 = ~a1308 & ~a1298;
assign a1312 = ~a1310 & ~l186;
assign a1314 = ~a1312 & ~a1296;
assign a1316 = ~a1314 & ~l184;
assign a1318 = ~a1316 & ~a1294;
assign a1320 = ~a1318 & ~l182;
assign a1322 = ~a1320 & ~a1292;
assign a1324 = ~a1322 & ~l180;
assign a1326 = ~a1324 & ~a1290;
assign a1328 = ~a1326 & a944;
assign a1330 = ~a1328 & a1288;
assign a1332 = ~a1218 & l170;
assign a1334 = ~a1332 & ~a1214;
assign a1338 = a1012 & ~l176;
assign a1340 = a1338 & i10;
assign a1342 = a1230 & ~a1204;
assign a1344 = a1342 & l174;
assign a1346 = ~a1344 & ~a1340;
assign a1348 = ~a1340 & ~a1204;
assign a1350 = a1228 & a1212;
assign a1352 = ~a1350 & a1342;
assign a1354 = ~a1352 & a1348;
assign a1356 = a618 & l204;
assign a1358 = a918 & l180;
assign a1360 = a810 & l182;
assign a1362 = a854 & l184;
assign a1364 = a898 & l186;
assign a1366 = ~a656 & l188;
assign a1368 = a1366 & ~l146;
assign a1370 = a906 & l190;
assign a1372 = a912 & ~l190;
assign a1374 = ~a1372 & ~a1370;
assign a1376 = ~a1374 & ~l188;
assign a1378 = ~a1376 & ~a1368;
assign a1380 = ~a1378 & ~l186;
assign a1382 = ~a1380 & ~a1364;
assign a1384 = ~a1382 & ~l184;
assign a1386 = ~a1384 & ~a1362;
assign a1388 = ~a1386 & ~l182;
assign a1390 = ~a1388 & ~a1360;
assign a1392 = ~a1390 & ~l180;
assign a1394 = ~a1392 & ~a1358;
assign a1396 = ~a1394 & a944;
assign a1398 = ~a1396 & ~a1356;
assign a1400 = a950 & a916;
assign a1402 = a954 & a808;
assign a1404 = a958 & a852;
assign a1406 = a1246 & a896;
assign a1408 = a966 & ~a766;
assign a1410 = a976 & a972;
assign a1412 = a910 & a656;
assign a1414 = a1412 & ~a972;
assign a1416 = ~a1414 & ~a1410;
assign a1418 = ~a1416 & ~l190;
assign a1420 = ~a1418 & ~a1408;
assign a1422 = ~a1420 & ~l188;
assign a1424 = ~a1422 & ~a1366;
assign a1426 = ~a1424 & ~l186;
assign a1428 = ~a1426 & ~a1406;
assign a1430 = ~a1428 & ~l184;
assign a1432 = ~a1430 & ~a1404;
assign a1434 = ~a1432 & ~l182;
assign a1436 = ~a1434 & ~a1402;
assign a1438 = ~a1436 & ~l180;
assign a1440 = ~a1438 & ~a1400;
assign a1442 = ~a1440 & a616;
assign a1444 = ~a1442 & a1398;
assign a1446 = a618 & l202;
assign a1448 = a912 & l180;
assign a1450 = a918 & l182;
assign a1452 = a810 & l184;
assign a1454 = a854 & l186;
assign a1456 = a898 & l188;
assign a1458 = ~a656 & l190;
assign a1460 = a1458 & ~l146;
assign a1462 = a906 & ~l190;
assign a1464 = ~a1462 & ~a1460;
assign a1466 = ~a1464 & ~l188;
assign a1468 = ~a1466 & ~a1456;
assign a1470 = ~a1468 & ~l186;
assign a1472 = ~a1470 & ~a1454;
assign a1474 = ~a1472 & ~l184;
assign a1476 = ~a1474 & ~a1452;
assign a1478 = ~a1476 & ~l182;
assign a1480 = ~a1478 & ~a1450;
assign a1482 = ~a1480 & ~l180;
assign a1484 = ~a1482 & ~a1448;
assign a1486 = ~a1484 & a944;
assign a1488 = ~a1486 & ~a1446;
assign a1490 = a950 & a910;
assign a1492 = a954 & a916;
assign a1494 = a958 & a808;
assign a1496 = a1246 & a852;
assign a1498 = a962 & a896;
assign a1500 = a1412 & a972;
assign a1502 = a1254 & ~a972;
assign a1504 = ~a1502 & ~a1500;
assign a1506 = ~a1504 & ~l190;
assign a1508 = ~a1506 & ~a1458;
assign a1510 = ~a1508 & ~l188;
assign a1512 = ~a1510 & ~a1498;
assign a1514 = ~a1512 & ~l186;
assign a1516 = ~a1514 & ~a1496;
assign a1518 = ~a1516 & ~l184;
assign a1520 = ~a1518 & ~a1494;
assign a1522 = ~a1520 & ~l182;
assign a1524 = ~a1522 & ~a1492;
assign a1526 = ~a1524 & ~l180;
assign a1528 = ~a1526 & ~a1490;
assign a1530 = ~a1528 & a616;
assign a1532 = ~a1530 & a1488;
assign a1534 = a1532 & a1444;
assign a1536 = a618 & l200;
assign a1538 = a854 & l180;
assign a1540 = a898 & l182;
assign a1542 = ~a656 & l184;
assign a1544 = a1542 & ~l146;
assign a1546 = a906 & l186;
assign a1548 = a912 & l188;
assign a1550 = a918 & l190;
assign a1552 = a810 & ~l190;
assign a1554 = ~a1552 & ~a1550;
assign a1556 = ~a1554 & ~l188;
assign a1558 = ~a1556 & ~a1548;
assign a1560 = ~a1558 & ~l186;
assign a1562 = ~a1560 & ~a1546;
assign a1564 = ~a1562 & ~l184;
assign a1566 = ~a1564 & ~a1544;
assign a1568 = ~a1566 & ~l182;
assign a1570 = ~a1568 & ~a1540;
assign a1572 = ~a1570 & ~l180;
assign a1574 = ~a1572 & ~a1538;
assign a1576 = ~a1574 & a944;
assign a1578 = ~a1576 & ~a1536;
assign a1580 = a950 & a852;
assign a1582 = a954 & a896;
assign a1584 = a1246 & ~a766;
assign a1586 = a962 & a910;
assign a1588 = a966 & a916;
assign a1590 = a852 & a656;
assign a1592 = a1590 & a972;
assign a1594 = ~a972 & a970;
assign a1596 = ~a1594 & ~a1592;
assign a1598 = ~a1596 & ~l190;
assign a1600 = ~a1598 & ~a1588;
assign a1602 = ~a1600 & ~l188;
assign a1604 = ~a1602 & ~a1586;
assign a1606 = ~a1604 & ~l186;
assign a1608 = ~a1606 & ~a1584;
assign a1610 = ~a1608 & ~l184;
assign a1612 = ~a1610 & ~a1542;
assign a1614 = ~a1612 & ~l182;
assign a1616 = ~a1614 & ~a1582;
assign a1618 = ~a1616 & ~l180;
assign a1620 = ~a1618 & ~a1580;
assign a1622 = ~a1620 & a616;
assign a1624 = ~a1622 & a1578;
assign a1626 = a1624 & a1534;
assign a1628 = a618 & l198;
assign a1630 = a898 & l180;
assign a1632 = ~a656 & l182;
assign a1634 = a1632 & ~l146;
assign a1636 = a906 & l184;
assign a1638 = a912 & l186;
assign a1640 = a918 & l188;
assign a1642 = a810 & l190;
assign a1644 = a854 & ~l190;
assign a1646 = ~a1644 & ~a1642;
assign a1648 = ~a1646 & ~l188;
assign a1650 = ~a1648 & ~a1640;
assign a1652 = ~a1650 & ~l186;
assign a1654 = ~a1652 & ~a1638;
assign a1656 = ~a1654 & ~l184;
assign a1658 = ~a1656 & ~a1636;
assign a1660 = ~a1658 & ~l182;
assign a1662 = ~a1660 & ~a1634;
assign a1664 = ~a1662 & ~l180;
assign a1666 = ~a1664 & ~a1630;
assign a1668 = ~a1666 & a944;
assign a1670 = ~a1668 & ~a1628;
assign a1672 = a950 & a896;
assign a1674 = a958 & ~a766;
assign a1676 = a1246 & a910;
assign a1678 = a962 & a916;
assign a1680 = a966 & a808;
assign a1682 = a896 & a656;
assign a1684 = a1682 & a972;
assign a1686 = a1590 & ~a972;
assign a1688 = ~a1686 & ~a1684;
assign a1690 = ~a1688 & ~l190;
assign a1692 = ~a1690 & ~a1680;
assign a1694 = ~a1692 & ~l188;
assign a1696 = ~a1694 & ~a1678;
assign a1698 = ~a1696 & ~l186;
assign a1700 = ~a1698 & ~a1676;
assign a1702 = ~a1700 & ~l184;
assign a1704 = ~a1702 & ~a1674;
assign a1706 = ~a1704 & ~l182;
assign a1708 = ~a1706 & ~a1632;
assign a1710 = ~a1708 & ~l180;
assign a1712 = ~a1710 & ~a1672;
assign a1714 = ~a1712 & a616;
assign a1716 = ~a1714 & a1670;
assign a1718 = a1716 & a1626;
assign a1720 = a1330 & a1008;
assign a1722 = a618 & l194;
assign a1724 = a1302 & l180;
assign a1726 = a906 & l182;
assign a1728 = a912 & l184;
assign a1730 = a918 & l186;
assign a1732 = a810 & l188;
assign a1734 = a854 & l190;
assign a1736 = a898 & ~l190;
assign a1738 = ~a1736 & ~a1734;
assign a1740 = ~a1738 & ~l188;
assign a1742 = ~a1740 & ~a1732;
assign a1744 = ~a1742 & ~l186;
assign a1746 = ~a1744 & ~a1730;
assign a1748 = ~a1746 & ~l184;
assign a1750 = ~a1748 & ~a1728;
assign a1752 = ~a1750 & ~l182;
assign a1754 = ~a1752 & ~a1726;
assign a1756 = ~a1754 & ~l180;
assign a1758 = ~a1756 & ~a1724;
assign a1760 = ~a1758 & a944;
assign a1762 = ~a1760 & ~a1722;
assign a1764 = a954 & ~a766;
assign a1766 = a958 & a910;
assign a1768 = a1246 & a916;
assign a1770 = a962 & a808;
assign a1772 = a966 & a852;
assign a1774 = a656 & l146;
assign a1776 = a1774 & a892;
assign a1778 = a1776 & a894;
assign a1780 = a1778 & a972;
assign a1782 = a1682 & ~a972;
assign a1784 = ~a1782 & ~a1780;
assign a1786 = ~a1784 & ~l190;
assign a1788 = ~a1786 & ~a1772;
assign a1790 = ~a1788 & ~l188;
assign a1792 = ~a1790 & ~a1770;
assign a1794 = ~a1792 & ~l186;
assign a1796 = ~a1794 & ~a1768;
assign a1798 = ~a1796 & ~l184;
assign a1800 = ~a1798 & ~a1766;
assign a1802 = ~a1800 & ~l182;
assign a1804 = ~a1802 & ~a1764;
assign a1806 = ~a1804 & ~l180;
assign a1808 = ~a1806 & ~a622;
assign a1810 = ~a1808 & a616;
assign a1812 = ~a1810 & a1762;
assign a1814 = a1812 & a1720;
assign a1816 = a1814 & a1718;
assign a1818 = ~a1816 & l114;
assign a1820 = ~a1818 & a614;
assign a1822 = a618 & l196;
assign a1824 = a944 & l146;
assign a1826 = ~a1824 & ~a1822;
assign a1828 = a1778 & a616;
assign a1830 = ~a1828 & a1826;
assign a1832 = ~a1830 & ~l110;
assign a1834 = a1832 & l114;
assign a1838 = ~a1832 & a1818;
assign a1840 = a1838 & ~a1716;
assign a1842 = ~a1838 & l180;
assign a1844 = ~a1842 & ~a1840;
assign a1846 = a1838 & ~a1624;
assign a1848 = ~a1838 & l182;
assign a1850 = ~a1848 & ~a1846;
assign a1852 = a1838 & ~a1008;
assign a1854 = ~a1838 & l184;
assign a1856 = ~a1854 & ~a1852;
assign a1858 = a1838 & ~a1444;
assign a1860 = ~a1838 & l186;
assign a1862 = ~a1860 & ~a1858;
assign a1864 = a1838 & ~a1532;
assign a1866 = ~a1838 & l188;
assign a1868 = ~a1866 & ~a1864;
assign a1870 = a1838 & ~a1330;
assign a1872 = ~a1838 & l190;
assign a1874 = ~a1872 & ~a1870;
assign a1876 = ~a1838 & ~a972;
assign a1878 = a1838 & ~a1812;
assign a1880 = ~a1878 & ~a1876;
assign a1882 = a1012 & l220;
assign a1884 = a1020 & l202;
assign a1886 = ~a1884 & a1882;
assign a1888 = ~a1886 & ~l218;
assign a1890 = ~l216 & ~l214;
assign a1892 = ~l218 & ~l212;
assign a1894 = ~a1892 & a1890;
assign a1896 = a1884 & l214;
assign a1898 = ~a1896 & ~a1894;
assign a1900 = ~a1884 & ~l214;
assign a1902 = a1900 & l212;
assign a1904 = ~a1902 & ~a1898;
assign a1906 = ~a1904 & l210;
assign a1908 = ~a1906 & a1888;
assign a1910 = ~a1902 & ~l218;
assign a1912 = a1012 & l222;
assign a1914 = a1912 & a1884;
assign a1916 = ~a1914 & l214;
assign a1918 = ~a1916 & ~a1886;
assign a1920 = ~a1900 & l216;
assign a1922 = ~a1920 & ~a1896;
assign a1926 = a1012 & ~l222;
assign a1928 = a1926 & i12;
assign a1930 = a1912 & ~a1886;
assign a1932 = a1930 & l220;
assign a1934 = ~a1932 & ~a1928;
assign a1936 = ~a1928 & ~a1886;
assign a1938 = a1910 & a1894;
assign a1940 = ~a1938 & a1930;
assign a1942 = ~a1940 & a1936;
assign a1944 = a1012 & l238;
assign a1946 = a1020 & l196;
assign a1948 = ~a1946 & a1944;
assign a1950 = ~a1948 & ~l236;
assign a1952 = ~l234 & ~l232;
assign a1954 = ~l236 & ~l230;
assign a1956 = ~a1954 & a1952;
assign a1958 = a1946 & l232;
assign a1960 = ~a1958 & ~a1956;
assign a1962 = ~a1946 & ~l232;
assign a1964 = a1962 & l230;
assign a1966 = ~a1964 & ~a1960;
assign a1968 = ~a1966 & l228;
assign a1970 = ~a1968 & a1950;
assign a1972 = ~a1964 & ~l236;
assign a1974 = a1012 & l240;
assign a1976 = a1974 & a1946;
assign a1978 = ~a1976 & l232;
assign a1980 = ~a1978 & ~a1948;
assign a1982 = ~a1962 & l234;
assign a1984 = ~a1982 & ~a1958;
assign a1988 = a1012 & ~l240;
assign a1990 = a1988 & i14;
assign a1992 = a1974 & ~a1948;
assign a1994 = a1992 & l238;
assign a1996 = ~a1994 & ~a1990;
assign a1998 = ~a1990 & ~a1948;
assign a2000 = a1972 & a1956;
assign a2002 = ~a2000 & a1992;
assign a2004 = ~a2002 & a1998;
assign a2006 = a1012 & l256;
assign a2008 = a1020 & l204;
assign a2010 = ~a2008 & a2006;
assign a2012 = ~a2010 & ~l254;
assign a2014 = ~l252 & ~l250;
assign a2016 = ~l254 & ~l248;
assign a2018 = ~a2016 & a2014;
assign a2020 = a2008 & l250;
assign a2022 = ~a2020 & ~a2018;
assign a2024 = ~a2008 & ~l250;
assign a2026 = a2024 & l248;
assign a2028 = ~a2026 & ~a2022;
assign a2030 = ~a2028 & l246;
assign a2032 = ~a2030 & a2012;
assign a2034 = ~a2026 & ~l254;
assign a2036 = a1012 & l258;
assign a2038 = a2036 & a2008;
assign a2040 = ~a2038 & l250;
assign a2042 = ~a2040 & ~a2010;
assign a2044 = ~a2024 & l252;
assign a2046 = ~a2044 & ~a2020;
assign a2050 = a1012 & ~l258;
assign a2052 = a2050 & i16;
assign a2054 = a2036 & ~a2010;
assign a2056 = a2054 & l256;
assign a2058 = ~a2056 & ~a2052;
assign a2060 = ~a2052 & ~a2010;
assign a2062 = a2034 & a2018;
assign a2064 = ~a2062 & a2054;
assign a2066 = ~a2064 & a2060;
assign a2068 = a1012 & l274;
assign a2070 = a1020 & l200;
assign a2072 = ~a2070 & a2068;
assign a2074 = ~a2072 & ~l272;
assign a2076 = ~l270 & ~l268;
assign a2078 = ~l272 & ~l266;
assign a2080 = ~a2078 & a2076;
assign a2082 = a2070 & l268;
assign a2084 = ~a2082 & ~a2080;
assign a2086 = ~a2070 & ~l268;
assign a2088 = a2086 & l266;
assign a2090 = ~a2088 & ~a2084;
assign a2092 = ~a2090 & l264;
assign a2094 = ~a2092 & a2074;
assign a2096 = ~a2088 & ~l272;
assign a2098 = a1012 & l276;
assign a2100 = a2098 & a2070;
assign a2102 = ~a2100 & l268;
assign a2104 = ~a2102 & ~a2072;
assign a2106 = ~a2086 & l270;
assign a2108 = ~a2106 & ~a2082;
assign a2112 = a1012 & ~l276;
assign a2114 = a2112 & i18;
assign a2116 = a2098 & ~a2072;
assign a2118 = a2116 & l274;
assign a2120 = ~a2118 & ~a2114;
assign a2122 = ~a2114 & ~a2072;
assign a2124 = a2096 & a2080;
assign a2126 = ~a2124 & a2116;
assign a2128 = ~a2126 & a2122;
assign a2130 = a1012 & l292;
assign a2132 = a1020 & l198;
assign a2134 = ~a2132 & a2130;
assign a2136 = ~a2134 & ~l290;
assign a2138 = ~l288 & ~l286;
assign a2140 = ~l290 & ~l284;
assign a2142 = ~a2140 & a2138;
assign a2144 = a2132 & l286;
assign a2146 = ~a2144 & ~a2142;
assign a2148 = ~a2132 & ~l286;
assign a2150 = a2148 & l284;
assign a2152 = ~a2150 & ~a2146;
assign a2154 = ~a2152 & l282;
assign a2156 = ~a2154 & a2136;
assign a2158 = ~a2150 & ~l290;
assign a2160 = a1012 & l294;
assign a2162 = a2160 & a2132;
assign a2164 = ~a2162 & l286;
assign a2166 = ~a2164 & ~a2134;
assign a2168 = ~a2148 & l288;
assign a2170 = ~a2168 & ~a2144;
assign a2174 = a1012 & ~l294;
assign a2176 = a2174 & i20;
assign a2178 = a2160 & ~a2134;
assign a2180 = a2178 & l292;
assign a2182 = ~a2180 & ~a2176;
assign a2184 = ~a2176 & ~a2134;
assign a2186 = a2158 & a2142;
assign a2188 = ~a2186 & a2178;
assign a2190 = ~a2188 & a2184;
assign a2192 = a1012 & l310;
assign a2194 = a1020 & l194;
assign a2196 = ~a2194 & a2192;
assign a2198 = ~a2196 & ~l308;
assign a2200 = ~l306 & ~l304;
assign a2202 = ~l308 & ~l302;
assign a2204 = ~a2202 & a2200;
assign a2206 = a2194 & l304;
assign a2208 = ~a2206 & ~a2204;
assign a2210 = ~a2194 & ~l304;
assign a2212 = a2210 & l302;
assign a2214 = ~a2212 & ~a2208;
assign a2216 = ~a2214 & l300;
assign a2218 = ~a2216 & a2198;
assign a2220 = ~a2212 & ~l308;
assign a2222 = a1012 & l312;
assign a2224 = a2222 & a2194;
assign a2226 = ~a2224 & l304;
assign a2228 = ~a2226 & ~a2196;
assign a2230 = ~a2210 & l306;
assign a2232 = ~a2230 & ~a2206;
assign a2236 = a1012 & ~l312;
assign a2238 = a2236 & i22;
assign a2240 = a2222 & ~a2196;
assign a2242 = a2240 & l310;
assign a2244 = ~a2242 & ~a2238;
assign a2246 = ~a2238 & ~a2196;
assign a2248 = a2220 & a2204;
assign a2250 = ~a2248 & a2240;
assign a2252 = ~a2250 & a2246;
assign a2256 = l338 & l96;
assign a2258 = l340 & l202;
assign a2260 = ~a2258 & ~a2256;
assign a2262 = l342 & l196;
assign a2264 = l344 & l168;
assign a2266 = ~a2264 & ~a2262;
assign a2268 = a2266 & a2260;
assign a2270 = l346 & l204;
assign a2272 = l348 & l194;
assign a2274 = ~a2272 & ~a2270;
assign a2276 = l350 & l200;
assign a2278 = l352 & l198;
assign a2280 = ~a2278 & ~a2276;
assign a2282 = a2280 & a2274;
assign a2284 = a2282 & a2268;
assign a2286 = l354 & l198;
assign a2288 = l356 & l194;
assign a2290 = ~a2288 & ~a2286;
assign a2292 = l358 & l96;
assign a2294 = l360 & l202;
assign a2296 = ~a2294 & ~a2292;
assign a2298 = a2296 & a2290;
assign a2300 = l362 & l196;
assign a2302 = l364 & l200;
assign a2304 = ~a2302 & ~a2300;
assign a2306 = l366 & l168;
assign a2308 = l368 & l204;
assign a2310 = ~a2308 & ~a2306;
assign a2312 = a2310 & a2304;
assign a2314 = a2312 & a2298;
assign a2316 = ~a2314 & a2284;
assign a2318 = l322 & l196;
assign a2320 = l324 & l96;
assign a2322 = ~a2320 & ~a2318;
assign a2324 = l326 & l168;
assign a2326 = l328 & l202;
assign a2328 = ~a2326 & ~a2324;
assign a2330 = a2328 & a2322;
assign a2332 = l330 & l198;
assign a2334 = l332 & l194;
assign a2336 = ~a2334 & ~a2332;
assign a2338 = l334 & l200;
assign a2340 = l336 & l204;
assign a2342 = ~a2340 & ~a2338;
assign a2344 = a2342 & a2336;
assign a2346 = a2344 & a2330;
assign a2348 = a2346 & l320;
assign a2350 = a2348 & a2316;
assign a2352 = a612 & ~l320;
assign a2354 = a2352 & l382;
assign a2356 = ~a2354 & ~a2350;
assign a2358 = a2314 & a2284;
assign a2360 = a2358 & a2348;
assign a2362 = a2352 & l380;
assign a2364 = ~a2362 & ~a2360;
assign a2366 = a2364 & a2356;
assign a2368 = ~a2346 & l320;
assign a2370 = a2368 & a2358;
assign a2372 = a2352 & l378;
assign a2374 = ~a2372 & ~a2370;
assign a2376 = a2348 & ~a2284;
assign a2378 = a2376 & a2314;
assign a2380 = a2352 & l376;
assign a2382 = ~a2380 & ~a2378;
assign a2384 = a2382 & a2374;
assign a2386 = a2384 & a2366;
assign a2388 = a2314 & ~a2284;
assign a2390 = a2388 & a2368;
assign a2392 = a2352 & l374;
assign a2394 = ~a2392 & ~a2390;
assign a2396 = a2394 & l320;
assign a2398 = a2376 & ~a2314;
assign a2400 = a2352 & l372;
assign a2402 = ~a2400 & ~a2398;
assign a2404 = a2368 & a2316;
assign a2406 = a2352 & l370;
assign a2408 = ~a2406 & ~a2404;
assign a2410 = a2408 & a2402;
assign a2412 = a2410 & a2396;
assign a2414 = a2412 & a2386;
assign a2416 = ~a2414 & ~l400;
assign a2418 = ~a1086 & l108;
assign a2420 = ~a1104 & ~l110;
assign a2422 = a2420 & ~a2418;
assign a2424 = a1098 & l400;
assign a2426 = ~a2424 & ~a1100;
assign a2428 = a2426 & a2422;
assign a2430 = a2428 & l316;
assign a2432 = ~a2430 & a2416;
assign a2434 = l384 & l370;
assign a2436 = l386 & l382;
assign a2438 = ~a2436 & ~a2434;
assign a2440 = l388 & l380;
assign a2442 = l390 & l372;
assign a2444 = ~a2442 & ~a2440;
assign a2446 = a2444 & a2438;
assign a2448 = ~l380 & ~l374;
assign a2450 = a2448 & ~l376;
assign a2452 = ~l382 & ~l370;
assign a2454 = ~l378 & ~l372;
assign a2456 = a2454 & a2452;
assign a2458 = a2456 & a2450;
assign a2460 = l392 & l378;
assign a2462 = l394 & l376;
assign a2464 = ~a2462 & ~a2460;
assign a2466 = l396 & l374;
assign a2468 = ~a2466 & a2464;
assign a2470 = a2468 & ~a2458;
assign a2472 = a2470 & a2446;
assign a2474 = ~l398 & ~l316;
assign a2476 = a2474 & a1094;
assign a2478 = a2476 & ~a2472;
assign a2480 = ~a2478 & l318;
assign a2482 = ~a2480 & ~l320;
assign a2486 = a2002 & l322;
assign a2488 = a1948 & l476;
assign a2490 = ~a2488 & ~a2486;
assign a2492 = a1170 & l324;
assign a2494 = a1024 & l474;
assign a2496 = ~a2494 & ~a2492;
assign a2498 = a1352 & l326;
assign a2500 = a1204 & l472;
assign a2502 = ~a2500 & ~a2498;
assign a2504 = a1940 & l328;
assign a2506 = a1886 & l470;
assign a2508 = ~a2506 & ~a2504;
assign a2510 = a2188 & l330;
assign a2512 = a2134 & l468;
assign a2514 = ~a2512 & ~a2510;
assign a2516 = a2250 & l332;
assign a2518 = a2196 & l466;
assign a2520 = ~a2518 & ~a2516;
assign a2522 = a2126 & l334;
assign a2524 = a2072 & l464;
assign a2526 = ~a2524 & ~a2522;
assign a2528 = a2064 & l336;
assign a2530 = a2010 & l462;
assign a2532 = ~a2530 & ~a2528;
assign a2534 = a1170 & l338;
assign a2536 = a1024 & l460;
assign a2538 = ~a2536 & ~a2534;
assign a2540 = a1940 & l340;
assign a2542 = a1886 & l458;
assign a2544 = ~a2542 & ~a2540;
assign a2546 = a2002 & l342;
assign a2548 = a1948 & l456;
assign a2550 = ~a2548 & ~a2546;
assign a2552 = a1352 & l344;
assign a2554 = a1204 & l454;
assign a2556 = ~a2554 & ~a2552;
assign a2558 = a2064 & l346;
assign a2560 = a2010 & l452;
assign a2562 = ~a2560 & ~a2558;
assign a2564 = a2250 & l348;
assign a2566 = a2196 & l450;
assign a2568 = ~a2566 & ~a2564;
assign a2570 = a2126 & l350;
assign a2572 = a2072 & l448;
assign a2574 = ~a2572 & ~a2570;
assign a2576 = a2188 & l352;
assign a2578 = a2134 & l446;
assign a2580 = ~a2578 & ~a2576;
assign a2582 = a2188 & l354;
assign a2584 = a2134 & l444;
assign a2586 = ~a2584 & ~a2582;
assign a2588 = a2250 & l356;
assign a2590 = a2196 & l442;
assign a2592 = ~a2590 & ~a2588;
assign a2594 = a1170 & l358;
assign a2596 = a1024 & l440;
assign a2598 = ~a2596 & ~a2594;
assign a2600 = a1940 & l360;
assign a2602 = a1886 & l438;
assign a2604 = ~a2602 & ~a2600;
assign a2606 = a2002 & l362;
assign a2608 = a1948 & l436;
assign a2610 = ~a2608 & ~a2606;
assign a2612 = a2126 & l364;
assign a2614 = a2072 & l434;
assign a2616 = ~a2614 & ~a2612;
assign a2618 = a1352 & l366;
assign a2620 = a1204 & l432;
assign a2622 = ~a2620 & ~a2618;
assign a2624 = a2064 & l368;
assign a2626 = a2010 & l430;
assign a2628 = ~a2626 & ~a2624;
assign a2630 = a1012 & ~l426;
assign a2632 = a1090 & ~l400;
assign a2634 = a2632 & a2474;
assign a2636 = ~a2634 & l370;
assign a2638 = a2630 & ~l428;
assign a2642 = ~a2640 & l384;
assign a2644 = ~a2642 & a2630;
assign a2646 = a1012 & ~l422;
assign a2648 = ~a2634 & l382;
assign a2650 = a2646 & ~l424;
assign a2654 = ~a2652 & l386;
assign a2656 = ~a2654 & a2646;
assign a2658 = a1012 & ~l418;
assign a2660 = ~a2634 & l380;
assign a2662 = a2658 & ~l420;
assign a2666 = ~a2664 & l388;
assign a2668 = ~a2666 & a2658;
assign a2670 = a1012 & ~l414;
assign a2672 = ~a2634 & l372;
assign a2674 = a2670 & ~l416;
assign a2678 = ~a2676 & l390;
assign a2680 = ~a2678 & a2670;
assign a2682 = a1012 & ~l410;
assign a2684 = ~a2634 & l378;
assign a2686 = a2682 & ~l412;
assign a2690 = ~a2688 & l392;
assign a2692 = ~a2690 & a2682;
assign a2694 = a1012 & ~l406;
assign a2696 = ~a2634 & l376;
assign a2698 = a2694 & ~l408;
assign a2702 = ~a2700 & l394;
assign a2704 = ~a2702 & a2694;
assign a2706 = a1012 & ~l402;
assign a2708 = ~a2634 & l374;
assign a2710 = a2706 & ~l404;
assign a2714 = ~a2712 & l396;
assign a2716 = ~a2714 & a2706;
assign a2718 = ~l400 & l398;
assign a2720 = a2718 & ~a2472;
assign a2722 = a2720 & a2428;
assign a2724 = a2478 & l318;
assign a2726 = ~a2724 & ~a2722;
assign a2730 = a2708 & l404;
assign a2732 = ~a2730 & ~l402;
assign a2734 = a2696 & l408;
assign a2736 = ~a2734 & ~l406;
assign a2738 = a2684 & l412;
assign a2740 = ~a2738 & ~l410;
assign a2742 = a2672 & l416;
assign a2744 = ~a2742 & ~l414;
assign a2746 = a2660 & l420;
assign a2748 = ~a2746 & ~l418;
assign a2750 = a2648 & l424;
assign a2752 = ~a2750 & ~l422;
assign a2754 = a2636 & l428;
assign a2756 = ~a2754 & ~l426;
assign a2758 = a2050 & i24;
assign a2760 = ~a2050 & l430;
assign a2762 = ~a2760 & ~a2758;
assign a2764 = a1338 & i26;
assign a2766 = ~a1338 & l432;
assign a2768 = ~a2766 & ~a2764;
assign a2770 = a2112 & i28;
assign a2772 = ~a2112 & l434;
assign a2774 = ~a2772 & ~a2770;
assign a2776 = a1988 & i30;
assign a2778 = ~a1988 & l436;
assign a2780 = ~a2778 & ~a2776;
assign a2782 = a1926 & i32;
assign a2784 = ~a1926 & l438;
assign a2786 = ~a2784 & ~a2782;
assign a2788 = a1156 & i34;
assign a2790 = ~a1156 & l440;
assign a2792 = ~a2790 & ~a2788;
assign a2794 = a2236 & i36;
assign a2796 = ~a2236 & l442;
assign a2798 = ~a2796 & ~a2794;
assign a2800 = a2174 & i38;
assign a2802 = ~a2174 & l444;
assign a2804 = ~a2802 & ~a2800;
assign a2806 = i40 & i38;
assign a2808 = ~a2806 & i42;
assign a2810 = a2808 & a2174;
assign a2812 = ~a2174 & l446;
assign a2814 = ~a2812 & ~a2810;
assign a2816 = i44 & i28;
assign a2818 = ~a2816 & i46;
assign a2820 = a2818 & a2112;
assign a2822 = ~a2112 & l448;
assign a2824 = ~a2822 & ~a2820;
assign a2826 = i48 & i36;
assign a2828 = ~a2826 & i50;
assign a2830 = a2828 & a2236;
assign a2832 = ~a2236 & l450;
assign a2834 = ~a2832 & ~a2830;
assign a2836 = i52 & i24;
assign a2838 = ~a2836 & i54;
assign a2840 = a2838 & a2050;
assign a2842 = ~a2050 & l452;
assign a2844 = ~a2842 & ~a2840;
assign a2846 = i56 & i26;
assign a2848 = ~a2846 & i58;
assign a2850 = a2848 & a1338;
assign a2852 = ~a1338 & l454;
assign a2854 = ~a2852 & ~a2850;
assign a2856 = i60 & i30;
assign a2858 = ~a2856 & i62;
assign a2860 = a2858 & a1988;
assign a2862 = ~a1988 & l456;
assign a2864 = ~a2862 & ~a2860;
assign a2866 = i64 & i32;
assign a2868 = ~a2866 & i66;
assign a2870 = a2868 & a1926;
assign a2872 = ~a1926 & l458;
assign a2874 = ~a2872 & ~a2870;
assign a2876 = i68 & i34;
assign a2878 = ~a2876 & i70;
assign a2880 = a2878 & a1156;
assign a2882 = ~a1156 & l460;
assign a2884 = ~a2882 & ~a2880;
assign a2886 = a2050 & i52;
assign a2888 = ~a2050 & l462;
assign a2890 = ~a2888 & ~a2886;
assign a2892 = a2112 & i44;
assign a2894 = ~a2112 & l464;
assign a2896 = ~a2894 & ~a2892;
assign a2898 = a2236 & i48;
assign a2900 = ~a2236 & l466;
assign a2902 = ~a2900 & ~a2898;
assign a2904 = a2174 & i40;
assign a2906 = ~a2174 & l468;
assign a2908 = ~a2906 & ~a2904;
assign a2910 = a1926 & i64;
assign a2912 = ~a1926 & l470;
assign a2914 = ~a2912 & ~a2910;
assign a2916 = a1338 & i56;
assign a2918 = ~a1338 & l472;
assign a2920 = ~a2918 & ~a2916;
assign a2922 = a1156 & i68;
assign a2924 = ~a1156 & l474;
assign a2926 = ~a2924 & ~a2922;
assign a2928 = a1988 & i60;
assign a2930 = ~a1988 & l476;
assign a2932 = ~a2930 & ~a2928;
assign a2934 = ~l484 & ~l482;
assign a2938 = l484 & l482;
assign a2940 = ~a2938 & ~l480;
assign a2942 = ~a2938 & ~a2934;
assign a2944 = ~a2942 & ~a550;
assign a2946 = ~a550 & l484;
assign p0 = l72;

assert property (~p0);

endmodule
