module m139444p (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474,i476,i478,i480,
i482,i484,i486,i488,i490,i492,i494,i496,i498,i500,i502,i504,i506,i508,i510,
i512,i514,i516,i518,i520,i522,i524,i526,i528,i530,i532,i534,i536,i538,i540,
i542,i544,i546,i548,i550,i552,i554,i556,i558,i560,i562,i564,i566,i568,i570,
i572,i574,i576,i578,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474,i476,i478,i480,
i482,i484,i486,i488,i490,i492,i494,i496,i498,i500,i502,i504,i506,i508,i510,
i512,i514,i516,i518,i520,i522,i524,i526,i528,i530,i532,i534,i536,i538,i540,
i542,i544,i546,i548,i550,i552,i554,i556,i558,i560,i562,i564,i566,i568,i570,
i572,i574,i576,i578;

output p0;

wire a1386,a1402,a1430,a1474,a1490,a1510,a1554,a1570,a1590,a1634,a1650,a1670,a1778,a1802,a1830,
a1842,a1996,a2006,a2016,a2026,a2084,a2100,a2128,a2172,a2188,a2208,a2252,a2268,a2288,a2332,
a2348,a2368,a2476,a2500,a2528,a2540,a2694,a2704,a2714,a2724,a2782,a2798,a2826,a2870,a2886,
a2906,a2950,a2966,a2986,a3030,a3046,a3066,a3174,a3198,a3226,a3238,a3392,a3402,a3412,a3422,
a3480,a3496,a3524,a3568,a3584,a3604,a3648,a3664,a3684,a3728,a3744,a3764,a3872,a3896,a3924,
a3936,a4090,a4100,a4110,a4120,a4126,a4134,a4144,a4152,a4154,a16876,c1,a1330,a1332,a1334,
a1336,a1338,a1340,a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,
a1366,a1368,a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1388,a1390,a1392,a1394,a1396,
a1398,a1400,a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1426,a1428,
a1432,a1434,a1436,a1438,a1440,a1442,a1444,a1446,a1448,a1450,a1452,a1454,a1456,a1458,a1460,
a1462,a1464,a1466,a1468,a1470,a1472,a1476,a1478,a1480,a1482,a1484,a1486,a1488,a1492,a1494,
a1496,a1498,a1500,a1502,a1504,a1506,a1508,a1512,a1514,a1516,a1518,a1520,a1522,a1524,a1526,
a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,a1548,a1550,a1552,a1556,a1558,
a1560,a1562,a1564,a1566,a1568,a1572,a1574,a1576,a1578,a1580,a1582,a1584,a1586,a1588,a1592,
a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,a1610,a1612,a1614,a1616,a1618,a1620,a1622,
a1624,a1626,a1628,a1630,a1632,a1636,a1638,a1640,a1642,a1644,a1646,a1648,a1652,a1654,a1656,
a1658,a1660,a1662,a1664,a1666,a1668,a1672,a1674,a1676,a1678,a1680,a1682,a1684,a1686,a1688,
a1690,a1692,a1694,a1696,a1698,a1700,a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,
a1720,a1722,a1724,a1726,a1728,a1730,a1732,a1734,a1736,a1738,a1740,a1742,a1744,a1746,a1748,
a1750,a1752,a1754,a1756,a1758,a1760,a1762,a1764,a1766,a1768,a1770,a1772,a1774,a1776,a1780,
a1782,a1784,a1786,a1788,a1790,a1792,a1794,a1796,a1798,a1800,a1804,a1806,a1808,a1810,a1812,
a1814,a1816,a1818,a1820,a1822,a1824,a1826,a1828,a1832,a1834,a1836,a1838,a1840,a1844,a1846,
a1848,a1850,a1852,a1854,a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,
a1878,a1880,a1882,a1884,a1886,a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,
a1908,a1910,a1912,a1914,a1916,a1918,a1920,a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,
a1938,a1940,a1942,a1944,a1946,a1948,a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,
a1968,a1970,a1972,a1974,a1976,a1978,a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1998,
a2000,a2002,a2004,a2008,a2010,a2012,a2014,a2018,a2020,a2022,a2024,a2028,a2030,a2032,a2034,
a2036,a2038,a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,a2058,a2060,a2062,a2064,
a2066,a2068,a2070,a2072,a2074,a2076,a2078,a2080,a2082,a2086,a2088,a2090,a2092,a2094,a2096,
a2098,a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,a2120,a2122,a2124,a2126,a2130,
a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,a2152,a2154,a2156,a2158,a2160,
a2162,a2164,a2166,a2168,a2170,a2174,a2176,a2178,a2180,a2182,a2184,a2186,a2190,a2192,a2194,
a2196,a2198,a2200,a2202,a2204,a2206,a2210,a2212,a2214,a2216,a2218,a2220,a2222,a2224,a2226,
a2228,a2230,a2232,a2234,a2236,a2238,a2240,a2242,a2244,a2246,a2248,a2250,a2254,a2256,a2258,
a2260,a2262,a2264,a2266,a2270,a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2290,a2292,
a2294,a2296,a2298,a2300,a2302,a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,
a2324,a2326,a2328,a2330,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2350,a2352,a2354,a2356,
a2358,a2360,a2362,a2364,a2366,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,a2388,
a2390,a2392,a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,
a2420,a2422,a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,a2448,
a2450,a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2478,a2480,
a2482,a2484,a2486,a2488,a2490,a2492,a2494,a2496,a2498,a2502,a2504,a2506,a2508,a2510,a2512,
a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2530,a2532,a2534,a2536,a2538,a2542,a2544,a2546,
a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,a2572,a2574,a2576,
a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,a2602,a2604,a2606,
a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,a2630,a2632,a2634,a2636,
a2638,a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,a2662,a2664,a2666,
a2668,a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,a2692,a2696,a2698,
a2700,a2702,a2706,a2708,a2710,a2712,a2716,a2718,a2720,a2722,a2726,a2728,a2730,a2732,a2734,
a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,a2752,a2754,a2756,a2758,a2760,a2762,a2764,
a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,a2784,a2786,a2788,a2790,a2792,a2794,a2796,
a2800,a2802,a2804,a2806,a2808,a2810,a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2828,a2830,
a2832,a2834,a2836,a2838,a2840,a2842,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,
a2862,a2864,a2866,a2868,a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2888,a2890,a2892,a2894,
a2896,a2898,a2900,a2902,a2904,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,
a2928,a2930,a2932,a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2952,a2954,a2956,a2958,
a2960,a2962,a2964,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2988,a2990,a2992,
a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,a3022,
a3024,a3026,a3028,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3048,a3050,a3052,a3054,a3056,
a3058,a3060,a3062,a3064,a3068,a3070,a3072,a3074,a3076,a3078,a3080,a3082,a3084,a3086,a3088,
a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,a3112,a3114,a3116,a3118,
a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,a3142,a3144,a3146,a3148,
a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,a3172,a3176,a3178,a3180,
a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3200,a3202,a3204,a3206,a3208,a3210,a3212,
a3214,a3216,a3218,a3220,a3222,a3224,a3228,a3230,a3232,a3234,a3236,a3240,a3242,a3244,a3246,
a3248,a3250,a3252,a3254,a3256,a3258,a3260,a3262,a3264,a3266,a3268,a3270,a3272,a3274,a3276,
a3278,a3280,a3282,a3284,a3286,a3288,a3290,a3292,a3294,a3296,a3298,a3300,a3302,a3304,a3306,
a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,a3324,a3326,a3328,a3330,a3332,a3334,a3336,
a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,a3354,a3356,a3358,a3360,a3362,a3364,a3366,
a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3382,a3384,a3386,a3388,a3390,a3394,a3396,a3398,
a3400,a3404,a3406,a3408,a3410,a3414,a3416,a3418,a3420,a3424,a3426,a3428,a3430,a3432,a3434,
a3436,a3438,a3440,a3442,a3444,a3446,a3448,a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,
a3466,a3468,a3470,a3472,a3474,a3476,a3478,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3498,
a3500,a3502,a3504,a3506,a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3526,a3528,a3530,
a3532,a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,a3558,a3560,
a3562,a3564,a3566,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3586,a3588,a3590,a3592,a3594,
a3596,a3598,a3600,a3602,a3606,a3608,a3610,a3612,a3614,a3616,a3618,a3620,a3622,a3624,a3626,
a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3650,a3652,a3654,a3656,a3658,
a3660,a3662,a3666,a3668,a3670,a3672,a3674,a3676,a3678,a3680,a3682,a3686,a3688,a3690,a3692,
a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,a3712,a3714,a3716,a3718,a3720,a3722,
a3724,a3726,a3730,a3732,a3734,a3736,a3738,a3740,a3742,a3746,a3748,a3750,a3752,a3754,a3756,
a3758,a3760,a3762,a3766,a3768,a3770,a3772,a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,
a3790,a3792,a3794,a3796,a3798,a3800,a3802,a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,
a3820,a3822,a3824,a3826,a3828,a3830,a3832,a3834,a3836,a3838,a3840,a3842,a3844,a3846,a3848,
a3850,a3852,a3854,a3856,a3858,a3860,a3862,a3864,a3866,a3868,a3870,a3874,a3876,a3878,a3880,
a3882,a3884,a3886,a3888,a3890,a3892,a3894,a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,
a3914,a3916,a3918,a3920,a3922,a3926,a3928,a3930,a3932,a3934,a3938,a3940,a3942,a3944,a3946,
a3948,a3950,a3952,a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,
a3978,a3980,a3982,a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,
a4008,a4010,a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,
a4038,a4040,a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,
a4068,a4070,a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4092,a4094,a4096,a4098,
a4102,a4104,a4106,a4108,a4112,a4114,a4116,a4118,a4122,a4124,a4128,a4130,a4132,a4136,a4138,
a4140,a4142,a4146,a4148,a4150,a4156,a4158,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,
a4176,a4178,a4180,a4182,a4184,a4186,a4188,a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,
a4206,a4208,a4210,a4212,a4214,a4216,a4218,a4220,a4222,a4224,a4226,a4228,a4230,a4232,a4234,
a4236,a4238,a4240,a4242,a4244,a4246,a4248,a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,
a4266,a4268,a4270,a4272,a4274,a4276,a4278,a4280,a4282,a4284,a4286,a4288,a4290,a4292,a4294,
a4296,a4298,a4300,a4302,a4304,a4306,a4308,a4310,a4312,a4314,a4316,a4318,a4320,a4322,a4324,
a4326,a4328,a4330,a4332,a4334,a4336,a4338,a4340,a4342,a4344,a4346,a4348,a4350,a4352,a4354,
a4356,a4358,a4360,a4362,a4364,a4366,a4368,a4370,a4372,a4374,a4376,a4378,a4380,a4382,a4384,
a4386,a4388,a4390,a4392,a4394,a4396,a4398,a4400,a4402,a4404,a4406,a4408,a4410,a4412,a4414,
a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,a4432,a4434,a4436,a4438,a4440,a4442,a4444,
a4446,a4448,a4450,a4452,a4454,a4456,a4458,a4460,a4462,a4464,a4466,a4468,a4470,a4472,a4474,
a4476,a4478,a4480,a4482,a4484,a4486,a4488,a4490,a4492,a4494,a4496,a4498,a4500,a4502,a4504,
a4506,a4508,a4510,a4512,a4514,a4516,a4518,a4520,a4522,a4524,a4526,a4528,a4530,a4532,a4534,
a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,a4554,a4556,a4558,a4560,a4562,a4564,
a4566,a4568,a4570,a4572,a4574,a4576,a4578,a4580,a4582,a4584,a4586,a4588,a4590,a4592,a4594,
a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,a4612,a4614,a4616,a4618,a4620,a4622,a4624,
a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,a4642,a4644,a4646,a4648,a4650,a4652,a4654,
a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,a4672,a4674,a4676,a4678,a4680,a4682,a4684,
a4686,a4688,a4690,a4692,a4694,a4696,a4698,a4700,a4702,a4704,a4706,a4708,a4710,a4712,a4714,
a4716,a4718,a4720,a4722,a4724,a4726,a4728,a4730,a4732,a4734,a4736,a4738,a4740,a4742,a4744,
a4746,a4748,a4750,a4752,a4754,a4756,a4758,a4760,a4762,a4764,a4766,a4768,a4770,a4772,a4774,
a4776,a4778,a4780,a4782,a4784,a4786,a4788,a4790,a4792,a4794,a4796,a4798,a4800,a4802,a4804,
a4806,a4808,a4810,a4812,a4814,a4816,a4818,a4820,a4822,a4824,a4826,a4828,a4830,a4832,a4834,
a4836,a4838,a4840,a4842,a4844,a4846,a4848,a4850,a4852,a4854,a4856,a4858,a4860,a4862,a4864,
a4866,a4868,a4870,a4872,a4874,a4876,a4878,a4880,a4882,a4884,a4886,a4888,a4890,a4892,a4894,
a4896,a4898,a4900,a4902,a4904,a4906,a4908,a4910,a4912,a4914,a4916,a4918,a4920,a4922,a4924,
a4926,a4928,a4930,a4932,a4934,a4936,a4938,a4940,a4942,a4944,a4946,a4948,a4950,a4952,a4954,
a4956,a4958,a4960,a4962,a4964,a4966,a4968,a4970,a4972,a4974,a4976,a4978,a4980,a4982,a4984,
a4986,a4988,a4990,a4992,a4994,a4996,a4998,a5000,a5002,a5004,a5006,a5008,a5010,a5012,a5014,
a5016,a5018,a5020,a5022,a5024,a5026,a5028,a5030,a5032,a5034,a5036,a5038,a5040,a5042,a5044,
a5046,a5048,a5050,a5052,a5054,a5056,a5058,a5060,a5062,a5064,a5066,a5068,a5070,a5072,a5074,
a5076,a5078,a5080,a5082,a5084,a5086,a5088,a5090,a5092,a5094,a5096,a5098,a5100,a5102,a5104,
a5106,a5108,a5110,a5112,a5114,a5116,a5118,a5120,a5122,a5124,a5126,a5128,a5130,a5132,a5134,
a5136,a5138,a5140,a5142,a5144,a5146,a5148,a5150,a5152,a5154,a5156,a5158,a5160,a5162,a5164,
a5166,a5168,a5170,a5172,a5174,a5176,a5178,a5180,a5182,a5184,a5186,a5188,a5190,a5192,a5194,
a5196,a5198,a5200,a5202,a5204,a5206,a5208,a5210,a5212,a5214,a5216,a5218,a5220,a5222,a5224,
a5226,a5228,a5230,a5232,a5234,a5236,a5238,a5240,a5242,a5244,a5246,a5248,a5250,a5252,a5254,
a5256,a5258,a5260,a5262,a5264,a5266,a5268,a5270,a5272,a5274,a5276,a5278,a5280,a5282,a5284,
a5286,a5288,a5290,a5292,a5294,a5296,a5298,a5300,a5302,a5304,a5306,a5308,a5310,a5312,a5314,
a5316,a5318,a5320,a5322,a5324,a5326,a5328,a5330,a5332,a5334,a5336,a5338,a5340,a5342,a5344,
a5346,a5348,a5350,a5352,a5354,a5356,a5358,a5360,a5362,a5364,a5366,a5368,a5370,a5372,a5374,
a5376,a5378,a5380,a5382,a5384,a5386,a5388,a5390,a5392,a5394,a5396,a5398,a5400,a5402,a5404,
a5406,a5408,a5410,a5412,a5414,a5416,a5418,a5420,a5422,a5424,a5426,a5428,a5430,a5432,a5434,
a5436,a5438,a5440,a5442,a5444,a5446,a5448,a5450,a5452,a5454,a5456,a5458,a5460,a5462,a5464,
a5466,a5468,a5470,a5472,a5474,a5476,a5478,a5480,a5482,a5484,a5486,a5488,a5490,a5492,a5494,
a5496,a5498,a5500,a5502,a5504,a5506,a5508,a5510,a5512,a5514,a5516,a5518,a5520,a5522,a5524,
a5526,a5528,a5530,a5532,a5534,a5536,a5538,a5540,a5542,a5544,a5546,a5548,a5550,a5552,a5554,
a5556,a5558,a5560,a5562,a5564,a5566,a5568,a5570,a5572,a5574,a5576,a5578,a5580,a5582,a5584,
a5586,a5588,a5590,a5592,a5594,a5596,a5598,a5600,a5602,a5604,a5606,a5608,a5610,a5612,a5614,
a5616,a5618,a5620,a5622,a5624,a5626,a5628,a5630,a5632,a5634,a5636,a5638,a5640,a5642,a5644,
a5646,a5648,a5650,a5652,a5654,a5656,a5658,a5660,a5662,a5664,a5666,a5668,a5670,a5672,a5674,
a5676,a5678,a5680,a5682,a5684,a5686,a5688,a5690,a5692,a5694,a5696,a5698,a5700,a5702,a5704,
a5706,a5708,a5710,a5712,a5714,a5716,a5718,a5720,a5722,a5724,a5726,a5728,a5730,a5732,a5734,
a5736,a5738,a5740,a5742,a5744,a5746,a5748,a5750,a5752,a5754,a5756,a5758,a5760,a5762,a5764,
a5766,a5768,a5770,a5772,a5774,a5776,a5778,a5780,a5782,a5784,a5786,a5788,a5790,a5792,a5794,
a5796,a5798,a5800,a5802,a5804,a5806,a5808,a5810,a5812,a5814,a5816,a5818,a5820,a5822,a5824,
a5826,a5828,a5830,a5832,a5834,a5836,a5838,a5840,a5842,a5844,a5846,a5848,a5850,a5852,a5854,
a5856,a5858,a5860,a5862,a5864,a5866,a5868,a5870,a5872,a5874,a5876,a5878,a5880,a5882,a5884,
a5886,a5888,a5890,a5892,a5894,a5896,a5898,a5900,a5902,a5904,a5906,a5908,a5910,a5912,a5914,
a5916,a5918,a5920,a5922,a5924,a5926,a5928,a5930,a5932,a5934,a5936,a5938,a5940,a5942,a5944,
a5946,a5948,a5950,a5952,a5954,a5956,a5958,a5960,a5962,a5964,a5966,a5968,a5970,a5972,a5974,
a5976,a5978,a5980,a5982,a5984,a5986,a5988,a5990,a5992,a5994,a5996,a5998,a6000,a6002,a6004,
a6006,a6008,a6010,a6012,a6014,a6016,a6018,a6020,a6022,a6024,a6026,a6028,a6030,a6032,a6034,
a6036,a6038,a6040,a6042,a6044,a6046,a6048,a6050,a6052,a6054,a6056,a6058,a6060,a6062,a6064,
a6066,a6068,a6070,a6072,a6074,a6076,a6078,a6080,a6082,a6084,a6086,a6088,a6090,a6092,a6094,
a6096,a6098,a6100,a6102,a6104,a6106,a6108,a6110,a6112,a6114,a6116,a6118,a6120,a6122,a6124,
a6126,a6128,a6130,a6132,a6134,a6136,a6138,a6140,a6142,a6144,a6146,a6148,a6150,a6152,a6154,
a6156,a6158,a6160,a6162,a6164,a6166,a6168,a6170,a6172,a6174,a6176,a6178,a6180,a6182,a6184,
a6186,a6188,a6190,a6192,a6194,a6196,a6198,a6200,a6202,a6204,a6206,a6208,a6210,a6212,a6214,
a6216,a6218,a6220,a6222,a6224,a6226,a6228,a6230,a6232,a6234,a6236,a6238,a6240,a6242,a6244,
a6246,a6248,a6250,a6252,a6254,a6256,a6258,a6260,a6262,a6264,a6266,a6268,a6270,a6272,a6274,
a6276,a6278,a6280,a6282,a6284,a6286,a6288,a6290,a6292,a6294,a6296,a6298,a6300,a6302,a6304,
a6306,a6308,a6310,a6312,a6314,a6316,a6318,a6320,a6322,a6324,a6326,a6328,a6330,a6332,a6334,
a6336,a6338,a6340,a6342,a6344,a6346,a6348,a6350,a6352,a6354,a6356,a6358,a6360,a6362,a6364,
a6366,a6368,a6370,a6372,a6374,a6376,a6378,a6380,a6382,a6384,a6386,a6388,a6390,a6392,a6394,
a6396,a6398,a6400,a6402,a6404,a6406,a6408,a6410,a6412,a6414,a6416,a6418,a6420,a6422,a6424,
a6426,a6428,a6430,a6432,a6434,a6436,a6438,a6440,a6442,a6444,a6446,a6448,a6450,a6452,a6454,
a6456,a6458,a6460,a6462,a6464,a6466,a6468,a6470,a6472,a6474,a6476,a6478,a6480,a6482,a6484,
a6486,a6488,a6490,a6492,a6494,a6496,a6498,a6500,a6502,a6504,a6506,a6508,a6510,a6512,a6514,
a6516,a6518,a6520,a6522,a6524,a6526,a6528,a6530,a6532,a6534,a6536,a6538,a6540,a6542,a6544,
a6546,a6548,a6550,a6552,a6554,a6556,a6558,a6560,a6562,a6564,a6566,a6568,a6570,a6572,a6574,
a6576,a6578,a6580,a6582,a6584,a6586,a6588,a6590,a6592,a6594,a6596,a6598,a6600,a6602,a6604,
a6606,a6608,a6610,a6612,a6614,a6616,a6618,a6620,a6622,a6624,a6626,a6628,a6630,a6632,a6634,
a6636,a6638,a6640,a6642,a6644,a6646,a6648,a6650,a6652,a6654,a6656,a6658,a6660,a6662,a6664,
a6666,a6668,a6670,a6672,a6674,a6676,a6678,a6680,a6682,a6684,a6686,a6688,a6690,a6692,a6694,
a6696,a6698,a6700,a6702,a6704,a6706,a6708,a6710,a6712,a6714,a6716,a6718,a6720,a6722,a6724,
a6726,a6728,a6730,a6732,a6734,a6736,a6738,a6740,a6742,a6744,a6746,a6748,a6750,a6752,a6754,
a6756,a6758,a6760,a6762,a6764,a6766,a6768,a6770,a6772,a6774,a6776,a6778,a6780,a6782,a6784,
a6786,a6788,a6790,a6792,a6794,a6796,a6798,a6800,a6802,a6804,a6806,a6808,a6810,a6812,a6814,
a6816,a6818,a6820,a6822,a6824,a6826,a6828,a6830,a6832,a6834,a6836,a6838,a6840,a6842,a6844,
a6846,a6848,a6850,a6852,a6854,a6856,a6858,a6860,a6862,a6864,a6866,a6868,a6870,a6872,a6874,
a6876,a6878,a6880,a6882,a6884,a6886,a6888,a6890,a6892,a6894,a6896,a6898,a6900,a6902,a6904,
a6906,a6908,a6910,a6912,a6914,a6916,a6918,a6920,a6922,a6924,a6926,a6928,a6930,a6932,a6934,
a6936,a6938,a6940,a6942,a6944,a6946,a6948,a6950,a6952,a6954,a6956,a6958,a6960,a6962,a6964,
a6966,a6968,a6970,a6972,a6974,a6976,a6978,a6980,a6982,a6984,a6986,a6988,a6990,a6992,a6994,
a6996,a6998,a7000,a7002,a7004,a7006,a7008,a7010,a7012,a7014,a7016,a7018,a7020,a7022,a7024,
a7026,a7028,a7030,a7032,a7034,a7036,a7038,a7040,a7042,a7044,a7046,a7048,a7050,a7052,a7054,
a7056,a7058,a7060,a7062,a7064,a7066,a7068,a7070,a7072,a7074,a7076,a7078,a7080,a7082,a7084,
a7086,a7088,a7090,a7092,a7094,a7096,a7098,a7100,a7102,a7104,a7106,a7108,a7110,a7112,a7114,
a7116,a7118,a7120,a7122,a7124,a7126,a7128,a7130,a7132,a7134,a7136,a7138,a7140,a7142,a7144,
a7146,a7148,a7150,a7152,a7154,a7156,a7158,a7160,a7162,a7164,a7166,a7168,a7170,a7172,a7174,
a7176,a7178,a7180,a7182,a7184,a7186,a7188,a7190,a7192,a7194,a7196,a7198,a7200,a7202,a7204,
a7206,a7208,a7210,a7212,a7214,a7216,a7218,a7220,a7222,a7224,a7226,a7228,a7230,a7232,a7234,
a7236,a7238,a7240,a7242,a7244,a7246,a7248,a7250,a7252,a7254,a7256,a7258,a7260,a7262,a7264,
a7266,a7268,a7270,a7272,a7274,a7276,a7278,a7280,a7282,a7284,a7286,a7288,a7290,a7292,a7294,
a7296,a7298,a7300,a7302,a7304,a7306,a7308,a7310,a7312,a7314,a7316,a7318,a7320,a7322,a7324,
a7326,a7328,a7330,a7332,a7334,a7336,a7338,a7340,a7342,a7344,a7346,a7348,a7350,a7352,a7354,
a7356,a7358,a7360,a7362,a7364,a7366,a7368,a7370,a7372,a7374,a7376,a7378,a7380,a7382,a7384,
a7386,a7388,a7390,a7392,a7394,a7396,a7398,a7400,a7402,a7404,a7406,a7408,a7410,a7412,a7414,
a7416,a7418,a7420,a7422,a7424,a7426,a7428,a7430,a7432,a7434,a7436,a7438,a7440,a7442,a7444,
a7446,a7448,a7450,a7452,a7454,a7456,a7458,a7460,a7462,a7464,a7466,a7468,a7470,a7472,a7474,
a7476,a7478,a7480,a7482,a7484,a7486,a7488,a7490,a7492,a7494,a7496,a7498,a7500,a7502,a7504,
a7506,a7508,a7510,a7512,a7514,a7516,a7518,a7520,a7522,a7524,a7526,a7528,a7530,a7532,a7534,
a7536,a7538,a7540,a7542,a7544,a7546,a7548,a7550,a7552,a7554,a7556,a7558,a7560,a7562,a7564,
a7566,a7568,a7570,a7572,a7574,a7576,a7578,a7580,a7582,a7584,a7586,a7588,a7590,a7592,a7594,
a7596,a7598,a7600,a7602,a7604,a7606,a7608,a7610,a7612,a7614,a7616,a7618,a7620,a7622,a7624,
a7626,a7628,a7630,a7632,a7634,a7636,a7638,a7640,a7642,a7644,a7646,a7648,a7650,a7652,a7654,
a7656,a7658,a7660,a7662,a7664,a7666,a7668,a7670,a7672,a7674,a7676,a7678,a7680,a7682,a7684,
a7686,a7688,a7690,a7692,a7694,a7696,a7698,a7700,a7702,a7704,a7706,a7708,a7710,a7712,a7714,
a7716,a7718,a7720,a7722,a7724,a7726,a7728,a7730,a7732,a7734,a7736,a7738,a7740,a7742,a7744,
a7746,a7748,a7750,a7752,a7754,a7756,a7758,a7760,a7762,a7764,a7766,a7768,a7770,a7772,a7774,
a7776,a7778,a7780,a7782,a7784,a7786,a7788,a7790,a7792,a7794,a7796,a7798,a7800,a7802,a7804,
a7806,a7808,a7810,a7812,a7814,a7816,a7818,a7820,a7822,a7824,a7826,a7828,a7830,a7832,a7834,
a7836,a7838,a7840,a7842,a7844,a7846,a7848,a7850,a7852,a7854,a7856,a7858,a7860,a7862,a7864,
a7866,a7868,a7870,a7872,a7874,a7876,a7878,a7880,a7882,a7884,a7886,a7888,a7890,a7892,a7894,
a7896,a7898,a7900,a7902,a7904,a7906,a7908,a7910,a7912,a7914,a7916,a7918,a7920,a7922,a7924,
a7926,a7928,a7930,a7932,a7934,a7936,a7938,a7940,a7942,a7944,a7946,a7948,a7950,a7952,a7954,
a7956,a7958,a7960,a7962,a7964,a7966,a7968,a7970,a7972,a7974,a7976,a7978,a7980,a7982,a7984,
a7986,a7988,a7990,a7992,a7994,a7996,a7998,a8000,a8002,a8004,a8006,a8008,a8010,a8012,a8014,
a8016,a8018,a8020,a8022,a8024,a8026,a8028,a8030,a8032,a8034,a8036,a8038,a8040,a8042,a8044,
a8046,a8048,a8050,a8052,a8054,a8056,a8058,a8060,a8062,a8064,a8066,a8068,a8070,a8072,a8074,
a8076,a8078,a8080,a8082,a8084,a8086,a8088,a8090,a8092,a8094,a8096,a8098,a8100,a8102,a8104,
a8106,a8108,a8110,a8112,a8114,a8116,a8118,a8120,a8122,a8124,a8126,a8128,a8130,a8132,a8134,
a8136,a8138,a8140,a8142,a8144,a8146,a8148,a8150,a8152,a8154,a8156,a8158,a8160,a8162,a8164,
a8166,a8168,a8170,a8172,a8174,a8176,a8178,a8180,a8182,a8184,a8186,a8188,a8190,a8192,a8194,
a8196,a8198,a8200,a8202,a8204,a8206,a8208,a8210,a8212,a8214,a8216,a8218,a8220,a8222,a8224,
a8226,a8228,a8230,a8232,a8234,a8236,a8238,a8240,a8242,a8244,a8246,a8248,a8250,a8252,a8254,
a8256,a8258,a8260,a8262,a8264,a8266,a8268,a8270,a8272,a8274,a8276,a8278,a8280,a8282,a8284,
a8286,a8288,a8290,a8292,a8294,a8296,a8298,a8300,a8302,a8304,a8306,a8308,a8310,a8312,a8314,
a8316,a8318,a8320,a8322,a8324,a8326,a8328,a8330,a8332,a8334,a8336,a8338,a8340,a8342,a8344,
a8346,a8348,a8350,a8352,a8354,a8356,a8358,a8360,a8362,a8364,a8366,a8368,a8370,a8372,a8374,
a8376,a8378,a8380,a8382,a8384,a8386,a8388,a8390,a8392,a8394,a8396,a8398,a8400,a8402,a8404,
a8406,a8408,a8410,a8412,a8414,a8416,a8418,a8420,a8422,a8424,a8426,a8428,a8430,a8432,a8434,
a8436,a8438,a8440,a8442,a8444,a8446,a8448,a8450,a8452,a8454,a8456,a8458,a8460,a8462,a8464,
a8466,a8468,a8470,a8472,a8474,a8476,a8478,a8480,a8482,a8484,a8486,a8488,a8490,a8492,a8494,
a8496,a8498,a8500,a8502,a8504,a8506,a8508,a8510,a8512,a8514,a8516,a8518,a8520,a8522,a8524,
a8526,a8528,a8530,a8532,a8534,a8536,a8538,a8540,a8542,a8544,a8546,a8548,a8550,a8552,a8554,
a8556,a8558,a8560,a8562,a8564,a8566,a8568,a8570,a8572,a8574,a8576,a8578,a8580,a8582,a8584,
a8586,a8588,a8590,a8592,a8594,a8596,a8598,a8600,a8602,a8604,a8606,a8608,a8610,a8612,a8614,
a8616,a8618,a8620,a8622,a8624,a8626,a8628,a8630,a8632,a8634,a8636,a8638,a8640,a8642,a8644,
a8646,a8648,a8650,a8652,a8654,a8656,a8658,a8660,a8662,a8664,a8666,a8668,a8670,a8672,a8674,
a8676,a8678,a8680,a8682,a8684,a8686,a8688,a8690,a8692,a8694,a8696,a8698,a8700,a8702,a8704,
a8706,a8708,a8710,a8712,a8714,a8716,a8718,a8720,a8722,a8724,a8726,a8728,a8730,a8732,a8734,
a8736,a8738,a8740,a8742,a8744,a8746,a8748,a8750,a8752,a8754,a8756,a8758,a8760,a8762,a8764,
a8766,a8768,a8770,a8772,a8774,a8776,a8778,a8780,a8782,a8784,a8786,a8788,a8790,a8792,a8794,
a8796,a8798,a8800,a8802,a8804,a8806,a8808,a8810,a8812,a8814,a8816,a8818,a8820,a8822,a8824,
a8826,a8828,a8830,a8832,a8834,a8836,a8838,a8840,a8842,a8844,a8846,a8848,a8850,a8852,a8854,
a8856,a8858,a8860,a8862,a8864,a8866,a8868,a8870,a8872,a8874,a8876,a8878,a8880,a8882,a8884,
a8886,a8888,a8890,a8892,a8894,a8896,a8898,a8900,a8902,a8904,a8906,a8908,a8910,a8912,a8914,
a8916,a8918,a8920,a8922,a8924,a8926,a8928,a8930,a8932,a8934,a8936,a8938,a8940,a8942,a8944,
a8946,a8948,a8950,a8952,a8954,a8956,a8958,a8960,a8962,a8964,a8966,a8968,a8970,a8972,a8974,
a8976,a8978,a8980,a8982,a8984,a8986,a8988,a8990,a8992,a8994,a8996,a8998,a9000,a9002,a9004,
a9006,a9008,a9010,a9012,a9014,a9016,a9018,a9020,a9022,a9024,a9026,a9028,a9030,a9032,a9034,
a9036,a9038,a9040,a9042,a9044,a9046,a9048,a9050,a9052,a9054,a9056,a9058,a9060,a9062,a9064,
a9066,a9068,a9070,a9072,a9074,a9076,a9078,a9080,a9082,a9084,a9086,a9088,a9090,a9092,a9094,
a9096,a9098,a9100,a9102,a9104,a9106,a9108,a9110,a9112,a9114,a9116,a9118,a9120,a9122,a9124,
a9126,a9128,a9130,a9132,a9134,a9136,a9138,a9140,a9142,a9144,a9146,a9148,a9150,a9152,a9154,
a9156,a9158,a9160,a9162,a9164,a9166,a9168,a9170,a9172,a9174,a9176,a9178,a9180,a9182,a9184,
a9186,a9188,a9190,a9192,a9194,a9196,a9198,a9200,a9202,a9204,a9206,a9208,a9210,a9212,a9214,
a9216,a9218,a9220,a9222,a9224,a9226,a9228,a9230,a9232,a9234,a9236,a9238,a9240,a9242,a9244,
a9246,a9248,a9250,a9252,a9254,a9256,a9258,a9260,a9262,a9264,a9266,a9268,a9270,a9272,a9274,
a9276,a9278,a9280,a9282,a9284,a9286,a9288,a9290,a9292,a9294,a9296,a9298,a9300,a9302,a9304,
a9306,a9308,a9310,a9312,a9314,a9316,a9318,a9320,a9322,a9324,a9326,a9328,a9330,a9332,a9334,
a9336,a9338,a9340,a9342,a9344,a9346,a9348,a9350,a9352,a9354,a9356,a9358,a9360,a9362,a9364,
a9366,a9368,a9370,a9372,a9374,a9376,a9378,a9380,a9382,a9384,a9386,a9388,a9390,a9392,a9394,
a9396,a9398,a9400,a9402,a9404,a9406,a9408,a9410,a9412,a9414,a9416,a9418,a9420,a9422,a9424,
a9426,a9428,a9430,a9432,a9434,a9436,a9438,a9440,a9442,a9444,a9446,a9448,a9450,a9452,a9454,
a9456,a9458,a9460,a9462,a9464,a9466,a9468,a9470,a9472,a9474,a9476,a9478,a9480,a9482,a9484,
a9486,a9488,a9490,a9492,a9494,a9496,a9498,a9500,a9502,a9504,a9506,a9508,a9510,a9512,a9514,
a9516,a9518,a9520,a9522,a9524,a9526,a9528,a9530,a9532,a9534,a9536,a9538,a9540,a9542,a9544,
a9546,a9548,a9550,a9552,a9554,a9556,a9558,a9560,a9562,a9564,a9566,a9568,a9570,a9572,a9574,
a9576,a9578,a9580,a9582,a9584,a9586,a9588,a9590,a9592,a9594,a9596,a9598,a9600,a9602,a9604,
a9606,a9608,a9610,a9612,a9614,a9616,a9618,a9620,a9622,a9624,a9626,a9628,a9630,a9632,a9634,
a9636,a9638,a9640,a9642,a9644,a9646,a9648,a9650,a9652,a9654,a9656,a9658,a9660,a9662,a9664,
a9666,a9668,a9670,a9672,a9674,a9676,a9678,a9680,a9682,a9684,a9686,a9688,a9690,a9692,a9694,
a9696,a9698,a9700,a9702,a9704,a9706,a9708,a9710,a9712,a9714,a9716,a9718,a9720,a9722,a9724,
a9726,a9728,a9730,a9732,a9734,a9736,a9738,a9740,a9742,a9744,a9746,a9748,a9750,a9752,a9754,
a9756,a9758,a9760,a9762,a9764,a9766,a9768,a9770,a9772,a9774,a9776,a9778,a9780,a9782,a9784,
a9786,a9788,a9790,a9792,a9794,a9796,a9798,a9800,a9802,a9804,a9806,a9808,a9810,a9812,a9814,
a9816,a9818,a9820,a9822,a9824,a9826,a9828,a9830,a9832,a9834,a9836,a9838,a9840,a9842,a9844,
a9846,a9848,a9850,a9852,a9854,a9856,a9858,a9860,a9862,a9864,a9866,a9868,a9870,a9872,a9874,
a9876,a9878,a9880,a9882,a9884,a9886,a9888,a9890,a9892,a9894,a9896,a9898,a9900,a9902,a9904,
a9906,a9908,a9910,a9912,a9914,a9916,a9918,a9920,a9922,a9924,a9926,a9928,a9930,a9932,a9934,
a9936,a9938,a9940,a9942,a9944,a9946,a9948,a9950,a9952,a9954,a9956,a9958,a9960,a9962,a9964,
a9966,a9968,a9970,a9972,a9974,a9976,a9978,a9980,a9982,a9984,a9986,a9988,a9990,a9992,a9994,
a9996,a9998,a10000,a10002,a10004,a10006,a10008,a10010,a10012,a10014,a10016,a10018,a10020,a10022,a10024,
a10026,a10028,a10030,a10032,a10034,a10036,a10038,a10040,a10042,a10044,a10046,a10048,a10050,a10052,a10054,
a10056,a10058,a10060,a10062,a10064,a10066,a10068,a10070,a10072,a10074,a10076,a10078,a10080,a10082,a10084,
a10086,a10088,a10090,a10092,a10094,a10096,a10098,a10100,a10102,a10104,a10106,a10108,a10110,a10112,a10114,
a10116,a10118,a10120,a10122,a10124,a10126,a10128,a10130,a10132,a10134,a10136,a10138,a10140,a10142,a10144,
a10146,a10148,a10150,a10152,a10154,a10156,a10158,a10160,a10162,a10164,a10166,a10168,a10170,a10172,a10174,
a10176,a10178,a10180,a10182,a10184,a10186,a10188,a10190,a10192,a10194,a10196,a10198,a10200,a10202,a10204,
a10206,a10208,a10210,a10212,a10214,a10216,a10218,a10220,a10222,a10224,a10226,a10228,a10230,a10232,a10234,
a10236,a10238,a10240,a10242,a10244,a10246,a10248,a10250,a10252,a10254,a10256,a10258,a10260,a10262,a10264,
a10266,a10268,a10270,a10272,a10274,a10276,a10278,a10280,a10282,a10284,a10286,a10288,a10290,a10292,a10294,
a10296,a10298,a10300,a10302,a10304,a10306,a10308,a10310,a10312,a10314,a10316,a10318,a10320,a10322,a10324,
a10326,a10328,a10330,a10332,a10334,a10336,a10338,a10340,a10342,a10344,a10346,a10348,a10350,a10352,a10354,
a10356,a10358,a10360,a10362,a10364,a10366,a10368,a10370,a10372,a10374,a10376,a10378,a10380,a10382,a10384,
a10386,a10388,a10390,a10392,a10394,a10396,a10398,a10400,a10402,a10404,a10406,a10408,a10410,a10412,a10414,
a10416,a10418,a10420,a10422,a10424,a10426,a10428,a10430,a10432,a10434,a10436,a10438,a10440,a10442,a10444,
a10446,a10448,a10450,a10452,a10454,a10456,a10458,a10460,a10462,a10464,a10466,a10468,a10470,a10472,a10474,
a10476,a10478,a10480,a10482,a10484,a10486,a10488,a10490,a10492,a10494,a10496,a10498,a10500,a10502,a10504,
a10506,a10508,a10510,a10512,a10514,a10516,a10518,a10520,a10522,a10524,a10526,a10528,a10530,a10532,a10534,
a10536,a10538,a10540,a10542,a10544,a10546,a10548,a10550,a10552,a10554,a10556,a10558,a10560,a10562,a10564,
a10566,a10568,a10570,a10572,a10574,a10576,a10578,a10580,a10582,a10584,a10586,a10588,a10590,a10592,a10594,
a10596,a10598,a10600,a10602,a10604,a10606,a10608,a10610,a10612,a10614,a10616,a10618,a10620,a10622,a10624,
a10626,a10628,a10630,a10632,a10634,a10636,a10638,a10640,a10642,a10644,a10646,a10648,a10650,a10652,a10654,
a10656,a10658,a10660,a10662,a10664,a10666,a10668,a10670,a10672,a10674,a10676,a10678,a10680,a10682,a10684,
a10686,a10688,a10690,a10692,a10694,a10696,a10698,a10700,a10702,a10704,a10706,a10708,a10710,a10712,a10714,
a10716,a10718,a10720,a10722,a10724,a10726,a10728,a10730,a10732,a10734,a10736,a10738,a10740,a10742,a10744,
a10746,a10748,a10750,a10752,a10754,a10756,a10758,a10760,a10762,a10764,a10766,a10768,a10770,a10772,a10774,
a10776,a10778,a10780,a10782,a10784,a10786,a10788,a10790,a10792,a10794,a10796,a10798,a10800,a10802,a10804,
a10806,a10808,a10810,a10812,a10814,a10816,a10818,a10820,a10822,a10824,a10826,a10828,a10830,a10832,a10834,
a10836,a10838,a10840,a10842,a10844,a10846,a10848,a10850,a10852,a10854,a10856,a10858,a10860,a10862,a10864,
a10866,a10868,a10870,a10872,a10874,a10876,a10878,a10880,a10882,a10884,a10886,a10888,a10890,a10892,a10894,
a10896,a10898,a10900,a10902,a10904,a10906,a10908,a10910,a10912,a10914,a10916,a10918,a10920,a10922,a10924,
a10926,a10928,a10930,a10932,a10934,a10936,a10938,a10940,a10942,a10944,a10946,a10948,a10950,a10952,a10954,
a10956,a10958,a10960,a10962,a10964,a10966,a10968,a10970,a10972,a10974,a10976,a10978,a10980,a10982,a10984,
a10986,a10988,a10990,a10992,a10994,a10996,a10998,a11000,a11002,a11004,a11006,a11008,a11010,a11012,a11014,
a11016,a11018,a11020,a11022,a11024,a11026,a11028,a11030,a11032,a11034,a11036,a11038,a11040,a11042,a11044,
a11046,a11048,a11050,a11052,a11054,a11056,a11058,a11060,a11062,a11064,a11066,a11068,a11070,a11072,a11074,
a11076,a11078,a11080,a11082,a11084,a11086,a11088,a11090,a11092,a11094,a11096,a11098,a11100,a11102,a11104,
a11106,a11108,a11110,a11112,a11114,a11116,a11118,a11120,a11122,a11124,a11126,a11128,a11130,a11132,a11134,
a11136,a11138,a11140,a11142,a11144,a11146,a11148,a11150,a11152,a11154,a11156,a11158,a11160,a11162,a11164,
a11166,a11168,a11170,a11172,a11174,a11176,a11178,a11180,a11182,a11184,a11186,a11188,a11190,a11192,a11194,
a11196,a11198,a11200,a11202,a11204,a11206,a11208,a11210,a11212,a11214,a11216,a11218,a11220,a11222,a11224,
a11226,a11228,a11230,a11232,a11234,a11236,a11238,a11240,a11242,a11244,a11246,a11248,a11250,a11252,a11254,
a11256,a11258,a11260,a11262,a11264,a11266,a11268,a11270,a11272,a11274,a11276,a11278,a11280,a11282,a11284,
a11286,a11288,a11290,a11292,a11294,a11296,a11298,a11300,a11302,a11304,a11306,a11308,a11310,a11312,a11314,
a11316,a11318,a11320,a11322,a11324,a11326,a11328,a11330,a11332,a11334,a11336,a11338,a11340,a11342,a11344,
a11346,a11348,a11350,a11352,a11354,a11356,a11358,a11360,a11362,a11364,a11366,a11368,a11370,a11372,a11374,
a11376,a11378,a11380,a11382,a11384,a11386,a11388,a11390,a11392,a11394,a11396,a11398,a11400,a11402,a11404,
a11406,a11408,a11410,a11412,a11414,a11416,a11418,a11420,a11422,a11424,a11426,a11428,a11430,a11432,a11434,
a11436,a11438,a11440,a11442,a11444,a11446,a11448,a11450,a11452,a11454,a11456,a11458,a11460,a11462,a11464,
a11466,a11468,a11470,a11472,a11474,a11476,a11478,a11480,a11482,a11484,a11486,a11488,a11490,a11492,a11494,
a11496,a11498,a11500,a11502,a11504,a11506,a11508,a11510,a11512,a11514,a11516,a11518,a11520,a11522,a11524,
a11526,a11528,a11530,a11532,a11534,a11536,a11538,a11540,a11542,a11544,a11546,a11548,a11550,a11552,a11554,
a11556,a11558,a11560,a11562,a11564,a11566,a11568,a11570,a11572,a11574,a11576,a11578,a11580,a11582,a11584,
a11586,a11588,a11590,a11592,a11594,a11596,a11598,a11600,a11602,a11604,a11606,a11608,a11610,a11612,a11614,
a11616,a11618,a11620,a11622,a11624,a11626,a11628,a11630,a11632,a11634,a11636,a11638,a11640,a11642,a11644,
a11646,a11648,a11650,a11652,a11654,a11656,a11658,a11660,a11662,a11664,a11666,a11668,a11670,a11672,a11674,
a11676,a11678,a11680,a11682,a11684,a11686,a11688,a11690,a11692,a11694,a11696,a11698,a11700,a11702,a11704,
a11706,a11708,a11710,a11712,a11714,a11716,a11718,a11720,a11722,a11724,a11726,a11728,a11730,a11732,a11734,
a11736,a11738,a11740,a11742,a11744,a11746,a11748,a11750,a11752,a11754,a11756,a11758,a11760,a11762,a11764,
a11766,a11768,a11770,a11772,a11774,a11776,a11778,a11780,a11782,a11784,a11786,a11788,a11790,a11792,a11794,
a11796,a11798,a11800,a11802,a11804,a11806,a11808,a11810,a11812,a11814,a11816,a11818,a11820,a11822,a11824,
a11826,a11828,a11830,a11832,a11834,a11836,a11838,a11840,a11842,a11844,a11846,a11848,a11850,a11852,a11854,
a11856,a11858,a11860,a11862,a11864,a11866,a11868,a11870,a11872,a11874,a11876,a11878,a11880,a11882,a11884,
a11886,a11888,a11890,a11892,a11894,a11896,a11898,a11900,a11902,a11904,a11906,a11908,a11910,a11912,a11914,
a11916,a11918,a11920,a11922,a11924,a11926,a11928,a11930,a11932,a11934,a11936,a11938,a11940,a11942,a11944,
a11946,a11948,a11950,a11952,a11954,a11956,a11958,a11960,a11962,a11964,a11966,a11968,a11970,a11972,a11974,
a11976,a11978,a11980,a11982,a11984,a11986,a11988,a11990,a11992,a11994,a11996,a11998,a12000,a12002,a12004,
a12006,a12008,a12010,a12012,a12014,a12016,a12018,a12020,a12022,a12024,a12026,a12028,a12030,a12032,a12034,
a12036,a12038,a12040,a12042,a12044,a12046,a12048,a12050,a12052,a12054,a12056,a12058,a12060,a12062,a12064,
a12066,a12068,a12070,a12072,a12074,a12076,a12078,a12080,a12082,a12084,a12086,a12088,a12090,a12092,a12094,
a12096,a12098,a12100,a12102,a12104,a12106,a12108,a12110,a12112,a12114,a12116,a12118,a12120,a12122,a12124,
a12126,a12128,a12130,a12132,a12134,a12136,a12138,a12140,a12142,a12144,a12146,a12148,a12150,a12152,a12154,
a12156,a12158,a12160,a12162,a12164,a12166,a12168,a12170,a12172,a12174,a12176,a12178,a12180,a12182,a12184,
a12186,a12188,a12190,a12192,a12194,a12196,a12198,a12200,a12202,a12204,a12206,a12208,a12210,a12212,a12214,
a12216,a12218,a12220,a12222,a12224,a12226,a12228,a12230,a12232,a12234,a12236,a12238,a12240,a12242,a12244,
a12246,a12248,a12250,a12252,a12254,a12256,a12258,a12260,a12262,a12264,a12266,a12268,a12270,a12272,a12274,
a12276,a12278,a12280,a12282,a12284,a12286,a12288,a12290,a12292,a12294,a12296,a12298,a12300,a12302,a12304,
a12306,a12308,a12310,a12312,a12314,a12316,a12318,a12320,a12322,a12324,a12326,a12328,a12330,a12332,a12334,
a12336,a12338,a12340,a12342,a12344,a12346,a12348,a12350,a12352,a12354,a12356,a12358,a12360,a12362,a12364,
a12366,a12368,a12370,a12372,a12374,a12376,a12378,a12380,a12382,a12384,a12386,a12388,a12390,a12392,a12394,
a12396,a12398,a12400,a12402,a12404,a12406,a12408,a12410,a12412,a12414,a12416,a12418,a12420,a12422,a12424,
a12426,a12428,a12430,a12432,a12434,a12436,a12438,a12440,a12442,a12444,a12446,a12448,a12450,a12452,a12454,
a12456,a12458,a12460,a12462,a12464,a12466,a12468,a12470,a12472,a12474,a12476,a12478,a12480,a12482,a12484,
a12486,a12488,a12490,a12492,a12494,a12496,a12498,a12500,a12502,a12504,a12506,a12508,a12510,a12512,a12514,
a12516,a12518,a12520,a12522,a12524,a12526,a12528,a12530,a12532,a12534,a12536,a12538,a12540,a12542,a12544,
a12546,a12548,a12550,a12552,a12554,a12556,a12558,a12560,a12562,a12564,a12566,a12568,a12570,a12572,a12574,
a12576,a12578,a12580,a12582,a12584,a12586,a12588,a12590,a12592,a12594,a12596,a12598,a12600,a12602,a12604,
a12606,a12608,a12610,a12612,a12614,a12616,a12618,a12620,a12622,a12624,a12626,a12628,a12630,a12632,a12634,
a12636,a12638,a12640,a12642,a12644,a12646,a12648,a12650,a12652,a12654,a12656,a12658,a12660,a12662,a12664,
a12666,a12668,a12670,a12672,a12674,a12676,a12678,a12680,a12682,a12684,a12686,a12688,a12690,a12692,a12694,
a12696,a12698,a12700,a12702,a12704,a12706,a12708,a12710,a12712,a12714,a12716,a12718,a12720,a12722,a12724,
a12726,a12728,a12730,a12732,a12734,a12736,a12738,a12740,a12742,a12744,a12746,a12748,a12750,a12752,a12754,
a12756,a12758,a12760,a12762,a12764,a12766,a12768,a12770,a12772,a12774,a12776,a12778,a12780,a12782,a12784,
a12786,a12788,a12790,a12792,a12794,a12796,a12798,a12800,a12802,a12804,a12806,a12808,a12810,a12812,a12814,
a12816,a12818,a12820,a12822,a12824,a12826,a12828,a12830,a12832,a12834,a12836,a12838,a12840,a12842,a12844,
a12846,a12848,a12850,a12852,a12854,a12856,a12858,a12860,a12862,a12864,a12866,a12868,a12870,a12872,a12874,
a12876,a12878,a12880,a12882,a12884,a12886,a12888,a12890,a12892,a12894,a12896,a12898,a12900,a12902,a12904,
a12906,a12908,a12910,a12912,a12914,a12916,a12918,a12920,a12922,a12924,a12926,a12928,a12930,a12932,a12934,
a12936,a12938,a12940,a12942,a12944,a12946,a12948,a12950,a12952,a12954,a12956,a12958,a12960,a12962,a12964,
a12966,a12968,a12970,a12972,a12974,a12976,a12978,a12980,a12982,a12984,a12986,a12988,a12990,a12992,a12994,
a12996,a12998,a13000,a13002,a13004,a13006,a13008,a13010,a13012,a13014,a13016,a13018,a13020,a13022,a13024,
a13026,a13028,a13030,a13032,a13034,a13036,a13038,a13040,a13042,a13044,a13046,a13048,a13050,a13052,a13054,
a13056,a13058,a13060,a13062,a13064,a13066,a13068,a13070,a13072,a13074,a13076,a13078,a13080,a13082,a13084,
a13086,a13088,a13090,a13092,a13094,a13096,a13098,a13100,a13102,a13104,a13106,a13108,a13110,a13112,a13114,
a13116,a13118,a13120,a13122,a13124,a13126,a13128,a13130,a13132,a13134,a13136,a13138,a13140,a13142,a13144,
a13146,a13148,a13150,a13152,a13154,a13156,a13158,a13160,a13162,a13164,a13166,a13168,a13170,a13172,a13174,
a13176,a13178,a13180,a13182,a13184,a13186,a13188,a13190,a13192,a13194,a13196,a13198,a13200,a13202,a13204,
a13206,a13208,a13210,a13212,a13214,a13216,a13218,a13220,a13222,a13224,a13226,a13228,a13230,a13232,a13234,
a13236,a13238,a13240,a13242,a13244,a13246,a13248,a13250,a13252,a13254,a13256,a13258,a13260,a13262,a13264,
a13266,a13268,a13270,a13272,a13274,a13276,a13278,a13280,a13282,a13284,a13286,a13288,a13290,a13292,a13294,
a13296,a13298,a13300,a13302,a13304,a13306,a13308,a13310,a13312,a13314,a13316,a13318,a13320,a13322,a13324,
a13326,a13328,a13330,a13332,a13334,a13336,a13338,a13340,a13342,a13344,a13346,a13348,a13350,a13352,a13354,
a13356,a13358,a13360,a13362,a13364,a13366,a13368,a13370,a13372,a13374,a13376,a13378,a13380,a13382,a13384,
a13386,a13388,a13390,a13392,a13394,a13396,a13398,a13400,a13402,a13404,a13406,a13408,a13410,a13412,a13414,
a13416,a13418,a13420,a13422,a13424,a13426,a13428,a13430,a13432,a13434,a13436,a13438,a13440,a13442,a13444,
a13446,a13448,a13450,a13452,a13454,a13456,a13458,a13460,a13462,a13464,a13466,a13468,a13470,a13472,a13474,
a13476,a13478,a13480,a13482,a13484,a13486,a13488,a13490,a13492,a13494,a13496,a13498,a13500,a13502,a13504,
a13506,a13508,a13510,a13512,a13514,a13516,a13518,a13520,a13522,a13524,a13526,a13528,a13530,a13532,a13534,
a13536,a13538,a13540,a13542,a13544,a13546,a13548,a13550,a13552,a13554,a13556,a13558,a13560,a13562,a13564,
a13566,a13568,a13570,a13572,a13574,a13576,a13578,a13580,a13582,a13584,a13586,a13588,a13590,a13592,a13594,
a13596,a13598,a13600,a13602,a13604,a13606,a13608,a13610,a13612,a13614,a13616,a13618,a13620,a13622,a13624,
a13626,a13628,a13630,a13632,a13634,a13636,a13638,a13640,a13642,a13644,a13646,a13648,a13650,a13652,a13654,
a13656,a13658,a13660,a13662,a13664,a13666,a13668,a13670,a13672,a13674,a13676,a13678,a13680,a13682,a13684,
a13686,a13688,a13690,a13692,a13694,a13696,a13698,a13700,a13702,a13704,a13706,a13708,a13710,a13712,a13714,
a13716,a13718,a13720,a13722,a13724,a13726,a13728,a13730,a13732,a13734,a13736,a13738,a13740,a13742,a13744,
a13746,a13748,a13750,a13752,a13754,a13756,a13758,a13760,a13762,a13764,a13766,a13768,a13770,a13772,a13774,
a13776,a13778,a13780,a13782,a13784,a13786,a13788,a13790,a13792,a13794,a13796,a13798,a13800,a13802,a13804,
a13806,a13808,a13810,a13812,a13814,a13816,a13818,a13820,a13822,a13824,a13826,a13828,a13830,a13832,a13834,
a13836,a13838,a13840,a13842,a13844,a13846,a13848,a13850,a13852,a13854,a13856,a13858,a13860,a13862,a13864,
a13866,a13868,a13870,a13872,a13874,a13876,a13878,a13880,a13882,a13884,a13886,a13888,a13890,a13892,a13894,
a13896,a13898,a13900,a13902,a13904,a13906,a13908,a13910,a13912,a13914,a13916,a13918,a13920,a13922,a13924,
a13926,a13928,a13930,a13932,a13934,a13936,a13938,a13940,a13942,a13944,a13946,a13948,a13950,a13952,a13954,
a13956,a13958,a13960,a13962,a13964,a13966,a13968,a13970,a13972,a13974,a13976,a13978,a13980,a13982,a13984,
a13986,a13988,a13990,a13992,a13994,a13996,a13998,a14000,a14002,a14004,a14006,a14008,a14010,a14012,a14014,
a14016,a14018,a14020,a14022,a14024,a14026,a14028,a14030,a14032,a14034,a14036,a14038,a14040,a14042,a14044,
a14046,a14048,a14050,a14052,a14054,a14056,a14058,a14060,a14062,a14064,a14066,a14068,a14070,a14072,a14074,
a14076,a14078,a14080,a14082,a14084,a14086,a14088,a14090,a14092,a14094,a14096,a14098,a14100,a14102,a14104,
a14106,a14108,a14110,a14112,a14114,a14116,a14118,a14120,a14122,a14124,a14126,a14128,a14130,a14132,a14134,
a14136,a14138,a14140,a14142,a14144,a14146,a14148,a14150,a14152,a14154,a14156,a14158,a14160,a14162,a14164,
a14166,a14168,a14170,a14172,a14174,a14176,a14178,a14180,a14182,a14184,a14186,a14188,a14190,a14192,a14194,
a14196,a14198,a14200,a14202,a14204,a14206,a14208,a14210,a14212,a14214,a14216,a14218,a14220,a14222,a14224,
a14226,a14228,a14230,a14232,a14234,a14236,a14238,a14240,a14242,a14244,a14246,a14248,a14250,a14252,a14254,
a14256,a14258,a14260,a14262,a14264,a14266,a14268,a14270,a14272,a14274,a14276,a14278,a14280,a14282,a14284,
a14286,a14288,a14290,a14292,a14294,a14296,a14298,a14300,a14302,a14304,a14306,a14308,a14310,a14312,a14314,
a14316,a14318,a14320,a14322,a14324,a14326,a14328,a14330,a14332,a14334,a14336,a14338,a14340,a14342,a14344,
a14346,a14348,a14350,a14352,a14354,a14356,a14358,a14360,a14362,a14364,a14366,a14368,a14370,a14372,a14374,
a14376,a14378,a14380,a14382,a14384,a14386,a14388,a14390,a14392,a14394,a14396,a14398,a14400,a14402,a14404,
a14406,a14408,a14410,a14412,a14414,a14416,a14418,a14420,a14422,a14424,a14426,a14428,a14430,a14432,a14434,
a14436,a14438,a14440,a14442,a14444,a14446,a14448,a14450,a14452,a14454,a14456,a14458,a14460,a14462,a14464,
a14466,a14468,a14470,a14472,a14474,a14476,a14478,a14480,a14482,a14484,a14486,a14488,a14490,a14492,a14494,
a14496,a14498,a14500,a14502,a14504,a14506,a14508,a14510,a14512,a14514,a14516,a14518,a14520,a14522,a14524,
a14526,a14528,a14530,a14532,a14534,a14536,a14538,a14540,a14542,a14544,a14546,a14548,a14550,a14552,a14554,
a14556,a14558,a14560,a14562,a14564,a14566,a14568,a14570,a14572,a14574,a14576,a14578,a14580,a14582,a14584,
a14586,a14588,a14590,a14592,a14594,a14596,a14598,a14600,a14602,a14604,a14606,a14608,a14610,a14612,a14614,
a14616,a14618,a14620,a14622,a14624,a14626,a14628,a14630,a14632,a14634,a14636,a14638,a14640,a14642,a14644,
a14646,a14648,a14650,a14652,a14654,a14656,a14658,a14660,a14662,a14664,a14666,a14668,a14670,a14672,a14674,
a14676,a14678,a14680,a14682,a14684,a14686,a14688,a14690,a14692,a14694,a14696,a14698,a14700,a14702,a14704,
a14706,a14708,a14710,a14712,a14714,a14716,a14718,a14720,a14722,a14724,a14726,a14728,a14730,a14732,a14734,
a14736,a14738,a14740,a14742,a14744,a14746,a14748,a14750,a14752,a14754,a14756,a14758,a14760,a14762,a14764,
a14766,a14768,a14770,a14772,a14774,a14776,a14778,a14780,a14782,a14784,a14786,a14788,a14790,a14792,a14794,
a14796,a14798,a14800,a14802,a14804,a14806,a14808,a14810,a14812,a14814,a14816,a14818,a14820,a14822,a14824,
a14826,a14828,a14830,a14832,a14834,a14836,a14838,a14840,a14842,a14844,a14846,a14848,a14850,a14852,a14854,
a14856,a14858,a14860,a14862,a14864,a14866,a14868,a14870,a14872,a14874,a14876,a14878,a14880,a14882,a14884,
a14886,a14888,a14890,a14892,a14894,a14896,a14898,a14900,a14902,a14904,a14906,a14908,a14910,a14912,a14914,
a14916,a14918,a14920,a14922,a14924,a14926,a14928,a14930,a14932,a14934,a14936,a14938,a14940,a14942,a14944,
a14946,a14948,a14950,a14952,a14954,a14956,a14958,a14960,a14962,a14964,a14966,a14968,a14970,a14972,a14974,
a14976,a14978,a14980,a14982,a14984,a14986,a14988,a14990,a14992,a14994,a14996,a14998,a15000,a15002,a15004,
a15006,a15008,a15010,a15012,a15014,a15016,a15018,a15020,a15022,a15024,a15026,a15028,a15030,a15032,a15034,
a15036,a15038,a15040,a15042,a15044,a15046,a15048,a15050,a15052,a15054,a15056,a15058,a15060,a15062,a15064,
a15066,a15068,a15070,a15072,a15074,a15076,a15078,a15080,a15082,a15084,a15086,a15088,a15090,a15092,a15094,
a15096,a15098,a15100,a15102,a15104,a15106,a15108,a15110,a15112,a15114,a15116,a15118,a15120,a15122,a15124,
a15126,a15128,a15130,a15132,a15134,a15136,a15138,a15140,a15142,a15144,a15146,a15148,a15150,a15152,a15154,
a15156,a15158,a15160,a15162,a15164,a15166,a15168,a15170,a15172,a15174,a15176,a15178,a15180,a15182,a15184,
a15186,a15188,a15190,a15192,a15194,a15196,a15198,a15200,a15202,a15204,a15206,a15208,a15210,a15212,a15214,
a15216,a15218,a15220,a15222,a15224,a15226,a15228,a15230,a15232,a15234,a15236,a15238,a15240,a15242,a15244,
a15246,a15248,a15250,a15252,a15254,a15256,a15258,a15260,a15262,a15264,a15266,a15268,a15270,a15272,a15274,
a15276,a15278,a15280,a15282,a15284,a15286,a15288,a15290,a15292,a15294,a15296,a15298,a15300,a15302,a15304,
a15306,a15308,a15310,a15312,a15314,a15316,a15318,a15320,a15322,a15324,a15326,a15328,a15330,a15332,a15334,
a15336,a15338,a15340,a15342,a15344,a15346,a15348,a15350,a15352,a15354,a15356,a15358,a15360,a15362,a15364,
a15366,a15368,a15370,a15372,a15374,a15376,a15378,a15380,a15382,a15384,a15386,a15388,a15390,a15392,a15394,
a15396,a15398,a15400,a15402,a15404,a15406,a15408,a15410,a15412,a15414,a15416,a15418,a15420,a15422,a15424,
a15426,a15428,a15430,a15432,a15434,a15436,a15438,a15440,a15442,a15444,a15446,a15448,a15450,a15452,a15454,
a15456,a15458,a15460,a15462,a15464,a15466,a15468,a15470,a15472,a15474,a15476,a15478,a15480,a15482,a15484,
a15486,a15488,a15490,a15492,a15494,a15496,a15498,a15500,a15502,a15504,a15506,a15508,a15510,a15512,a15514,
a15516,a15518,a15520,a15522,a15524,a15526,a15528,a15530,a15532,a15534,a15536,a15538,a15540,a15542,a15544,
a15546,a15548,a15550,a15552,a15554,a15556,a15558,a15560,a15562,a15564,a15566,a15568,a15570,a15572,a15574,
a15576,a15578,a15580,a15582,a15584,a15586,a15588,a15590,a15592,a15594,a15596,a15598,a15600,a15602,a15604,
a15606,a15608,a15610,a15612,a15614,a15616,a15618,a15620,a15622,a15624,a15626,a15628,a15630,a15632,a15634,
a15636,a15638,a15640,a15642,a15644,a15646,a15648,a15650,a15652,a15654,a15656,a15658,a15660,a15662,a15664,
a15666,a15668,a15670,a15672,a15674,a15676,a15678,a15680,a15682,a15684,a15686,a15688,a15690,a15692,a15694,
a15696,a15698,a15700,a15702,a15704,a15706,a15708,a15710,a15712,a15714,a15716,a15718,a15720,a15722,a15724,
a15726,a15728,a15730,a15732,a15734,a15736,a15738,a15740,a15742,a15744,a15746,a15748,a15750,a15752,a15754,
a15756,a15758,a15760,a15762,a15764,a15766,a15768,a15770,a15772,a15774,a15776,a15778,a15780,a15782,a15784,
a15786,a15788,a15790,a15792,a15794,a15796,a15798,a15800,a15802,a15804,a15806,a15808,a15810,a15812,a15814,
a15816,a15818,a15820,a15822,a15824,a15826,a15828,a15830,a15832,a15834,a15836,a15838,a15840,a15842,a15844,
a15846,a15848,a15850,a15852,a15854,a15856,a15858,a15860,a15862,a15864,a15866,a15868,a15870,a15872,a15874,
a15876,a15878,a15880,a15882,a15884,a15886,a15888,a15890,a15892,a15894,a15896,a15898,a15900,a15902,a15904,
a15906,a15908,a15910,a15912,a15914,a15916,a15918,a15920,a15922,a15924,a15926,a15928,a15930,a15932,a15934,
a15936,a15938,a15940,a15942,a15944,a15946,a15948,a15950,a15952,a15954,a15956,a15958,a15960,a15962,a15964,
a15966,a15968,a15970,a15972,a15974,a15976,a15978,a15980,a15982,a15984,a15986,a15988,a15990,a15992,a15994,
a15996,a15998,a16000,a16002,a16004,a16006,a16008,a16010,a16012,a16014,a16016,a16018,a16020,a16022,a16024,
a16026,a16028,a16030,a16032,a16034,a16036,a16038,a16040,a16042,a16044,a16046,a16048,a16050,a16052,a16054,
a16056,a16058,a16060,a16062,a16064,a16066,a16068,a16070,a16072,a16074,a16076,a16078,a16080,a16082,a16084,
a16086,a16088,a16090,a16092,a16094,a16096,a16098,a16100,a16102,a16104,a16106,a16108,a16110,a16112,a16114,
a16116,a16118,a16120,a16122,a16124,a16126,a16128,a16130,a16132,a16134,a16136,a16138,a16140,a16142,a16144,
a16146,a16148,a16150,a16152,a16154,a16156,a16158,a16160,a16162,a16164,a16166,a16168,a16170,a16172,a16174,
a16176,a16178,a16180,a16182,a16184,a16186,a16188,a16190,a16192,a16194,a16196,a16198,a16200,a16202,a16204,
a16206,a16208,a16210,a16212,a16214,a16216,a16218,a16220,a16222,a16224,a16226,a16228,a16230,a16232,a16234,
a16236,a16238,a16240,a16242,a16244,a16246,a16248,a16250,a16252,a16254,a16256,a16258,a16260,a16262,a16264,
a16266,a16268,a16270,a16272,a16274,a16276,a16278,a16280,a16282,a16284,a16286,a16288,a16290,a16292,a16294,
a16296,a16298,a16300,a16302,a16304,a16306,a16308,a16310,a16312,a16314,a16316,a16318,a16320,a16322,a16324,
a16326,a16328,a16330,a16332,a16334,a16336,a16338,a16340,a16342,a16344,a16346,a16348,a16350,a16352,a16354,
a16356,a16358,a16360,a16362,a16364,a16366,a16368,a16370,a16372,a16374,a16376,a16378,a16380,a16382,a16384,
a16386,a16388,a16390,a16392,a16394,a16396,a16398,a16400,a16402,a16404,a16406,a16408,a16410,a16412,a16414,
a16416,a16418,a16420,a16422,a16424,a16426,a16428,a16430,a16432,a16434,a16436,a16438,a16440,a16442,a16444,
a16446,a16448,a16450,a16452,a16454,a16456,a16458,a16460,a16462,a16464,a16466,a16468,a16470,a16472,a16474,
a16476,a16478,a16480,a16482,a16484,a16486,a16488,a16490,a16492,a16494,a16496,a16498,a16500,a16502,a16504,
a16506,a16508,a16510,a16512,a16514,a16516,a16518,a16520,a16522,a16524,a16526,a16528,a16530,a16532,a16534,
a16536,a16538,a16540,a16542,a16544,a16546,a16548,a16550,a16552,a16554,a16556,a16558,a16560,a16562,a16564,
a16566,a16568,a16570,a16572,a16574,a16576,a16578,a16580,a16582,a16584,a16586,a16588,a16590,a16592,a16594,
a16596,a16598,a16600,a16602,a16604,a16606,a16608,a16610,a16612,a16614,a16616,a16618,a16620,a16622,a16624,
a16626,a16628,a16630,a16632,a16634,a16636,a16638,a16640,a16642,a16644,a16646,a16648,a16650,a16652,a16654,
a16656,a16658,a16660,a16662,a16664,a16666,a16668,a16670,a16672,a16674,a16676,a16678,a16680,a16682,a16684,
a16686,a16688,a16690,a16692,a16694,a16696,a16698,a16700,a16702,a16704,a16706,a16708,a16710,a16712,a16714,
a16716,a16718,a16720,a16722,a16724,a16726,a16728,a16730,a16732,a16734,a16736,a16738,a16740,a16742,a16744,
a16746,a16748,a16750,a16752,a16754,a16756,a16758,a16760,a16762,a16764,a16766,a16768,a16770,a16772,a16774,
a16776,a16778,a16780,a16782,a16784,a16786,a16788,a16790,a16792,a16794,a16796,a16798,a16800,a16802,a16804,
a16806,a16808,a16810,a16812,a16814,a16816,a16818,a16820,a16822,a16824,a16826,a16828,a16830,a16832,a16834,
a16836,a16838,a16840,a16842,a16844,a16846,a16848,a16850,a16852,a16854,a16856,a16858,a16860,a16862,a16864,
a16866,a16868,a16870,a16872,a16874,a16878,p0;

reg l580,l582,l584,l586,l588,l590,l592,l594,l596,l598,l600,l602,l604,l606,l608,
l610,l612,l614,l616,l618,l620,l622,l624,l626,l628,l630,l632,l634,l636,l638,
l640,l642,l644,l646,l648,l650,l652,l654,l656,l658,l660,l662,l664,l666,l668,
l670,l672,l674,l676,l678,l680,l682,l684,l686,l688,l690,l692,l694,l696,l698,
l700,l702,l704,l706,l708,l710,l712,l714,l716,l718,l720,l722,l724,l726,l728,
l730,l732,l734,l736,l738,l740,l742,l744,l746,l748,l750,l752,l754,l756,l758,
l760,l762,l764,l766,l768,l770,l772,l774,l776,l778,l780,l782,l784,l786,l788,
l790,l792,l794,l796,l798,l800,l802,l804,l806,l808,l810,l812,l814,l816,l818,
l820,l822,l824,l826,l828,l830,l832,l834,l836,l838,l840,l842,l844,l846,l848,
l850,l852,l854,l856,l858,l860,l862,l864,l866,l868,l870,l872,l874,l876,l878,
l880,l882,l884,l886,l888,l890,l892,l894,l896,l898,l900,l902,l904,l906,l908,
l910,l912,l914,l916,l918,l920,l922,l924,l926,l928,l930,l932,l934,l936,l938,
l940,l942,l944,l946,l948,l950,l952,l954,l956,l958,l960,l962,l964,l966,l968,
l970,l972,l974,l976,l978,l980,l982,l984,l986,l988,l990,l992,l994,l996,l998,
l1000,l1002,l1004,l1006,l1008,l1010,l1012,l1014,l1016,l1018,l1020,l1022,l1024,l1026,l1028,
l1030,l1032,l1034,l1036,l1038,l1040,l1042,l1044,l1046,l1048,l1050,l1052,l1054,l1056,l1058,
l1060,l1062,l1064,l1066,l1068,l1070,l1072,l1074,l1076,l1078,l1080,l1082,l1084,l1086,l1088,
l1090,l1092,l1094,l1096,l1098,l1100,l1102,l1104,l1106,l1108,l1110,l1112,l1114,l1116,l1118,
l1120,l1122,l1124,l1126,l1128,l1130,l1132,l1134,l1136,l1138,l1140,l1142,l1144,l1146,l1148,
l1150,l1152,l1154,l1156,l1158,l1160,l1162,l1164,l1166,l1168,l1170,l1172,l1174,l1176,l1178,
l1180,l1182,l1184,l1186,l1188,l1190,l1192,l1194,l1196,l1198,l1200,l1202,l1204,l1206,l1208,
l1210,l1212,l1214,l1216,l1218,l1220,l1222,l1224,l1226,l1228,l1230,l1232,l1234,l1236,l1238,
l1240,l1242,l1244,l1246,l1248,l1250,l1252,l1254,l1256,l1258,l1260,l1262,l1264,l1266,l1268,
l1270,l1272,l1274,l1276,l1278,l1280,l1282,l1284,l1286,l1288,l1290,l1292,l1294,l1296,l1298,
l1300,l1302,l1304,l1306,l1308,l1310,l1312,l1314,l1316,l1318,l1320,l1322,l1324,l1326,l1328;

initial
begin
   l580 = 0;
   l582 = 0;
   l584 = 0;
   l586 = 0;
   l588 = 0;
   l590 = 0;
   l592 = 0;
   l594 = 0;
   l596 = 0;
   l598 = 0;
   l600 = 0;
   l602 = 0;
   l604 = 0;
   l606 = 0;
   l608 = 0;
   l610 = 0;
   l612 = 0;
   l614 = 0;
   l616 = 0;
   l618 = 0;
   l620 = 0;
   l622 = 0;
   l624 = 0;
   l626 = 0;
   l628 = 0;
   l630 = 0;
   l632 = 0;
   l634 = 0;
   l636 = 0;
   l638 = 0;
   l640 = 0;
   l642 = 0;
   l644 = 0;
   l646 = 0;
   l648 = 0;
   l650 = 0;
   l652 = 0;
   l654 = 0;
   l656 = 0;
   l658 = 0;
   l660 = 0;
   l662 = 0;
   l664 = 0;
   l666 = 0;
   l668 = 0;
   l670 = 0;
   l672 = 0;
   l674 = 0;
   l676 = 0;
   l678 = 0;
   l680 = 0;
   l682 = 0;
   l684 = 0;
   l686 = 0;
   l688 = 0;
   l690 = 0;
   l692 = 0;
   l694 = 0;
   l696 = 0;
   l698 = 0;
   l700 = 0;
   l702 = 0;
   l704 = 0;
   l706 = 0;
   l708 = 0;
   l710 = 0;
   l712 = 0;
   l714 = 0;
   l716 = 0;
   l718 = 0;
   l720 = 0;
   l722 = 0;
   l724 = 0;
   l726 = 0;
   l728 = 0;
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
   l802 = 0;
   l804 = 0;
   l806 = 0;
   l808 = 0;
   l810 = 0;
   l812 = 0;
   l814 = 0;
   l816 = 0;
   l818 = 0;
   l820 = 0;
   l822 = 0;
   l824 = 0;
   l826 = 0;
   l828 = 0;
   l830 = 0;
   l832 = 0;
   l834 = 0;
   l836 = 0;
   l838 = 0;
   l840 = 0;
   l842 = 0;
   l844 = 0;
   l846 = 0;
   l848 = 0;
   l850 = 0;
   l852 = 0;
   l854 = 0;
   l856 = 0;
   l858 = 0;
   l860 = 0;
   l862 = 0;
   l864 = 0;
   l866 = 0;
   l868 = 0;
   l870 = 0;
   l872 = 0;
   l874 = 0;
   l876 = 0;
   l878 = 0;
   l880 = 0;
   l882 = 0;
   l884 = 0;
   l886 = 0;
   l888 = 0;
   l890 = 0;
   l892 = 0;
   l894 = 0;
   l896 = 0;
   l898 = 0;
   l900 = 0;
   l902 = 0;
   l904 = 0;
   l906 = 0;
   l908 = 0;
   l910 = 0;
   l912 = 0;
   l914 = 0;
   l916 = 0;
   l918 = 0;
   l920 = 0;
   l922 = 0;
   l924 = 0;
   l926 = 0;
   l928 = 0;
   l930 = 0;
   l932 = 0;
   l934 = 0;
   l936 = 0;
   l938 = 0;
   l940 = 0;
   l942 = 0;
   l944 = 0;
   l946 = 0;
   l948 = 0;
   l950 = 0;
   l952 = 0;
   l954 = 0;
   l956 = 0;
   l958 = 0;
   l960 = 0;
   l962 = 0;
   l964 = 0;
   l966 = 0;
   l968 = 0;
   l970 = 0;
   l972 = 0;
   l974 = 0;
   l976 = 0;
   l978 = 0;
   l980 = 0;
   l982 = 0;
   l984 = 0;
   l986 = 0;
   l988 = 0;
   l990 = 0;
   l992 = 0;
   l994 = 0;
   l996 = 0;
   l998 = 0;
   l1000 = 0;
   l1002 = 0;
   l1004 = 0;
   l1006 = 0;
   l1008 = 0;
   l1010 = 0;
   l1012 = 0;
   l1014 = 0;
   l1016 = 0;
   l1018 = 0;
   l1020 = 0;
   l1022 = 0;
   l1024 = 0;
   l1026 = 0;
   l1028 = 0;
   l1030 = 0;
   l1032 = 0;
   l1034 = 0;
   l1036 = 0;
   l1038 = 0;
   l1040 = 0;
   l1042 = 0;
   l1044 = 0;
   l1046 = 0;
   l1048 = 0;
   l1050 = 0;
   l1052 = 0;
   l1054 = 0;
   l1056 = 0;
   l1058 = 0;
   l1060 = 0;
   l1062 = 0;
   l1064 = 0;
   l1066 = 0;
   l1068 = 0;
   l1070 = 0;
   l1072 = 0;
   l1074 = 0;
   l1076 = 0;
   l1078 = 0;
   l1080 = 0;
   l1082 = 0;
   l1084 = 0;
   l1086 = 0;
   l1088 = 0;
   l1090 = 0;
   l1092 = 0;
   l1094 = 0;
   l1096 = 0;
   l1098 = 0;
   l1100 = 0;
   l1102 = 0;
   l1104 = 0;
   l1106 = 0;
   l1108 = 0;
   l1110 = 0;
   l1112 = 0;
   l1114 = 0;
   l1116 = 0;
   l1118 = 0;
   l1120 = 0;
   l1122 = 0;
   l1124 = 0;
   l1126 = 0;
   l1128 = 0;
   l1130 = 0;
   l1132 = 0;
   l1134 = 0;
   l1136 = 0;
   l1138 = 0;
   l1140 = 0;
   l1142 = 0;
   l1144 = 0;
   l1146 = 0;
   l1148 = 0;
   l1150 = 0;
   l1152 = 0;
   l1154 = 0;
   l1156 = 0;
   l1158 = 0;
   l1160 = 0;
   l1162 = 0;
   l1164 = 0;
   l1166 = 0;
   l1168 = 0;
   l1170 = 0;
   l1172 = 0;
   l1174 = 0;
   l1176 = 0;
   l1178 = 0;
   l1180 = 0;
   l1182 = 0;
   l1184 = 0;
   l1186 = 0;
   l1188 = 0;
   l1190 = 0;
   l1192 = 0;
   l1194 = 0;
   l1196 = 0;
   l1198 = 0;
   l1200 = 0;
   l1202 = 0;
   l1204 = 0;
   l1206 = 0;
   l1208 = 0;
   l1210 = 0;
   l1212 = 0;
   l1214 = 0;
   l1216 = 0;
   l1218 = 0;
   l1220 = 0;
   l1222 = 0;
   l1224 = 0;
   l1226 = 0;
   l1228 = 0;
   l1230 = 0;
   l1232 = 0;
   l1234 = 0;
   l1236 = 0;
   l1238 = 0;
   l1240 = 0;
   l1242 = 0;
   l1244 = 0;
   l1246 = 0;
   l1248 = 0;
   l1250 = 0;
   l1252 = 0;
   l1254 = 0;
   l1256 = 0;
   l1258 = 0;
   l1260 = 0;
   l1262 = 0;
   l1264 = 0;
   l1266 = 0;
   l1268 = 0;
   l1270 = 0;
   l1272 = 0;
   l1274 = 0;
   l1276 = 0;
   l1278 = 0;
   l1280 = 0;
   l1282 = 0;
   l1284 = 0;
   l1286 = 0;
   l1288 = 0;
   l1290 = 0;
   l1292 = 0;
   l1294 = 0;
   l1296 = 0;
   l1298 = 0;
   l1300 = 0;
   l1302 = 0;
   l1304 = 0;
   l1306 = 0;
   l1308 = 0;
   l1310 = 0;
   l1312 = 0;
   l1314 = 0;
   l1316 = 0;
   l1318 = 0;
   l1320 = 0;
   l1322 = 0;
   l1324 = 0;
   l1326 = 0;
   l1328 = 0;
end

always @(posedge i2)
   l580 <= i2;

always @(posedge i4)
   l582 <= i4;

always @(posedge i6)
   l584 <= i6;

always @(posedge i8)
   l586 <= i8;

always @(posedge i10)
   l588 <= i10;

always @(posedge i12)
   l590 <= i12;

always @(posedge i14)
   l592 <= i14;

always @(posedge i16)
   l594 <= i16;

always @(posedge i18)
   l596 <= i18;

always @(posedge i20)
   l598 <= i20;

always @(posedge i22)
   l600 <= i22;

always @(posedge i24)
   l602 <= i24;

always @(posedge i26)
   l604 <= i26;

always @(posedge i28)
   l606 <= i28;

always @(posedge i30)
   l608 <= i30;

always @(posedge i32)
   l610 <= i32;

always @(posedge i34)
   l612 <= i34;

always @(posedge i36)
   l614 <= i36;

always @(posedge i38)
   l616 <= i38;

always @(posedge i40)
   l618 <= i40;

always @(posedge i42)
   l620 <= i42;

always @(posedge i44)
   l622 <= i44;

always @(posedge i46)
   l624 <= i46;

always @(posedge i48)
   l626 <= i48;

always @(posedge i50)
   l628 <= i50;

always @(posedge i52)
   l630 <= i52;

always @(posedge i54)
   l632 <= i54;

always @(posedge i56)
   l634 <= i56;

always @(posedge i58)
   l636 <= i58;

always @(posedge i60)
   l638 <= i60;

always @(posedge i62)
   l640 <= i62;

always @(posedge i64)
   l642 <= i64;

always @(posedge i66)
   l644 <= i66;

always @(posedge i68)
   l646 <= i68;

always @(posedge i70)
   l648 <= i70;

always @(posedge i72)
   l650 <= i72;

always @(posedge i74)
   l652 <= i74;

always @(posedge i76)
   l654 <= i76;

always @(posedge i78)
   l656 <= i78;

always @(posedge i80)
   l658 <= i80;

always @(posedge i82)
   l660 <= i82;

always @(posedge i84)
   l662 <= i84;

always @(posedge i86)
   l664 <= i86;

always @(posedge i88)
   l666 <= i88;

always @(posedge i90)
   l668 <= i90;

always @(posedge i92)
   l670 <= i92;

always @(posedge i94)
   l672 <= i94;

always @(posedge i96)
   l674 <= i96;

always @(posedge i98)
   l676 <= i98;

always @(posedge i100)
   l678 <= i100;

always @(posedge i102)
   l680 <= i102;

always @(posedge i104)
   l682 <= i104;

always @(posedge i106)
   l684 <= i106;

always @(posedge i108)
   l686 <= i108;

always @(posedge i110)
   l688 <= i110;

always @(posedge i112)
   l690 <= i112;

always @(posedge i114)
   l692 <= i114;

always @(posedge i116)
   l694 <= i116;

always @(posedge i118)
   l696 <= i118;

always @(posedge i120)
   l698 <= i120;

always @(posedge i122)
   l700 <= i122;

always @(posedge i124)
   l702 <= i124;

always @(posedge i126)
   l704 <= i126;

always @(posedge i128)
   l706 <= i128;

always @(posedge i130)
   l708 <= i130;

always @(posedge i132)
   l710 <= i132;

always @(posedge i134)
   l712 <= i134;

always @(posedge i136)
   l714 <= i136;

always @(posedge i138)
   l716 <= i138;

always @(posedge i140)
   l718 <= i140;

always @(posedge i142)
   l720 <= i142;

always @(posedge i144)
   l722 <= i144;

always @(posedge i146)
   l724 <= i146;

always @(posedge i148)
   l726 <= i148;

always @(posedge i150)
   l728 <= i150;

always @(posedge i152)
   l730 <= i152;

always @(posedge i154)
   l732 <= i154;

always @(posedge i156)
   l734 <= i156;

always @(posedge i158)
   l736 <= i158;

always @(posedge i160)
   l738 <= i160;

always @(posedge i162)
   l740 <= i162;

always @(posedge i164)
   l742 <= i164;

always @(posedge a1386)
   l744 <= a1386;

always @(posedge a1402)
   l746 <= a1402;

always @(posedge i166)
   l748 <= i166;

always @(posedge i168)
   l750 <= i168;

always @(posedge a1430)
   l752 <= a1430;

always @(posedge i170)
   l754 <= i170;

always @(posedge i172)
   l756 <= i172;

always @(posedge a1474)
   l758 <= a1474;

always @(posedge a1490)
   l760 <= a1490;

always @(posedge i174)
   l762 <= i174;

always @(posedge i176)
   l764 <= i176;

always @(posedge a1510)
   l766 <= a1510;

always @(posedge i178)
   l768 <= i178;

always @(posedge i180)
   l770 <= i180;

always @(posedge a1554)
   l772 <= a1554;

always @(posedge a1570)
   l774 <= a1570;

always @(posedge i182)
   l776 <= i182;

always @(posedge i184)
   l778 <= i184;

always @(posedge a1590)
   l780 <= a1590;

always @(posedge i186)
   l782 <= i186;

always @(posedge i188)
   l784 <= i188;

always @(posedge a1634)
   l786 <= a1634;

always @(posedge a1650)
   l788 <= a1650;

always @(posedge i190)
   l790 <= i190;

always @(posedge i192)
   l792 <= i192;

always @(posedge a1670)
   l794 <= a1670;

always @(posedge a1778)
   l796 <= a1778;

always @(posedge a1802)
   l798 <= a1802;

always @(posedge a1830)
   l800 <= a1830;

always @(posedge i194)
   l802 <= i194;

always @(posedge i196)
   l804 <= i196;

always @(posedge i198)
   l806 <= i198;

always @(posedge i200)
   l808 <= i200;

always @(posedge i202)
   l810 <= i202;

always @(posedge a1842)
   l812 <= a1842;

always @(posedge a1996)
   l814 <= a1996;

always @(posedge a2006)
   l816 <= a2006;

always @(posedge a2016)
   l818 <= a2016;

always @(posedge a2026)
   l820 <= a2026;

always @(posedge i204)
   l822 <= i204;

always @(posedge i206)
   l824 <= i206;

always @(posedge a2084)
   l826 <= a2084;

always @(posedge a2100)
   l828 <= a2100;

always @(posedge i208)
   l830 <= i208;

always @(posedge i210)
   l832 <= i210;

always @(posedge a2128)
   l834 <= a2128;

always @(posedge i212)
   l836 <= i212;

always @(posedge i214)
   l838 <= i214;

always @(posedge a2172)
   l840 <= a2172;

always @(posedge a2188)
   l842 <= a2188;

always @(posedge i216)
   l844 <= i216;

always @(posedge i218)
   l846 <= i218;

always @(posedge a2208)
   l848 <= a2208;

always @(posedge i220)
   l850 <= i220;

always @(posedge i222)
   l852 <= i222;

always @(posedge a2252)
   l854 <= a2252;

always @(posedge a2268)
   l856 <= a2268;

always @(posedge i224)
   l858 <= i224;

always @(posedge i226)
   l860 <= i226;

always @(posedge a2288)
   l862 <= a2288;

always @(posedge i228)
   l864 <= i228;

always @(posedge i230)
   l866 <= i230;

always @(posedge a2332)
   l868 <= a2332;

always @(posedge a2348)
   l870 <= a2348;

always @(posedge i232)
   l872 <= i232;

always @(posedge i234)
   l874 <= i234;

always @(posedge a2368)
   l876 <= a2368;

always @(posedge a2476)
   l878 <= a2476;

always @(posedge a2500)
   l880 <= a2500;

always @(posedge a2528)
   l882 <= a2528;

always @(posedge i236)
   l884 <= i236;

always @(posedge i238)
   l886 <= i238;

always @(posedge i240)
   l888 <= i240;

always @(posedge i242)
   l890 <= i242;

always @(posedge i244)
   l892 <= i244;

always @(posedge a2540)
   l894 <= a2540;

always @(posedge a2694)
   l896 <= a2694;

always @(posedge a2704)
   l898 <= a2704;

always @(posedge a2714)
   l900 <= a2714;

always @(posedge a2724)
   l902 <= a2724;

always @(posedge i246)
   l904 <= i246;

always @(posedge i248)
   l906 <= i248;

always @(posedge a2782)
   l908 <= a2782;

always @(posedge a2798)
   l910 <= a2798;

always @(posedge i250)
   l912 <= i250;

always @(posedge i252)
   l914 <= i252;

always @(posedge a2826)
   l916 <= a2826;

always @(posedge i254)
   l918 <= i254;

always @(posedge i256)
   l920 <= i256;

always @(posedge a2870)
   l922 <= a2870;

always @(posedge a2886)
   l924 <= a2886;

always @(posedge i258)
   l926 <= i258;

always @(posedge i260)
   l928 <= i260;

always @(posedge a2906)
   l930 <= a2906;

always @(posedge i262)
   l932 <= i262;

always @(posedge i264)
   l934 <= i264;

always @(posedge a2950)
   l936 <= a2950;

always @(posedge a2966)
   l938 <= a2966;

always @(posedge i266)
   l940 <= i266;

always @(posedge i268)
   l942 <= i268;

always @(posedge a2986)
   l944 <= a2986;

always @(posedge i270)
   l946 <= i270;

always @(posedge i272)
   l948 <= i272;

always @(posedge a3030)
   l950 <= a3030;

always @(posedge a3046)
   l952 <= a3046;

always @(posedge i274)
   l954 <= i274;

always @(posedge i276)
   l956 <= i276;

always @(posedge a3066)
   l958 <= a3066;

always @(posedge a3174)
   l960 <= a3174;

always @(posedge a3198)
   l962 <= a3198;

always @(posedge a3226)
   l964 <= a3226;

always @(posedge i278)
   l966 <= i278;

always @(posedge i280)
   l968 <= i280;

always @(posedge i282)
   l970 <= i282;

always @(posedge i284)
   l972 <= i284;

always @(posedge i286)
   l974 <= i286;

always @(posedge a3238)
   l976 <= a3238;

always @(posedge a3392)
   l978 <= a3392;

always @(posedge a3402)
   l980 <= a3402;

always @(posedge a3412)
   l982 <= a3412;

always @(posedge a3422)
   l984 <= a3422;

always @(posedge i288)
   l986 <= i288;

always @(posedge i290)
   l988 <= i290;

always @(posedge a3480)
   l990 <= a3480;

always @(posedge a3496)
   l992 <= a3496;

always @(posedge i292)
   l994 <= i292;

always @(posedge i294)
   l996 <= i294;

always @(posedge a3524)
   l998 <= a3524;

always @(posedge i296)
   l1000 <= i296;

always @(posedge i298)
   l1002 <= i298;

always @(posedge a3568)
   l1004 <= a3568;

always @(posedge a3584)
   l1006 <= a3584;

always @(posedge i300)
   l1008 <= i300;

always @(posedge i302)
   l1010 <= i302;

always @(posedge a3604)
   l1012 <= a3604;

always @(posedge i304)
   l1014 <= i304;

always @(posedge i306)
   l1016 <= i306;

always @(posedge a3648)
   l1018 <= a3648;

always @(posedge a3664)
   l1020 <= a3664;

always @(posedge i308)
   l1022 <= i308;

always @(posedge i310)
   l1024 <= i310;

always @(posedge a3684)
   l1026 <= a3684;

always @(posedge i312)
   l1028 <= i312;

always @(posedge i314)
   l1030 <= i314;

always @(posedge a3728)
   l1032 <= a3728;

always @(posedge a3744)
   l1034 <= a3744;

always @(posedge i316)
   l1036 <= i316;

always @(posedge i318)
   l1038 <= i318;

always @(posedge a3764)
   l1040 <= a3764;

always @(posedge a3872)
   l1042 <= a3872;

always @(posedge a3896)
   l1044 <= a3896;

always @(posedge a3924)
   l1046 <= a3924;

always @(posedge i320)
   l1048 <= i320;

always @(posedge i322)
   l1050 <= i322;

always @(posedge i324)
   l1052 <= i324;

always @(posedge i326)
   l1054 <= i326;

always @(posedge i328)
   l1056 <= i328;

always @(posedge a3936)
   l1058 <= a3936;

always @(posedge a4090)
   l1060 <= a4090;

always @(posedge a4100)
   l1062 <= a4100;

always @(posedge a4110)
   l1064 <= a4110;

always @(posedge a4120)
   l1066 <= a4120;

always @(posedge i330)
   l1068 <= i330;

always @(posedge a4126)
   l1070 <= a4126;

always @(posedge i332)
   l1072 <= i332;

always @(posedge i334)
   l1074 <= i334;

always @(posedge i336)
   l1076 <= i336;

always @(posedge i338)
   l1078 <= i338;

always @(posedge i340)
   l1080 <= i340;

always @(posedge i342)
   l1082 <= i342;

always @(posedge i344)
   l1084 <= i344;

always @(posedge i346)
   l1086 <= i346;

always @(posedge i348)
   l1088 <= i348;

always @(posedge i350)
   l1090 <= i350;

always @(posedge i352)
   l1092 <= i352;

always @(posedge i354)
   l1094 <= i354;

always @(posedge i356)
   l1096 <= i356;

always @(posedge i358)
   l1098 <= i358;

always @(posedge i360)
   l1100 <= i360;

always @(posedge i362)
   l1102 <= i362;

always @(posedge i364)
   l1104 <= i364;

always @(posedge i366)
   l1106 <= i366;

always @(posedge i368)
   l1108 <= i368;

always @(posedge i370)
   l1110 <= i370;

always @(posedge i372)
   l1112 <= i372;

always @(posedge i374)
   l1114 <= i374;

always @(posedge i376)
   l1116 <= i376;

always @(posedge i378)
   l1118 <= i378;

always @(posedge i380)
   l1120 <= i380;

always @(posedge i382)
   l1122 <= i382;

always @(posedge i384)
   l1124 <= i384;

always @(posedge i386)
   l1126 <= i386;

always @(posedge i388)
   l1128 <= i388;

always @(posedge i390)
   l1130 <= i390;

always @(posedge i392)
   l1132 <= i392;

always @(posedge i394)
   l1134 <= i394;

always @(posedge i396)
   l1136 <= i396;

always @(posedge i398)
   l1138 <= i398;

always @(posedge i400)
   l1140 <= i400;

always @(posedge i402)
   l1142 <= i402;

always @(posedge i404)
   l1144 <= i404;

always @(posedge i406)
   l1146 <= i406;

always @(posedge i408)
   l1148 <= i408;

always @(posedge i410)
   l1150 <= i410;

always @(posedge i412)
   l1152 <= i412;

always @(posedge i414)
   l1154 <= i414;

always @(posedge i416)
   l1156 <= i416;

always @(posedge i418)
   l1158 <= i418;

always @(posedge i420)
   l1160 <= i420;

always @(posedge i422)
   l1162 <= i422;

always @(posedge i424)
   l1164 <= i424;

always @(posedge i426)
   l1166 <= i426;

always @(posedge i428)
   l1168 <= i428;

always @(posedge i430)
   l1170 <= i430;

always @(posedge i432)
   l1172 <= i432;

always @(posedge i434)
   l1174 <= i434;

always @(posedge i436)
   l1176 <= i436;

always @(posedge i438)
   l1178 <= i438;

always @(posedge i440)
   l1180 <= i440;

always @(posedge i442)
   l1182 <= i442;

always @(posedge i444)
   l1184 <= i444;

always @(posedge i446)
   l1186 <= i446;

always @(posedge i448)
   l1188 <= i448;

always @(posedge i450)
   l1190 <= i450;

always @(posedge i452)
   l1192 <= i452;

always @(posedge i454)
   l1194 <= i454;

always @(posedge i456)
   l1196 <= i456;

always @(posedge i458)
   l1198 <= i458;

always @(posedge i460)
   l1200 <= i460;

always @(posedge i462)
   l1202 <= i462;

always @(posedge i464)
   l1204 <= i464;

always @(posedge i466)
   l1206 <= i466;

always @(posedge i468)
   l1208 <= i468;

always @(posedge i470)
   l1210 <= i470;

always @(posedge i472)
   l1212 <= i472;

always @(posedge i474)
   l1214 <= i474;

always @(posedge i476)
   l1216 <= i476;

always @(posedge i478)
   l1218 <= i478;

always @(posedge i480)
   l1220 <= i480;

always @(posedge i482)
   l1222 <= i482;

always @(posedge i484)
   l1224 <= i484;

always @(posedge i486)
   l1226 <= i486;

always @(posedge i488)
   l1228 <= i488;

always @(posedge i490)
   l1230 <= i490;

always @(posedge i492)
   l1232 <= i492;

always @(posedge i494)
   l1234 <= i494;

always @(posedge i496)
   l1236 <= i496;

always @(posedge i498)
   l1238 <= i498;

always @(posedge i500)
   l1240 <= i500;

always @(posedge i502)
   l1242 <= i502;

always @(posedge i504)
   l1244 <= i504;

always @(posedge i506)
   l1246 <= i506;

always @(posedge i508)
   l1248 <= i508;

always @(posedge i510)
   l1250 <= i510;

always @(posedge i512)
   l1252 <= i512;

always @(posedge i514)
   l1254 <= i514;

always @(posedge i516)
   l1256 <= i516;

always @(posedge i518)
   l1258 <= i518;

always @(posedge i520)
   l1260 <= i520;

always @(posedge i522)
   l1262 <= i522;

always @(posedge i524)
   l1264 <= i524;

always @(posedge i526)
   l1266 <= i526;

always @(posedge i528)
   l1268 <= i528;

always @(posedge i530)
   l1270 <= i530;

always @(posedge i532)
   l1272 <= i532;

always @(posedge i534)
   l1274 <= i534;

always @(posedge i536)
   l1276 <= i536;

always @(posedge i538)
   l1278 <= i538;

always @(posedge i540)
   l1280 <= i540;

always @(posedge i542)
   l1282 <= i542;

always @(posedge i544)
   l1284 <= i544;

always @(posedge i546)
   l1286 <= i546;

always @(posedge i548)
   l1288 <= i548;

always @(posedge i550)
   l1290 <= i550;

always @(posedge i552)
   l1292 <= i552;

always @(posedge i554)
   l1294 <= i554;

always @(posedge i556)
   l1296 <= i556;

always @(posedge i558)
   l1298 <= i558;

always @(posedge i560)
   l1300 <= i560;

always @(posedge i562)
   l1302 <= i562;

always @(posedge i564)
   l1304 <= i564;

always @(posedge i566)
   l1306 <= i566;

always @(posedge a4134)
   l1308 <= a4134;

always @(posedge a4144)
   l1310 <= a4144;

always @(posedge a4152)
   l1312 <= a4152;

always @(posedge i568)
   l1314 <= i568;

always @(posedge a4154)
   l1316 <= a4154;

always @(posedge i572)
   l1318 <= i572;

always @(posedge i574)
   l1320 <= i574;

always @(posedge i576)
   l1322 <= i576;

always @(posedge i578)
   l1324 <= i578;

always @(posedge a16876)
   l1326 <= a16876;

always @(posedge c1)
   l1328 <= c1;


assign a1386 = a1384 & l1328;
assign a1402 = ~a1400 & l1328;
assign a1430 = ~a1428 & l1328;
assign a1474 = a1472 & l1328;
assign a1490 = ~a1488 & l1328;
assign a1510 = ~a1508 & l1328;
assign a1554 = a1552 & l1328;
assign a1570 = ~a1568 & l1328;
assign a1590 = ~a1588 & l1328;
assign a1634 = a1632 & l1328;
assign a1650 = ~a1648 & l1328;
assign a1670 = ~a1668 & l1328;
assign a1778 = a1776 & l1328;
assign a1802 = ~a1800 & l1328;
assign a1830 = ~a1828 & l1328;
assign a1842 = ~a1840 & l1328;
assign a1996 = a1994 & l1328;
assign a2006 = a2004 & l1328;
assign a2016 = a2014 & l1328;
assign a2026 = a2024 & l1328;
assign a2084 = a2082 & l1328;
assign a2100 = ~a2098 & l1328;
assign a2128 = ~a2126 & l1328;
assign a2172 = a2170 & l1328;
assign a2188 = ~a2186 & l1328;
assign a2208 = ~a2206 & l1328;
assign a2252 = a2250 & l1328;
assign a2268 = ~a2266 & l1328;
assign a2288 = ~a2286 & l1328;
assign a2332 = a2330 & l1328;
assign a2348 = ~a2346 & l1328;
assign a2368 = ~a2366 & l1328;
assign a2476 = a2474 & l1328;
assign a2500 = ~a2498 & l1328;
assign a2528 = ~a2526 & l1328;
assign a2540 = ~a2538 & l1328;
assign a2694 = a2692 & l1328;
assign a2704 = a2702 & l1328;
assign a2714 = a2712 & l1328;
assign a2724 = a2722 & l1328;
assign a2782 = a2780 & l1328;
assign a2798 = ~a2796 & l1328;
assign a2826 = ~a2824 & l1328;
assign a2870 = a2868 & l1328;
assign a2886 = ~a2884 & l1328;
assign a2906 = ~a2904 & l1328;
assign a2950 = a2948 & l1328;
assign a2966 = ~a2964 & l1328;
assign a2986 = ~a2984 & l1328;
assign a3030 = a3028 & l1328;
assign a3046 = ~a3044 & l1328;
assign a3066 = ~a3064 & l1328;
assign a3174 = a3172 & l1328;
assign a3198 = ~a3196 & l1328;
assign a3226 = ~a3224 & l1328;
assign a3238 = ~a3236 & l1328;
assign a3392 = a3390 & l1328;
assign a3402 = a3400 & l1328;
assign a3412 = a3410 & l1328;
assign a3422 = a3420 & l1328;
assign a3480 = a3478 & l1328;
assign a3496 = ~a3494 & l1328;
assign a3524 = ~a3522 & l1328;
assign a3568 = a3566 & l1328;
assign a3584 = ~a3582 & l1328;
assign a3604 = ~a3602 & l1328;
assign a3648 = a3646 & l1328;
assign a3664 = ~a3662 & l1328;
assign a3684 = ~a3682 & l1328;
assign a3728 = a3726 & l1328;
assign a3744 = ~a3742 & l1328;
assign a3764 = ~a3762 & l1328;
assign a3872 = a3870 & l1328;
assign a3896 = ~a3894 & l1328;
assign a3924 = ~a3922 & l1328;
assign a3936 = ~a3934 & l1328;
assign a4090 = a4088 & l1328;
assign a4100 = a4098 & l1328;
assign a4110 = a4108 & l1328;
assign a4120 = a4118 & l1328;
assign a4126 = ~a4124 & l1328;
assign a4134 = ~a4132 & l1328;
assign a4144 = ~a4142 & l1328;
assign a4152 = ~a4150 & l1328;
assign a4154 = ~a4128 & l1328;
assign a16876 = a16874 & l1328;
assign c1 = 1;
assign a1330 = l752 & ~l750;
assign a1332 = l800 & l798;
assign a1334 = a1332 & ~l796;
assign a1336 = a1334 & a1330;
assign a1338 = ~l752 & l750;
assign a1340 = a1338 & a1334;
assign a1342 = l800 & ~l798;
assign a1344 = a1342 & l796;
assign a1346 = a1344 & a1338;
assign a1348 = l742 & ~l740;
assign a1350 = a1332 & l796;
assign a1352 = a1350 & a1338;
assign a1354 = a1352 & a1348;
assign a1356 = ~l742 & ~l740;
assign a1358 = l752 & l750;
assign a1360 = a1342 & ~l796;
assign a1362 = a1360 & a1358;
assign a1364 = a1362 & a1356;
assign a1366 = a1360 & a1330;
assign a1368 = a1366 & a1348;
assign a1370 = a1360 & l802;
assign a1372 = ~a1370 & l744;
assign a1374 = a1372 & ~a1368;
assign a1376 = a1374 & ~a1364;
assign a1378 = ~a1376 & ~a1354;
assign a1380 = ~a1378 & ~a1346;
assign a1382 = ~a1380 & ~a1340;
assign a1384 = ~a1382 & ~a1336;
assign a1388 = ~a1370 & l746;
assign a1390 = a1388 & ~a1368;
assign a1392 = a1390 & ~a1364;
assign a1394 = ~a1392 & ~a1354;
assign a1396 = ~a1394 & ~a1346;
assign a1398 = ~a1396 & ~a1340;
assign a1400 = a1398 & ~a1336;
assign a1404 = ~l742 & l740;
assign a1406 = ~l800 & ~l798;
assign a1408 = a1406 & ~l796;
assign a1410 = a1408 & a1338;
assign a1412 = a1410 & a1404;
assign a1414 = ~l800 & l798;
assign a1416 = a1414 & ~l796;
assign a1418 = a1416 & a1338;
assign a1420 = a1418 & a1356;
assign a1422 = a1404 & a1352;
assign a1424 = ~a1422 & ~l752;
assign a1426 = a1424 & ~a1420;
assign a1428 = a1426 & ~a1412;
assign a1432 = l766 & ~l764;
assign a1434 = a1432 & a1334;
assign a1436 = ~l766 & l764;
assign a1438 = a1436 & a1334;
assign a1440 = a1436 & a1344;
assign a1442 = l756 & ~l754;
assign a1444 = a1436 & a1350;
assign a1446 = a1444 & a1442;
assign a1448 = ~l756 & ~l754;
assign a1450 = l766 & l764;
assign a1452 = a1450 & a1360;
assign a1454 = a1452 & a1448;
assign a1456 = a1432 & a1360;
assign a1458 = a1456 & a1442;
assign a1460 = ~a1370 & l758;
assign a1462 = a1460 & ~a1458;
assign a1464 = a1462 & ~a1454;
assign a1466 = ~a1464 & ~a1446;
assign a1468 = ~a1466 & ~a1440;
assign a1470 = ~a1468 & ~a1438;
assign a1472 = ~a1470 & ~a1434;
assign a1476 = ~a1370 & l760;
assign a1478 = a1476 & ~a1458;
assign a1480 = a1478 & ~a1454;
assign a1482 = ~a1480 & ~a1446;
assign a1484 = ~a1482 & ~a1440;
assign a1486 = ~a1484 & ~a1438;
assign a1488 = a1486 & ~a1434;
assign a1492 = ~l756 & l754;
assign a1494 = a1436 & a1408;
assign a1496 = a1494 & a1492;
assign a1498 = a1436 & a1416;
assign a1500 = a1498 & a1448;
assign a1502 = a1492 & a1444;
assign a1504 = ~a1502 & ~l766;
assign a1506 = a1504 & ~a1500;
assign a1508 = a1506 & ~a1496;
assign a1512 = l780 & ~l778;
assign a1514 = a1512 & a1334;
assign a1516 = ~l780 & l778;
assign a1518 = a1516 & a1334;
assign a1520 = a1516 & a1344;
assign a1522 = l770 & ~l768;
assign a1524 = a1516 & a1350;
assign a1526 = a1524 & a1522;
assign a1528 = ~l770 & ~l768;
assign a1530 = l780 & l778;
assign a1532 = a1530 & a1360;
assign a1534 = a1532 & a1528;
assign a1536 = a1512 & a1360;
assign a1538 = a1536 & a1522;
assign a1540 = ~a1370 & l772;
assign a1542 = a1540 & ~a1538;
assign a1544 = a1542 & ~a1534;
assign a1546 = ~a1544 & ~a1526;
assign a1548 = ~a1546 & ~a1520;
assign a1550 = ~a1548 & ~a1518;
assign a1552 = ~a1550 & ~a1514;
assign a1556 = ~a1370 & l774;
assign a1558 = a1556 & ~a1538;
assign a1560 = a1558 & ~a1534;
assign a1562 = ~a1560 & ~a1526;
assign a1564 = ~a1562 & ~a1520;
assign a1566 = ~a1564 & ~a1518;
assign a1568 = a1566 & ~a1514;
assign a1572 = ~l770 & l768;
assign a1574 = a1516 & a1408;
assign a1576 = a1574 & a1572;
assign a1578 = a1516 & a1416;
assign a1580 = a1578 & a1528;
assign a1582 = a1572 & a1524;
assign a1584 = ~a1582 & ~l780;
assign a1586 = a1584 & ~a1580;
assign a1588 = a1586 & ~a1576;
assign a1592 = l794 & ~l792;
assign a1594 = a1592 & a1334;
assign a1596 = ~l794 & l792;
assign a1598 = a1596 & a1334;
assign a1600 = a1596 & a1344;
assign a1602 = l784 & ~l782;
assign a1604 = a1596 & a1350;
assign a1606 = a1604 & a1602;
assign a1608 = ~l784 & ~l782;
assign a1610 = l794 & l792;
assign a1612 = a1610 & a1360;
assign a1614 = a1612 & a1608;
assign a1616 = a1592 & a1360;
assign a1618 = a1616 & a1602;
assign a1620 = ~a1370 & l786;
assign a1622 = a1620 & ~a1618;
assign a1624 = a1622 & ~a1614;
assign a1626 = ~a1624 & ~a1606;
assign a1628 = ~a1626 & ~a1600;
assign a1630 = ~a1628 & ~a1598;
assign a1632 = ~a1630 & ~a1594;
assign a1636 = ~a1370 & l788;
assign a1638 = a1636 & ~a1618;
assign a1640 = a1638 & ~a1614;
assign a1642 = ~a1640 & ~a1606;
assign a1644 = ~a1642 & ~a1600;
assign a1646 = ~a1644 & ~a1598;
assign a1648 = a1646 & ~a1594;
assign a1652 = ~l784 & l782;
assign a1654 = a1596 & a1408;
assign a1656 = a1654 & a1652;
assign a1658 = a1596 & a1416;
assign a1660 = a1658 & a1608;
assign a1662 = a1652 & a1604;
assign a1664 = ~a1662 & ~l794;
assign a1666 = a1664 & ~a1660;
assign a1668 = a1666 & ~a1656;
assign a1672 = ~l814 & l808;
assign a1674 = ~a1436 & ~a1338;
assign a1676 = a1674 & ~a1516;
assign a1678 = a1436 & a1338;
assign a1680 = ~a1678 & ~a1516;
assign a1682 = ~a1680 & ~a1674;
assign a1684 = ~a1682 & ~a1596;
assign a1686 = ~a1684 & ~a1676;
assign a1688 = ~a1686 & a1408;
assign a1690 = a1688 & ~a1672;
assign a1692 = ~a1348 & a1330;
assign a1694 = ~a1692 & a1334;
assign a1696 = ~a1442 & a1432;
assign a1698 = ~a1696 & a1694;
assign a1700 = ~a1522 & a1512;
assign a1702 = ~a1700 & a1698;
assign a1704 = ~a1602 & a1592;
assign a1706 = ~a1704 & a1702;
assign a1708 = ~a1356 & a1338;
assign a1710 = ~a1708 & a1416;
assign a1712 = ~a1448 & a1436;
assign a1714 = ~a1712 & a1710;
assign a1716 = ~a1528 & a1516;
assign a1718 = ~a1716 & a1714;
assign a1720 = ~a1608 & a1596;
assign a1722 = ~a1720 & a1718;
assign a1724 = ~a1652 & a1596;
assign a1726 = ~a1572 & a1516;
assign a1728 = ~a1492 & a1436;
assign a1730 = ~a1404 & a1338;
assign a1732 = ~a1730 & a1416;
assign a1734 = a1732 & ~a1728;
assign a1736 = a1734 & ~a1726;
assign a1738 = a1736 & ~a1724;
assign a1740 = ~a1602 & a1596;
assign a1742 = ~a1522 & a1516;
assign a1744 = ~a1348 & a1338;
assign a1746 = ~a1442 & a1436;
assign a1748 = ~a1746 & ~a1744;
assign a1750 = a1748 & ~a1742;
assign a1752 = a1750 & ~a1740;
assign a1754 = ~a1730 & ~a1728;
assign a1756 = a1754 & ~a1726;
assign a1758 = a1756 & ~a1724;
assign a1760 = ~a1758 & ~a1752;
assign a1762 = ~a1760 & ~a1342;
assign a1764 = a1762 & a1350;
assign a1766 = a1764 & ~a1406;
assign a1768 = ~a1766 & l796;
assign a1770 = ~a1768 & ~a1738;
assign a1772 = ~a1770 & ~a1722;
assign a1774 = a1772 & ~a1706;
assign a1776 = a1774 & ~a1690;
assign a1780 = a1344 & ~l810;
assign a1782 = a1406 & l796;
assign a1784 = l800 & l796;
assign a1786 = a1784 & l810;
assign a1788 = ~a1786 & a1782;
assign a1790 = ~a1788 & ~l798;
assign a1792 = a1790 & ~a1780;
assign a1794 = ~a1792 & ~a1738;
assign a1796 = a1794 & ~a1722;
assign a1798 = ~a1796 & ~a1706;
assign a1800 = a1798 & ~a1690;
assign a1804 = a1344 & l810;
assign a1806 = ~a1742 & ~a1740;
assign a1808 = a1806 & ~a1746;
assign a1810 = a1808 & ~a1744;
assign a1812 = a1810 & a1350;
assign a1814 = ~a1812 & l800;
assign a1816 = ~a1814 & ~a1782;
assign a1818 = ~a1816 & ~a1804;
assign a1820 = ~a1818 & ~a1780;
assign a1822 = a1820 & ~a1738;
assign a1824 = a1822 & ~a1722;
assign a1826 = ~a1824 & ~a1706;
assign a1828 = ~a1826 & ~a1690;
assign a1832 = ~l820 & ~l818;
assign a1834 = ~a1832 & l816;
assign a1836 = a1834 & l814;
assign a1838 = a1836 & a1408;
assign a1840 = ~a1838 & ~l812;
assign a1844 = ~l818 & ~l816;
assign a1846 = a1844 & ~l814;
assign a1848 = l820 & ~l818;
assign a1850 = a1848 & ~l816;
assign a1852 = a1850 & ~l814;
assign a1854 = l818 & ~l816;
assign a1856 = a1854 & ~l814;
assign a1858 = l820 & l818;
assign a1860 = a1858 & ~l816;
assign a1862 = a1860 & ~l814;
assign a1864 = ~l818 & l816;
assign a1866 = a1864 & ~l814;
assign a1868 = a1848 & l816;
assign a1870 = a1868 & ~l814;
assign a1872 = l818 & l816;
assign a1874 = a1872 & ~l814;
assign a1876 = a1850 & l814;
assign a1878 = a1860 & l814;
assign a1880 = ~a1878 & a1864;
assign a1882 = ~a1880 & ~a1854;
assign a1884 = ~a1882 & ~a1876;
assign a1886 = ~a1884 & ~a1844;
assign a1888 = ~a1886 & l814;
assign a1890 = ~a1888 & ~a1874;
assign a1892 = ~a1890 & ~a1870;
assign a1894 = ~a1892 & ~a1866;
assign a1896 = ~a1894 & ~a1862;
assign a1898 = ~a1896 & ~a1856;
assign a1900 = ~a1898 & ~a1852;
assign a1902 = ~a1900 & ~a1846;
assign a1904 = ~a1902 & ~l820;
assign a1906 = a1832 & ~l816;
assign a1908 = a1906 & ~l814;
assign a1910 = l820 & ~l816;
assign a1912 = a1910 & ~l814;
assign a1914 = a1832 & l816;
assign a1916 = a1914 & ~l814;
assign a1918 = l820 & l816;
assign a1920 = a1918 & ~l814;
assign a1922 = a1906 & l814;
assign a1924 = ~l816 & l814;
assign a1926 = a1924 & ~a1848;
assign a1928 = a1926 & ~a1922;
assign a1930 = ~a1928 & ~a1920;
assign a1932 = ~l820 & l816;
assign a1934 = a1932 & ~l814;
assign a1936 = ~a1934 & a1930;
assign a1938 = ~a1936 & ~a1870;
assign a1940 = a1938 & ~a1916;
assign a1942 = ~a1940 & ~a1912;
assign a1944 = ~l820 & ~l816;
assign a1946 = a1944 & ~l814;
assign a1948 = ~a1946 & a1942;
assign a1950 = ~a1948 & l818;
assign a1952 = a1950 & ~a1852;
assign a1954 = a1952 & ~a1908;
assign a1956 = a1954 & a1904;
assign a1958 = ~l820 & l818;
assign a1960 = ~a1858 & ~l814;
assign a1962 = a1960 & ~a1958;
assign a1964 = a1848 & ~l814;
assign a1966 = ~a1964 & a1962;
assign a1968 = a1832 & ~l814;
assign a1970 = ~a1968 & a1966;
assign a1972 = ~a1970 & ~l816;
assign a1974 = ~a1972 & a1956;
assign a1976 = ~a1858 & ~l816;
assign a1978 = a1976 & ~a1958;
assign a1980 = a1978 & ~a1850;
assign a1982 = a1980 & ~a1906;
assign a1984 = ~a1982 & ~l814;
assign a1986 = ~a1984 & a1974;
assign a1988 = ~a1986 & l814;
assign a1990 = ~a1988 & a1408;
assign a1992 = ~a1408 & ~l814;
assign a1994 = ~a1992 & ~a1990;
assign a1998 = ~a1986 & l816;
assign a2000 = ~a1998 & a1408;
assign a2002 = ~a1408 & ~l816;
assign a2004 = ~a2002 & ~a2000;
assign a2008 = ~a1986 & l818;
assign a2010 = ~a2008 & a1408;
assign a2012 = ~a1408 & ~l818;
assign a2014 = ~a2012 & ~a2010;
assign a2018 = ~a1986 & ~l820;
assign a2020 = ~a2018 & a1408;
assign a2022 = ~a1408 & ~l820;
assign a2024 = ~a2022 & ~a2020;
assign a2028 = l834 & ~l832;
assign a2030 = l882 & l880;
assign a2032 = a2030 & ~l878;
assign a2034 = a2032 & a2028;
assign a2036 = ~l834 & l832;
assign a2038 = a2036 & a2032;
assign a2040 = l882 & ~l880;
assign a2042 = a2040 & l878;
assign a2044 = a2042 & a2036;
assign a2046 = l824 & ~l822;
assign a2048 = a2030 & l878;
assign a2050 = a2048 & a2036;
assign a2052 = a2050 & a2046;
assign a2054 = ~l824 & ~l822;
assign a2056 = l834 & l832;
assign a2058 = a2040 & ~l878;
assign a2060 = a2058 & a2056;
assign a2062 = a2060 & a2054;
assign a2064 = a2058 & a2028;
assign a2066 = a2064 & a2046;
assign a2068 = a2058 & l884;
assign a2070 = ~a2068 & l826;
assign a2072 = a2070 & ~a2066;
assign a2074 = a2072 & ~a2062;
assign a2076 = ~a2074 & ~a2052;
assign a2078 = ~a2076 & ~a2044;
assign a2080 = ~a2078 & ~a2038;
assign a2082 = ~a2080 & ~a2034;
assign a2086 = ~a2068 & l828;
assign a2088 = a2086 & ~a2066;
assign a2090 = a2088 & ~a2062;
assign a2092 = ~a2090 & ~a2052;
assign a2094 = ~a2092 & ~a2044;
assign a2096 = ~a2094 & ~a2038;
assign a2098 = a2096 & ~a2034;
assign a2102 = ~l824 & l822;
assign a2104 = ~l882 & ~l880;
assign a2106 = a2104 & ~l878;
assign a2108 = a2106 & a2036;
assign a2110 = a2108 & a2102;
assign a2112 = ~l882 & l880;
assign a2114 = a2112 & ~l878;
assign a2116 = a2114 & a2036;
assign a2118 = a2116 & a2054;
assign a2120 = a2102 & a2050;
assign a2122 = ~a2120 & ~l834;
assign a2124 = a2122 & ~a2118;
assign a2126 = a2124 & ~a2110;
assign a2130 = l848 & ~l846;
assign a2132 = a2130 & a2032;
assign a2134 = ~l848 & l846;
assign a2136 = a2134 & a2032;
assign a2138 = a2134 & a2042;
assign a2140 = l838 & ~l836;
assign a2142 = a2134 & a2048;
assign a2144 = a2142 & a2140;
assign a2146 = ~l838 & ~l836;
assign a2148 = l848 & l846;
assign a2150 = a2148 & a2058;
assign a2152 = a2150 & a2146;
assign a2154 = a2130 & a2058;
assign a2156 = a2154 & a2140;
assign a2158 = ~a2068 & l840;
assign a2160 = a2158 & ~a2156;
assign a2162 = a2160 & ~a2152;
assign a2164 = ~a2162 & ~a2144;
assign a2166 = ~a2164 & ~a2138;
assign a2168 = ~a2166 & ~a2136;
assign a2170 = ~a2168 & ~a2132;
assign a2174 = ~a2068 & l842;
assign a2176 = a2174 & ~a2156;
assign a2178 = a2176 & ~a2152;
assign a2180 = ~a2178 & ~a2144;
assign a2182 = ~a2180 & ~a2138;
assign a2184 = ~a2182 & ~a2136;
assign a2186 = a2184 & ~a2132;
assign a2190 = ~l838 & l836;
assign a2192 = a2134 & a2106;
assign a2194 = a2192 & a2190;
assign a2196 = a2134 & a2114;
assign a2198 = a2196 & a2146;
assign a2200 = a2190 & a2142;
assign a2202 = ~a2200 & ~l848;
assign a2204 = a2202 & ~a2198;
assign a2206 = a2204 & ~a2194;
assign a2210 = l862 & ~l860;
assign a2212 = a2210 & a2032;
assign a2214 = ~l862 & l860;
assign a2216 = a2214 & a2032;
assign a2218 = a2214 & a2042;
assign a2220 = l852 & ~l850;
assign a2222 = a2214 & a2048;
assign a2224 = a2222 & a2220;
assign a2226 = ~l852 & ~l850;
assign a2228 = l862 & l860;
assign a2230 = a2228 & a2058;
assign a2232 = a2230 & a2226;
assign a2234 = a2210 & a2058;
assign a2236 = a2234 & a2220;
assign a2238 = ~a2068 & l854;
assign a2240 = a2238 & ~a2236;
assign a2242 = a2240 & ~a2232;
assign a2244 = ~a2242 & ~a2224;
assign a2246 = ~a2244 & ~a2218;
assign a2248 = ~a2246 & ~a2216;
assign a2250 = ~a2248 & ~a2212;
assign a2254 = ~a2068 & l856;
assign a2256 = a2254 & ~a2236;
assign a2258 = a2256 & ~a2232;
assign a2260 = ~a2258 & ~a2224;
assign a2262 = ~a2260 & ~a2218;
assign a2264 = ~a2262 & ~a2216;
assign a2266 = a2264 & ~a2212;
assign a2270 = ~l852 & l850;
assign a2272 = a2214 & a2106;
assign a2274 = a2272 & a2270;
assign a2276 = a2214 & a2114;
assign a2278 = a2276 & a2226;
assign a2280 = a2270 & a2222;
assign a2282 = ~a2280 & ~l862;
assign a2284 = a2282 & ~a2278;
assign a2286 = a2284 & ~a2274;
assign a2290 = l876 & ~l874;
assign a2292 = a2290 & a2032;
assign a2294 = ~l876 & l874;
assign a2296 = a2294 & a2032;
assign a2298 = a2294 & a2042;
assign a2300 = l866 & ~l864;
assign a2302 = a2294 & a2048;
assign a2304 = a2302 & a2300;
assign a2306 = ~l866 & ~l864;
assign a2308 = l876 & l874;
assign a2310 = a2308 & a2058;
assign a2312 = a2310 & a2306;
assign a2314 = a2290 & a2058;
assign a2316 = a2314 & a2300;
assign a2318 = ~a2068 & l868;
assign a2320 = a2318 & ~a2316;
assign a2322 = a2320 & ~a2312;
assign a2324 = ~a2322 & ~a2304;
assign a2326 = ~a2324 & ~a2298;
assign a2328 = ~a2326 & ~a2296;
assign a2330 = ~a2328 & ~a2292;
assign a2334 = ~a2068 & l870;
assign a2336 = a2334 & ~a2316;
assign a2338 = a2336 & ~a2312;
assign a2340 = ~a2338 & ~a2304;
assign a2342 = ~a2340 & ~a2298;
assign a2344 = ~a2342 & ~a2296;
assign a2346 = a2344 & ~a2292;
assign a2350 = ~l866 & l864;
assign a2352 = a2294 & a2106;
assign a2354 = a2352 & a2350;
assign a2356 = a2294 & a2114;
assign a2358 = a2356 & a2306;
assign a2360 = a2350 & a2302;
assign a2362 = ~a2360 & ~l876;
assign a2364 = a2362 & ~a2358;
assign a2366 = a2364 & ~a2354;
assign a2370 = ~l896 & l890;
assign a2372 = ~a2134 & ~a2036;
assign a2374 = a2372 & ~a2214;
assign a2376 = a2134 & a2036;
assign a2378 = ~a2376 & ~a2214;
assign a2380 = ~a2378 & ~a2372;
assign a2382 = ~a2380 & ~a2294;
assign a2384 = ~a2382 & ~a2374;
assign a2386 = ~a2384 & a2106;
assign a2388 = a2386 & ~a2370;
assign a2390 = ~a2046 & a2028;
assign a2392 = ~a2390 & a2032;
assign a2394 = ~a2140 & a2130;
assign a2396 = ~a2394 & a2392;
assign a2398 = ~a2220 & a2210;
assign a2400 = ~a2398 & a2396;
assign a2402 = ~a2300 & a2290;
assign a2404 = ~a2402 & a2400;
assign a2406 = ~a2054 & a2036;
assign a2408 = ~a2406 & a2114;
assign a2410 = ~a2146 & a2134;
assign a2412 = ~a2410 & a2408;
assign a2414 = ~a2226 & a2214;
assign a2416 = ~a2414 & a2412;
assign a2418 = ~a2306 & a2294;
assign a2420 = ~a2418 & a2416;
assign a2422 = ~a2350 & a2294;
assign a2424 = ~a2270 & a2214;
assign a2426 = ~a2190 & a2134;
assign a2428 = ~a2102 & a2036;
assign a2430 = ~a2428 & a2114;
assign a2432 = a2430 & ~a2426;
assign a2434 = a2432 & ~a2424;
assign a2436 = a2434 & ~a2422;
assign a2438 = ~a2300 & a2294;
assign a2440 = ~a2220 & a2214;
assign a2442 = ~a2046 & a2036;
assign a2444 = ~a2140 & a2134;
assign a2446 = ~a2444 & ~a2442;
assign a2448 = a2446 & ~a2440;
assign a2450 = a2448 & ~a2438;
assign a2452 = ~a2428 & ~a2426;
assign a2454 = a2452 & ~a2424;
assign a2456 = a2454 & ~a2422;
assign a2458 = ~a2456 & ~a2450;
assign a2460 = ~a2458 & ~a2040;
assign a2462 = a2460 & a2048;
assign a2464 = a2462 & ~a2104;
assign a2466 = ~a2464 & l878;
assign a2468 = ~a2466 & ~a2436;
assign a2470 = ~a2468 & ~a2420;
assign a2472 = a2470 & ~a2404;
assign a2474 = a2472 & ~a2388;
assign a2478 = a2042 & ~l892;
assign a2480 = a2104 & l878;
assign a2482 = l882 & l878;
assign a2484 = a2482 & l892;
assign a2486 = ~a2484 & a2480;
assign a2488 = ~a2486 & ~l880;
assign a2490 = a2488 & ~a2478;
assign a2492 = ~a2490 & ~a2436;
assign a2494 = a2492 & ~a2420;
assign a2496 = ~a2494 & ~a2404;
assign a2498 = a2496 & ~a2388;
assign a2502 = a2042 & l892;
assign a2504 = ~a2440 & ~a2438;
assign a2506 = a2504 & ~a2444;
assign a2508 = a2506 & ~a2442;
assign a2510 = a2508 & a2048;
assign a2512 = ~a2510 & l882;
assign a2514 = ~a2512 & ~a2480;
assign a2516 = ~a2514 & ~a2502;
assign a2518 = ~a2516 & ~a2478;
assign a2520 = a2518 & ~a2436;
assign a2522 = a2520 & ~a2420;
assign a2524 = ~a2522 & ~a2404;
assign a2526 = ~a2524 & ~a2388;
assign a2530 = ~l902 & ~l900;
assign a2532 = ~a2530 & l898;
assign a2534 = a2532 & l896;
assign a2536 = a2534 & a2106;
assign a2538 = ~a2536 & ~l894;
assign a2542 = ~l900 & ~l898;
assign a2544 = a2542 & ~l896;
assign a2546 = l902 & ~l900;
assign a2548 = a2546 & ~l898;
assign a2550 = a2548 & ~l896;
assign a2552 = l900 & ~l898;
assign a2554 = a2552 & ~l896;
assign a2556 = l902 & l900;
assign a2558 = a2556 & ~l898;
assign a2560 = a2558 & ~l896;
assign a2562 = ~l900 & l898;
assign a2564 = a2562 & ~l896;
assign a2566 = a2546 & l898;
assign a2568 = a2566 & ~l896;
assign a2570 = l900 & l898;
assign a2572 = a2570 & ~l896;
assign a2574 = a2548 & l896;
assign a2576 = a2558 & l896;
assign a2578 = ~a2576 & a2562;
assign a2580 = ~a2578 & ~a2552;
assign a2582 = ~a2580 & ~a2574;
assign a2584 = ~a2582 & ~a2542;
assign a2586 = ~a2584 & l896;
assign a2588 = ~a2586 & ~a2572;
assign a2590 = ~a2588 & ~a2568;
assign a2592 = ~a2590 & ~a2564;
assign a2594 = ~a2592 & ~a2560;
assign a2596 = ~a2594 & ~a2554;
assign a2598 = ~a2596 & ~a2550;
assign a2600 = ~a2598 & ~a2544;
assign a2602 = ~a2600 & ~l902;
assign a2604 = a2530 & ~l898;
assign a2606 = a2604 & ~l896;
assign a2608 = l902 & ~l898;
assign a2610 = a2608 & ~l896;
assign a2612 = a2530 & l898;
assign a2614 = a2612 & ~l896;
assign a2616 = l902 & l898;
assign a2618 = a2616 & ~l896;
assign a2620 = a2604 & l896;
assign a2622 = ~l898 & l896;
assign a2624 = a2622 & ~a2546;
assign a2626 = a2624 & ~a2620;
assign a2628 = ~a2626 & ~a2618;
assign a2630 = ~l902 & l898;
assign a2632 = a2630 & ~l896;
assign a2634 = ~a2632 & a2628;
assign a2636 = ~a2634 & ~a2568;
assign a2638 = a2636 & ~a2614;
assign a2640 = ~a2638 & ~a2610;
assign a2642 = ~l902 & ~l898;
assign a2644 = a2642 & ~l896;
assign a2646 = ~a2644 & a2640;
assign a2648 = ~a2646 & l900;
assign a2650 = a2648 & ~a2550;
assign a2652 = a2650 & ~a2606;
assign a2654 = a2652 & a2602;
assign a2656 = ~l902 & l900;
assign a2658 = ~a2556 & ~l896;
assign a2660 = a2658 & ~a2656;
assign a2662 = a2546 & ~l896;
assign a2664 = ~a2662 & a2660;
assign a2666 = a2530 & ~l896;
assign a2668 = ~a2666 & a2664;
assign a2670 = ~a2668 & ~l898;
assign a2672 = ~a2670 & a2654;
assign a2674 = ~a2556 & ~l898;
assign a2676 = a2674 & ~a2656;
assign a2678 = a2676 & ~a2548;
assign a2680 = a2678 & ~a2604;
assign a2682 = ~a2680 & ~l896;
assign a2684 = ~a2682 & a2672;
assign a2686 = ~a2684 & l896;
assign a2688 = ~a2686 & a2106;
assign a2690 = ~a2106 & ~l896;
assign a2692 = ~a2690 & ~a2688;
assign a2696 = ~a2684 & l898;
assign a2698 = ~a2696 & a2106;
assign a2700 = ~a2106 & ~l898;
assign a2702 = ~a2700 & ~a2698;
assign a2706 = ~a2684 & l900;
assign a2708 = ~a2706 & a2106;
assign a2710 = ~a2106 & ~l900;
assign a2712 = ~a2710 & ~a2708;
assign a2716 = ~a2684 & ~l902;
assign a2718 = ~a2716 & a2106;
assign a2720 = ~a2106 & ~l902;
assign a2722 = ~a2720 & ~a2718;
assign a2726 = l916 & ~l914;
assign a2728 = l964 & l962;
assign a2730 = a2728 & ~l960;
assign a2732 = a2730 & a2726;
assign a2734 = ~l916 & l914;
assign a2736 = a2734 & a2730;
assign a2738 = l964 & ~l962;
assign a2740 = a2738 & l960;
assign a2742 = a2740 & a2734;
assign a2744 = l906 & ~l904;
assign a2746 = a2728 & l960;
assign a2748 = a2746 & a2734;
assign a2750 = a2748 & a2744;
assign a2752 = ~l906 & ~l904;
assign a2754 = l916 & l914;
assign a2756 = a2738 & ~l960;
assign a2758 = a2756 & a2754;
assign a2760 = a2758 & a2752;
assign a2762 = a2756 & a2726;
assign a2764 = a2762 & a2744;
assign a2766 = a2756 & l966;
assign a2768 = ~a2766 & l908;
assign a2770 = a2768 & ~a2764;
assign a2772 = a2770 & ~a2760;
assign a2774 = ~a2772 & ~a2750;
assign a2776 = ~a2774 & ~a2742;
assign a2778 = ~a2776 & ~a2736;
assign a2780 = ~a2778 & ~a2732;
assign a2784 = ~a2766 & l910;
assign a2786 = a2784 & ~a2764;
assign a2788 = a2786 & ~a2760;
assign a2790 = ~a2788 & ~a2750;
assign a2792 = ~a2790 & ~a2742;
assign a2794 = ~a2792 & ~a2736;
assign a2796 = a2794 & ~a2732;
assign a2800 = ~l906 & l904;
assign a2802 = ~l964 & ~l962;
assign a2804 = a2802 & ~l960;
assign a2806 = a2804 & a2734;
assign a2808 = a2806 & a2800;
assign a2810 = ~l964 & l962;
assign a2812 = a2810 & ~l960;
assign a2814 = a2812 & a2734;
assign a2816 = a2814 & a2752;
assign a2818 = a2800 & a2748;
assign a2820 = ~a2818 & ~l916;
assign a2822 = a2820 & ~a2816;
assign a2824 = a2822 & ~a2808;
assign a2828 = l930 & ~l928;
assign a2830 = a2828 & a2730;
assign a2832 = ~l930 & l928;
assign a2834 = a2832 & a2730;
assign a2836 = a2832 & a2740;
assign a2838 = l920 & ~l918;
assign a2840 = a2832 & a2746;
assign a2842 = a2840 & a2838;
assign a2844 = ~l920 & ~l918;
assign a2846 = l930 & l928;
assign a2848 = a2846 & a2756;
assign a2850 = a2848 & a2844;
assign a2852 = a2828 & a2756;
assign a2854 = a2852 & a2838;
assign a2856 = ~a2766 & l922;
assign a2858 = a2856 & ~a2854;
assign a2860 = a2858 & ~a2850;
assign a2862 = ~a2860 & ~a2842;
assign a2864 = ~a2862 & ~a2836;
assign a2866 = ~a2864 & ~a2834;
assign a2868 = ~a2866 & ~a2830;
assign a2872 = ~a2766 & l924;
assign a2874 = a2872 & ~a2854;
assign a2876 = a2874 & ~a2850;
assign a2878 = ~a2876 & ~a2842;
assign a2880 = ~a2878 & ~a2836;
assign a2882 = ~a2880 & ~a2834;
assign a2884 = a2882 & ~a2830;
assign a2888 = ~l920 & l918;
assign a2890 = a2832 & a2804;
assign a2892 = a2890 & a2888;
assign a2894 = a2832 & a2812;
assign a2896 = a2894 & a2844;
assign a2898 = a2888 & a2840;
assign a2900 = ~a2898 & ~l930;
assign a2902 = a2900 & ~a2896;
assign a2904 = a2902 & ~a2892;
assign a2908 = l944 & ~l942;
assign a2910 = a2908 & a2730;
assign a2912 = ~l944 & l942;
assign a2914 = a2912 & a2730;
assign a2916 = a2912 & a2740;
assign a2918 = l934 & ~l932;
assign a2920 = a2912 & a2746;
assign a2922 = a2920 & a2918;
assign a2924 = ~l934 & ~l932;
assign a2926 = l944 & l942;
assign a2928 = a2926 & a2756;
assign a2930 = a2928 & a2924;
assign a2932 = a2908 & a2756;
assign a2934 = a2932 & a2918;
assign a2936 = ~a2766 & l936;
assign a2938 = a2936 & ~a2934;
assign a2940 = a2938 & ~a2930;
assign a2942 = ~a2940 & ~a2922;
assign a2944 = ~a2942 & ~a2916;
assign a2946 = ~a2944 & ~a2914;
assign a2948 = ~a2946 & ~a2910;
assign a2952 = ~a2766 & l938;
assign a2954 = a2952 & ~a2934;
assign a2956 = a2954 & ~a2930;
assign a2958 = ~a2956 & ~a2922;
assign a2960 = ~a2958 & ~a2916;
assign a2962 = ~a2960 & ~a2914;
assign a2964 = a2962 & ~a2910;
assign a2968 = ~l934 & l932;
assign a2970 = a2912 & a2804;
assign a2972 = a2970 & a2968;
assign a2974 = a2912 & a2812;
assign a2976 = a2974 & a2924;
assign a2978 = a2968 & a2920;
assign a2980 = ~a2978 & ~l944;
assign a2982 = a2980 & ~a2976;
assign a2984 = a2982 & ~a2972;
assign a2988 = l958 & ~l956;
assign a2990 = a2988 & a2730;
assign a2992 = ~l958 & l956;
assign a2994 = a2992 & a2730;
assign a2996 = a2992 & a2740;
assign a2998 = l948 & ~l946;
assign a3000 = a2992 & a2746;
assign a3002 = a3000 & a2998;
assign a3004 = ~l948 & ~l946;
assign a3006 = l958 & l956;
assign a3008 = a3006 & a2756;
assign a3010 = a3008 & a3004;
assign a3012 = a2988 & a2756;
assign a3014 = a3012 & a2998;
assign a3016 = ~a2766 & l950;
assign a3018 = a3016 & ~a3014;
assign a3020 = a3018 & ~a3010;
assign a3022 = ~a3020 & ~a3002;
assign a3024 = ~a3022 & ~a2996;
assign a3026 = ~a3024 & ~a2994;
assign a3028 = ~a3026 & ~a2990;
assign a3032 = ~a2766 & l952;
assign a3034 = a3032 & ~a3014;
assign a3036 = a3034 & ~a3010;
assign a3038 = ~a3036 & ~a3002;
assign a3040 = ~a3038 & ~a2996;
assign a3042 = ~a3040 & ~a2994;
assign a3044 = a3042 & ~a2990;
assign a3048 = ~l948 & l946;
assign a3050 = a2992 & a2804;
assign a3052 = a3050 & a3048;
assign a3054 = a2992 & a2812;
assign a3056 = a3054 & a3004;
assign a3058 = a3048 & a3000;
assign a3060 = ~a3058 & ~l958;
assign a3062 = a3060 & ~a3056;
assign a3064 = a3062 & ~a3052;
assign a3068 = ~l978 & l972;
assign a3070 = ~a2832 & ~a2734;
assign a3072 = a3070 & ~a2912;
assign a3074 = a2832 & a2734;
assign a3076 = ~a3074 & ~a2912;
assign a3078 = ~a3076 & ~a3070;
assign a3080 = ~a3078 & ~a2992;
assign a3082 = ~a3080 & ~a3072;
assign a3084 = ~a3082 & a2804;
assign a3086 = a3084 & ~a3068;
assign a3088 = ~a2744 & a2726;
assign a3090 = ~a3088 & a2730;
assign a3092 = ~a2838 & a2828;
assign a3094 = ~a3092 & a3090;
assign a3096 = ~a2918 & a2908;
assign a3098 = ~a3096 & a3094;
assign a3100 = ~a2998 & a2988;
assign a3102 = ~a3100 & a3098;
assign a3104 = ~a2752 & a2734;
assign a3106 = ~a3104 & a2812;
assign a3108 = ~a2844 & a2832;
assign a3110 = ~a3108 & a3106;
assign a3112 = ~a2924 & a2912;
assign a3114 = ~a3112 & a3110;
assign a3116 = ~a3004 & a2992;
assign a3118 = ~a3116 & a3114;
assign a3120 = ~a3048 & a2992;
assign a3122 = ~a2968 & a2912;
assign a3124 = ~a2888 & a2832;
assign a3126 = ~a2800 & a2734;
assign a3128 = ~a3126 & a2812;
assign a3130 = a3128 & ~a3124;
assign a3132 = a3130 & ~a3122;
assign a3134 = a3132 & ~a3120;
assign a3136 = ~a2998 & a2992;
assign a3138 = ~a2918 & a2912;
assign a3140 = ~a2744 & a2734;
assign a3142 = ~a2838 & a2832;
assign a3144 = ~a3142 & ~a3140;
assign a3146 = a3144 & ~a3138;
assign a3148 = a3146 & ~a3136;
assign a3150 = ~a3126 & ~a3124;
assign a3152 = a3150 & ~a3122;
assign a3154 = a3152 & ~a3120;
assign a3156 = ~a3154 & ~a3148;
assign a3158 = ~a3156 & ~a2738;
assign a3160 = a3158 & a2746;
assign a3162 = a3160 & ~a2802;
assign a3164 = ~a3162 & l960;
assign a3166 = ~a3164 & ~a3134;
assign a3168 = ~a3166 & ~a3118;
assign a3170 = a3168 & ~a3102;
assign a3172 = a3170 & ~a3086;
assign a3176 = a2740 & ~l974;
assign a3178 = a2802 & l960;
assign a3180 = l964 & l960;
assign a3182 = a3180 & l974;
assign a3184 = ~a3182 & a3178;
assign a3186 = ~a3184 & ~l962;
assign a3188 = a3186 & ~a3176;
assign a3190 = ~a3188 & ~a3134;
assign a3192 = a3190 & ~a3118;
assign a3194 = ~a3192 & ~a3102;
assign a3196 = a3194 & ~a3086;
assign a3200 = a2740 & l974;
assign a3202 = ~a3138 & ~a3136;
assign a3204 = a3202 & ~a3142;
assign a3206 = a3204 & ~a3140;
assign a3208 = a3206 & a2746;
assign a3210 = ~a3208 & l964;
assign a3212 = ~a3210 & ~a3178;
assign a3214 = ~a3212 & ~a3200;
assign a3216 = ~a3214 & ~a3176;
assign a3218 = a3216 & ~a3134;
assign a3220 = a3218 & ~a3118;
assign a3222 = ~a3220 & ~a3102;
assign a3224 = ~a3222 & ~a3086;
assign a3228 = ~l984 & ~l982;
assign a3230 = ~a3228 & l980;
assign a3232 = a3230 & l978;
assign a3234 = a3232 & a2804;
assign a3236 = ~a3234 & ~l976;
assign a3240 = ~l982 & ~l980;
assign a3242 = a3240 & ~l978;
assign a3244 = l984 & ~l982;
assign a3246 = a3244 & ~l980;
assign a3248 = a3246 & ~l978;
assign a3250 = l982 & ~l980;
assign a3252 = a3250 & ~l978;
assign a3254 = l984 & l982;
assign a3256 = a3254 & ~l980;
assign a3258 = a3256 & ~l978;
assign a3260 = ~l982 & l980;
assign a3262 = a3260 & ~l978;
assign a3264 = a3244 & l980;
assign a3266 = a3264 & ~l978;
assign a3268 = l982 & l980;
assign a3270 = a3268 & ~l978;
assign a3272 = a3246 & l978;
assign a3274 = a3256 & l978;
assign a3276 = ~a3274 & a3260;
assign a3278 = ~a3276 & ~a3250;
assign a3280 = ~a3278 & ~a3272;
assign a3282 = ~a3280 & ~a3240;
assign a3284 = ~a3282 & l978;
assign a3286 = ~a3284 & ~a3270;
assign a3288 = ~a3286 & ~a3266;
assign a3290 = ~a3288 & ~a3262;
assign a3292 = ~a3290 & ~a3258;
assign a3294 = ~a3292 & ~a3252;
assign a3296 = ~a3294 & ~a3248;
assign a3298 = ~a3296 & ~a3242;
assign a3300 = ~a3298 & ~l984;
assign a3302 = a3228 & ~l980;
assign a3304 = a3302 & ~l978;
assign a3306 = l984 & ~l980;
assign a3308 = a3306 & ~l978;
assign a3310 = a3228 & l980;
assign a3312 = a3310 & ~l978;
assign a3314 = l984 & l980;
assign a3316 = a3314 & ~l978;
assign a3318 = a3302 & l978;
assign a3320 = ~l980 & l978;
assign a3322 = a3320 & ~a3244;
assign a3324 = a3322 & ~a3318;
assign a3326 = ~a3324 & ~a3316;
assign a3328 = ~l984 & l980;
assign a3330 = a3328 & ~l978;
assign a3332 = ~a3330 & a3326;
assign a3334 = ~a3332 & ~a3266;
assign a3336 = a3334 & ~a3312;
assign a3338 = ~a3336 & ~a3308;
assign a3340 = ~l984 & ~l980;
assign a3342 = a3340 & ~l978;
assign a3344 = ~a3342 & a3338;
assign a3346 = ~a3344 & l982;
assign a3348 = a3346 & ~a3248;
assign a3350 = a3348 & ~a3304;
assign a3352 = a3350 & a3300;
assign a3354 = ~l984 & l982;
assign a3356 = ~a3254 & ~l978;
assign a3358 = a3356 & ~a3354;
assign a3360 = a3244 & ~l978;
assign a3362 = ~a3360 & a3358;
assign a3364 = a3228 & ~l978;
assign a3366 = ~a3364 & a3362;
assign a3368 = ~a3366 & ~l980;
assign a3370 = ~a3368 & a3352;
assign a3372 = ~a3254 & ~l980;
assign a3374 = a3372 & ~a3354;
assign a3376 = a3374 & ~a3246;
assign a3378 = a3376 & ~a3302;
assign a3380 = ~a3378 & ~l978;
assign a3382 = ~a3380 & a3370;
assign a3384 = ~a3382 & l978;
assign a3386 = ~a3384 & a2804;
assign a3388 = ~a2804 & ~l978;
assign a3390 = ~a3388 & ~a3386;
assign a3394 = ~a3382 & l980;
assign a3396 = ~a3394 & a2804;
assign a3398 = ~a2804 & ~l980;
assign a3400 = ~a3398 & ~a3396;
assign a3404 = ~a3382 & l982;
assign a3406 = ~a3404 & a2804;
assign a3408 = ~a2804 & ~l982;
assign a3410 = ~a3408 & ~a3406;
assign a3414 = ~a3382 & ~l984;
assign a3416 = ~a3414 & a2804;
assign a3418 = ~a2804 & ~l984;
assign a3420 = ~a3418 & ~a3416;
assign a3424 = l998 & ~l996;
assign a3426 = l1046 & l1044;
assign a3428 = a3426 & ~l1042;
assign a3430 = a3428 & a3424;
assign a3432 = ~l998 & l996;
assign a3434 = a3432 & a3428;
assign a3436 = l1046 & ~l1044;
assign a3438 = a3436 & l1042;
assign a3440 = a3438 & a3432;
assign a3442 = l988 & ~l986;
assign a3444 = a3426 & l1042;
assign a3446 = a3444 & a3432;
assign a3448 = a3446 & a3442;
assign a3450 = ~l988 & ~l986;
assign a3452 = l998 & l996;
assign a3454 = a3436 & ~l1042;
assign a3456 = a3454 & a3452;
assign a3458 = a3456 & a3450;
assign a3460 = a3454 & a3424;
assign a3462 = a3460 & a3442;
assign a3464 = a3454 & l1048;
assign a3466 = ~a3464 & l990;
assign a3468 = a3466 & ~a3462;
assign a3470 = a3468 & ~a3458;
assign a3472 = ~a3470 & ~a3448;
assign a3474 = ~a3472 & ~a3440;
assign a3476 = ~a3474 & ~a3434;
assign a3478 = ~a3476 & ~a3430;
assign a3482 = ~a3464 & l992;
assign a3484 = a3482 & ~a3462;
assign a3486 = a3484 & ~a3458;
assign a3488 = ~a3486 & ~a3448;
assign a3490 = ~a3488 & ~a3440;
assign a3492 = ~a3490 & ~a3434;
assign a3494 = a3492 & ~a3430;
assign a3498 = ~l988 & l986;
assign a3500 = ~l1046 & ~l1044;
assign a3502 = a3500 & ~l1042;
assign a3504 = a3502 & a3432;
assign a3506 = a3504 & a3498;
assign a3508 = ~l1046 & l1044;
assign a3510 = a3508 & ~l1042;
assign a3512 = a3510 & a3432;
assign a3514 = a3512 & a3450;
assign a3516 = a3498 & a3446;
assign a3518 = ~a3516 & ~l998;
assign a3520 = a3518 & ~a3514;
assign a3522 = a3520 & ~a3506;
assign a3526 = l1012 & ~l1010;
assign a3528 = a3526 & a3428;
assign a3530 = ~l1012 & l1010;
assign a3532 = a3530 & a3428;
assign a3534 = a3530 & a3438;
assign a3536 = l1002 & ~l1000;
assign a3538 = a3530 & a3444;
assign a3540 = a3538 & a3536;
assign a3542 = ~l1002 & ~l1000;
assign a3544 = l1012 & l1010;
assign a3546 = a3544 & a3454;
assign a3548 = a3546 & a3542;
assign a3550 = a3526 & a3454;
assign a3552 = a3550 & a3536;
assign a3554 = ~a3464 & l1004;
assign a3556 = a3554 & ~a3552;
assign a3558 = a3556 & ~a3548;
assign a3560 = ~a3558 & ~a3540;
assign a3562 = ~a3560 & ~a3534;
assign a3564 = ~a3562 & ~a3532;
assign a3566 = ~a3564 & ~a3528;
assign a3570 = ~a3464 & l1006;
assign a3572 = a3570 & ~a3552;
assign a3574 = a3572 & ~a3548;
assign a3576 = ~a3574 & ~a3540;
assign a3578 = ~a3576 & ~a3534;
assign a3580 = ~a3578 & ~a3532;
assign a3582 = a3580 & ~a3528;
assign a3586 = ~l1002 & l1000;
assign a3588 = a3530 & a3502;
assign a3590 = a3588 & a3586;
assign a3592 = a3530 & a3510;
assign a3594 = a3592 & a3542;
assign a3596 = a3586 & a3538;
assign a3598 = ~a3596 & ~l1012;
assign a3600 = a3598 & ~a3594;
assign a3602 = a3600 & ~a3590;
assign a3606 = l1026 & ~l1024;
assign a3608 = a3606 & a3428;
assign a3610 = ~l1026 & l1024;
assign a3612 = a3610 & a3428;
assign a3614 = a3610 & a3438;
assign a3616 = l1016 & ~l1014;
assign a3618 = a3610 & a3444;
assign a3620 = a3618 & a3616;
assign a3622 = ~l1016 & ~l1014;
assign a3624 = l1026 & l1024;
assign a3626 = a3624 & a3454;
assign a3628 = a3626 & a3622;
assign a3630 = a3606 & a3454;
assign a3632 = a3630 & a3616;
assign a3634 = ~a3464 & l1018;
assign a3636 = a3634 & ~a3632;
assign a3638 = a3636 & ~a3628;
assign a3640 = ~a3638 & ~a3620;
assign a3642 = ~a3640 & ~a3614;
assign a3644 = ~a3642 & ~a3612;
assign a3646 = ~a3644 & ~a3608;
assign a3650 = ~a3464 & l1020;
assign a3652 = a3650 & ~a3632;
assign a3654 = a3652 & ~a3628;
assign a3656 = ~a3654 & ~a3620;
assign a3658 = ~a3656 & ~a3614;
assign a3660 = ~a3658 & ~a3612;
assign a3662 = a3660 & ~a3608;
assign a3666 = ~l1016 & l1014;
assign a3668 = a3610 & a3502;
assign a3670 = a3668 & a3666;
assign a3672 = a3610 & a3510;
assign a3674 = a3672 & a3622;
assign a3676 = a3666 & a3618;
assign a3678 = ~a3676 & ~l1026;
assign a3680 = a3678 & ~a3674;
assign a3682 = a3680 & ~a3670;
assign a3686 = l1040 & ~l1038;
assign a3688 = a3686 & a3428;
assign a3690 = ~l1040 & l1038;
assign a3692 = a3690 & a3428;
assign a3694 = a3690 & a3438;
assign a3696 = l1030 & ~l1028;
assign a3698 = a3690 & a3444;
assign a3700 = a3698 & a3696;
assign a3702 = ~l1030 & ~l1028;
assign a3704 = l1040 & l1038;
assign a3706 = a3704 & a3454;
assign a3708 = a3706 & a3702;
assign a3710 = a3686 & a3454;
assign a3712 = a3710 & a3696;
assign a3714 = ~a3464 & l1032;
assign a3716 = a3714 & ~a3712;
assign a3718 = a3716 & ~a3708;
assign a3720 = ~a3718 & ~a3700;
assign a3722 = ~a3720 & ~a3694;
assign a3724 = ~a3722 & ~a3692;
assign a3726 = ~a3724 & ~a3688;
assign a3730 = ~a3464 & l1034;
assign a3732 = a3730 & ~a3712;
assign a3734 = a3732 & ~a3708;
assign a3736 = ~a3734 & ~a3700;
assign a3738 = ~a3736 & ~a3694;
assign a3740 = ~a3738 & ~a3692;
assign a3742 = a3740 & ~a3688;
assign a3746 = ~l1030 & l1028;
assign a3748 = a3690 & a3502;
assign a3750 = a3748 & a3746;
assign a3752 = a3690 & a3510;
assign a3754 = a3752 & a3702;
assign a3756 = a3746 & a3698;
assign a3758 = ~a3756 & ~l1040;
assign a3760 = a3758 & ~a3754;
assign a3762 = a3760 & ~a3750;
assign a3766 = ~l1060 & l1054;
assign a3768 = ~a3530 & ~a3432;
assign a3770 = a3768 & ~a3610;
assign a3772 = a3530 & a3432;
assign a3774 = ~a3772 & ~a3610;
assign a3776 = ~a3774 & ~a3768;
assign a3778 = ~a3776 & ~a3690;
assign a3780 = ~a3778 & ~a3770;
assign a3782 = ~a3780 & a3502;
assign a3784 = a3782 & ~a3766;
assign a3786 = ~a3442 & a3424;
assign a3788 = ~a3786 & a3428;
assign a3790 = ~a3536 & a3526;
assign a3792 = ~a3790 & a3788;
assign a3794 = ~a3616 & a3606;
assign a3796 = ~a3794 & a3792;
assign a3798 = ~a3696 & a3686;
assign a3800 = ~a3798 & a3796;
assign a3802 = ~a3450 & a3432;
assign a3804 = ~a3802 & a3510;
assign a3806 = ~a3542 & a3530;
assign a3808 = ~a3806 & a3804;
assign a3810 = ~a3622 & a3610;
assign a3812 = ~a3810 & a3808;
assign a3814 = ~a3702 & a3690;
assign a3816 = ~a3814 & a3812;
assign a3818 = ~a3746 & a3690;
assign a3820 = ~a3666 & a3610;
assign a3822 = ~a3586 & a3530;
assign a3824 = ~a3498 & a3432;
assign a3826 = ~a3824 & a3510;
assign a3828 = a3826 & ~a3822;
assign a3830 = a3828 & ~a3820;
assign a3832 = a3830 & ~a3818;
assign a3834 = ~a3696 & a3690;
assign a3836 = ~a3616 & a3610;
assign a3838 = ~a3442 & a3432;
assign a3840 = ~a3536 & a3530;
assign a3842 = ~a3840 & ~a3838;
assign a3844 = a3842 & ~a3836;
assign a3846 = a3844 & ~a3834;
assign a3848 = ~a3824 & ~a3822;
assign a3850 = a3848 & ~a3820;
assign a3852 = a3850 & ~a3818;
assign a3854 = ~a3852 & ~a3846;
assign a3856 = ~a3854 & ~a3436;
assign a3858 = a3856 & a3444;
assign a3860 = a3858 & ~a3500;
assign a3862 = ~a3860 & l1042;
assign a3864 = ~a3862 & ~a3832;
assign a3866 = ~a3864 & ~a3816;
assign a3868 = a3866 & ~a3800;
assign a3870 = a3868 & ~a3784;
assign a3874 = a3438 & ~l1056;
assign a3876 = a3500 & l1042;
assign a3878 = l1046 & l1042;
assign a3880 = a3878 & l1056;
assign a3882 = ~a3880 & a3876;
assign a3884 = ~a3882 & ~l1044;
assign a3886 = a3884 & ~a3874;
assign a3888 = ~a3886 & ~a3832;
assign a3890 = a3888 & ~a3816;
assign a3892 = ~a3890 & ~a3800;
assign a3894 = a3892 & ~a3784;
assign a3898 = a3438 & l1056;
assign a3900 = ~a3836 & ~a3834;
assign a3902 = a3900 & ~a3840;
assign a3904 = a3902 & ~a3838;
assign a3906 = a3904 & a3444;
assign a3908 = ~a3906 & l1046;
assign a3910 = ~a3908 & ~a3876;
assign a3912 = ~a3910 & ~a3898;
assign a3914 = ~a3912 & ~a3874;
assign a3916 = a3914 & ~a3832;
assign a3918 = a3916 & ~a3816;
assign a3920 = ~a3918 & ~a3800;
assign a3922 = ~a3920 & ~a3784;
assign a3926 = ~l1066 & ~l1064;
assign a3928 = ~a3926 & l1062;
assign a3930 = a3928 & l1060;
assign a3932 = a3930 & a3502;
assign a3934 = ~a3932 & ~l1058;
assign a3938 = ~l1064 & ~l1062;
assign a3940 = a3938 & ~l1060;
assign a3942 = l1066 & ~l1064;
assign a3944 = a3942 & ~l1062;
assign a3946 = a3944 & ~l1060;
assign a3948 = l1064 & ~l1062;
assign a3950 = a3948 & ~l1060;
assign a3952 = l1066 & l1064;
assign a3954 = a3952 & ~l1062;
assign a3956 = a3954 & ~l1060;
assign a3958 = ~l1064 & l1062;
assign a3960 = a3958 & ~l1060;
assign a3962 = a3942 & l1062;
assign a3964 = a3962 & ~l1060;
assign a3966 = l1064 & l1062;
assign a3968 = a3966 & ~l1060;
assign a3970 = a3944 & l1060;
assign a3972 = a3954 & l1060;
assign a3974 = ~a3972 & a3958;
assign a3976 = ~a3974 & ~a3948;
assign a3978 = ~a3976 & ~a3970;
assign a3980 = ~a3978 & ~a3938;
assign a3982 = ~a3980 & l1060;
assign a3984 = ~a3982 & ~a3968;
assign a3986 = ~a3984 & ~a3964;
assign a3988 = ~a3986 & ~a3960;
assign a3990 = ~a3988 & ~a3956;
assign a3992 = ~a3990 & ~a3950;
assign a3994 = ~a3992 & ~a3946;
assign a3996 = ~a3994 & ~a3940;
assign a3998 = ~a3996 & ~l1066;
assign a4000 = a3926 & ~l1062;
assign a4002 = a4000 & ~l1060;
assign a4004 = l1066 & ~l1062;
assign a4006 = a4004 & ~l1060;
assign a4008 = a3926 & l1062;
assign a4010 = a4008 & ~l1060;
assign a4012 = l1066 & l1062;
assign a4014 = a4012 & ~l1060;
assign a4016 = a4000 & l1060;
assign a4018 = ~l1062 & l1060;
assign a4020 = a4018 & ~a3942;
assign a4022 = a4020 & ~a4016;
assign a4024 = ~a4022 & ~a4014;
assign a4026 = ~l1066 & l1062;
assign a4028 = a4026 & ~l1060;
assign a4030 = ~a4028 & a4024;
assign a4032 = ~a4030 & ~a3964;
assign a4034 = a4032 & ~a4010;
assign a4036 = ~a4034 & ~a4006;
assign a4038 = ~l1066 & ~l1062;
assign a4040 = a4038 & ~l1060;
assign a4042 = ~a4040 & a4036;
assign a4044 = ~a4042 & l1064;
assign a4046 = a4044 & ~a3946;
assign a4048 = a4046 & ~a4002;
assign a4050 = a4048 & a3998;
assign a4052 = ~l1066 & l1064;
assign a4054 = ~a3952 & ~l1060;
assign a4056 = a4054 & ~a4052;
assign a4058 = a3942 & ~l1060;
assign a4060 = ~a4058 & a4056;
assign a4062 = a3926 & ~l1060;
assign a4064 = ~a4062 & a4060;
assign a4066 = ~a4064 & ~l1062;
assign a4068 = ~a4066 & a4050;
assign a4070 = ~a3952 & ~l1062;
assign a4072 = a4070 & ~a4052;
assign a4074 = a4072 & ~a3944;
assign a4076 = a4074 & ~a4000;
assign a4078 = ~a4076 & ~l1060;
assign a4080 = ~a4078 & a4068;
assign a4082 = ~a4080 & l1060;
assign a4084 = ~a4082 & a3502;
assign a4086 = ~a3502 & ~l1060;
assign a4088 = ~a4086 & ~a4084;
assign a4092 = ~a4080 & l1062;
assign a4094 = ~a4092 & a3502;
assign a4096 = ~a3502 & ~l1062;
assign a4098 = ~a4096 & ~a4094;
assign a4102 = ~a4080 & l1064;
assign a4104 = ~a4102 & a3502;
assign a4106 = ~a3502 & ~l1064;
assign a4108 = ~a4106 & ~a4104;
assign a4112 = ~a4080 & ~l1066;
assign a4114 = ~a4112 & a3502;
assign a4116 = ~a3502 & ~l1066;
assign a4118 = ~a4116 & ~a4114;
assign a4122 = ~a2480 & l1070;
assign a4124 = ~a4122 & ~a1782;
assign a4128 = ~l1316 & ~l1314;
assign a4130 = ~a4128 & l1068;
assign a4132 = ~a4130 & ~l1308;
assign a4136 = ~l1072 & l884;
assign a4138 = ~a4136 & l1074;
assign a4140 = ~a4138 & ~a4128;
assign a4142 = ~a4140 & ~l1310;
assign a4146 = l1072 & l884;
assign a4148 = ~a4146 & ~a4128;
assign a4150 = ~a4148 & ~l1312;
assign a4156 = ~l1072 & ~l884;
assign a4158 = l1068 & ~i330;
assign a4160 = a4136 & ~l1074;
assign a4162 = ~a4160 & ~a4158;
assign a4164 = a4162 & ~a4156;
assign a4166 = l580 & ~i2;
assign a4168 = ~l580 & i2;
assign a4170 = ~a4168 & ~a4166;
assign a4172 = a4170 & a4164;
assign a4174 = l582 & ~i4;
assign a4176 = ~l582 & i4;
assign a4178 = ~a4176 & ~a4174;
assign a4180 = a4178 & a4172;
assign a4182 = l584 & ~i6;
assign a4184 = ~l584 & i6;
assign a4186 = ~a4184 & ~a4182;
assign a4188 = a4186 & a4180;
assign a4190 = l586 & ~i8;
assign a4192 = ~l586 & i8;
assign a4194 = ~a4192 & ~a4190;
assign a4196 = a4194 & a4188;
assign a4198 = l588 & ~i10;
assign a4200 = ~l588 & i10;
assign a4202 = ~a4200 & ~a4198;
assign a4204 = a4202 & a4196;
assign a4206 = l590 & ~i12;
assign a4208 = ~l590 & i12;
assign a4210 = ~a4208 & ~a4206;
assign a4212 = a4210 & a4204;
assign a4214 = l592 & ~i14;
assign a4216 = ~l592 & i14;
assign a4218 = ~a4216 & ~a4214;
assign a4220 = a4218 & a4212;
assign a4222 = l594 & ~i16;
assign a4224 = ~l594 & i16;
assign a4226 = ~a4224 & ~a4222;
assign a4228 = a4226 & a4220;
assign a4230 = l596 & ~i18;
assign a4232 = ~l596 & i18;
assign a4234 = ~a4232 & ~a4230;
assign a4236 = a4234 & a4228;
assign a4238 = l598 & ~i20;
assign a4240 = ~l598 & i20;
assign a4242 = ~a4240 & ~a4238;
assign a4244 = a4242 & a4236;
assign a4246 = l600 & ~i22;
assign a4248 = ~l600 & i22;
assign a4250 = ~a4248 & ~a4246;
assign a4252 = a4250 & a4244;
assign a4254 = l602 & ~i24;
assign a4256 = ~l602 & i24;
assign a4258 = ~a4256 & ~a4254;
assign a4260 = a4258 & a4252;
assign a4262 = l604 & ~i26;
assign a4264 = ~l604 & i26;
assign a4266 = ~a4264 & ~a4262;
assign a4268 = a4266 & a4260;
assign a4270 = l606 & ~i28;
assign a4272 = ~l606 & i28;
assign a4274 = ~a4272 & ~a4270;
assign a4276 = a4274 & a4268;
assign a4278 = l608 & ~i30;
assign a4280 = ~l608 & i30;
assign a4282 = ~a4280 & ~a4278;
assign a4284 = a4282 & a4276;
assign a4286 = l610 & ~i32;
assign a4288 = ~l610 & i32;
assign a4290 = ~a4288 & ~a4286;
assign a4292 = a4290 & a4284;
assign a4294 = l612 & ~i34;
assign a4296 = ~l612 & i34;
assign a4298 = ~a4296 & ~a4294;
assign a4300 = a4298 & a4292;
assign a4302 = l614 & ~i36;
assign a4304 = ~l614 & i36;
assign a4306 = ~a4304 & ~a4302;
assign a4308 = a4306 & a4300;
assign a4310 = l616 & ~i38;
assign a4312 = ~l616 & i38;
assign a4314 = ~a4312 & ~a4310;
assign a4316 = a4314 & a4308;
assign a4318 = l618 & ~i40;
assign a4320 = ~l618 & i40;
assign a4322 = ~a4320 & ~a4318;
assign a4324 = a4322 & a4316;
assign a4326 = l620 & ~i42;
assign a4328 = ~l620 & i42;
assign a4330 = ~a4328 & ~a4326;
assign a4332 = a4330 & a4324;
assign a4334 = l622 & ~i44;
assign a4336 = ~l622 & i44;
assign a4338 = ~a4336 & ~a4334;
assign a4340 = a4338 & a4332;
assign a4342 = l624 & ~i46;
assign a4344 = ~l624 & i46;
assign a4346 = ~a4344 & ~a4342;
assign a4348 = a4346 & a4340;
assign a4350 = l626 & ~i48;
assign a4352 = ~l626 & i48;
assign a4354 = ~a4352 & ~a4350;
assign a4356 = a4354 & a4348;
assign a4358 = l628 & ~i50;
assign a4360 = ~l628 & i50;
assign a4362 = ~a4360 & ~a4358;
assign a4364 = a4362 & a4356;
assign a4366 = l630 & ~i52;
assign a4368 = ~l630 & i52;
assign a4370 = ~a4368 & ~a4366;
assign a4372 = a4370 & a4364;
assign a4374 = l632 & ~i54;
assign a4376 = ~l632 & i54;
assign a4378 = ~a4376 & ~a4374;
assign a4380 = a4378 & a4372;
assign a4382 = l634 & ~i56;
assign a4384 = ~l634 & i56;
assign a4386 = ~a4384 & ~a4382;
assign a4388 = a4386 & a4380;
assign a4390 = l636 & ~i58;
assign a4392 = ~l636 & i58;
assign a4394 = ~a4392 & ~a4390;
assign a4396 = a4394 & a4388;
assign a4398 = l638 & ~i60;
assign a4400 = ~l638 & i60;
assign a4402 = ~a4400 & ~a4398;
assign a4404 = a4402 & a4396;
assign a4406 = l640 & ~i62;
assign a4408 = ~l640 & i62;
assign a4410 = ~a4408 & ~a4406;
assign a4412 = a4410 & a4404;
assign a4414 = l642 & ~i64;
assign a4416 = ~l642 & i64;
assign a4418 = ~a4416 & ~a4414;
assign a4420 = a4418 & a4412;
assign a4422 = l644 & ~i66;
assign a4424 = ~l644 & i66;
assign a4426 = ~a4424 & ~a4422;
assign a4428 = a4426 & a4420;
assign a4430 = l646 & ~i68;
assign a4432 = ~l646 & i68;
assign a4434 = ~a4432 & ~a4430;
assign a4436 = a4434 & a4428;
assign a4438 = l648 & ~i70;
assign a4440 = ~l648 & i70;
assign a4442 = ~a4440 & ~a4438;
assign a4444 = a4442 & a4436;
assign a4446 = l650 & ~i72;
assign a4448 = ~l650 & i72;
assign a4450 = ~a4448 & ~a4446;
assign a4452 = a4450 & a4444;
assign a4454 = l652 & ~i74;
assign a4456 = ~l652 & i74;
assign a4458 = ~a4456 & ~a4454;
assign a4460 = a4458 & a4452;
assign a4462 = l654 & ~i76;
assign a4464 = ~l654 & i76;
assign a4466 = ~a4464 & ~a4462;
assign a4468 = a4466 & a4460;
assign a4470 = l656 & ~i78;
assign a4472 = ~l656 & i78;
assign a4474 = ~a4472 & ~a4470;
assign a4476 = a4474 & a4468;
assign a4478 = l658 & ~i80;
assign a4480 = ~l658 & i80;
assign a4482 = ~a4480 & ~a4478;
assign a4484 = a4482 & a4476;
assign a4486 = l660 & ~i82;
assign a4488 = ~l660 & i82;
assign a4490 = ~a4488 & ~a4486;
assign a4492 = a4490 & a4484;
assign a4494 = l662 & ~i84;
assign a4496 = ~l662 & i84;
assign a4498 = ~a4496 & ~a4494;
assign a4500 = a4498 & a4492;
assign a4502 = l664 & ~i86;
assign a4504 = ~l664 & i86;
assign a4506 = ~a4504 & ~a4502;
assign a4508 = a4506 & a4500;
assign a4510 = l666 & ~i88;
assign a4512 = ~l666 & i88;
assign a4514 = ~a4512 & ~a4510;
assign a4516 = a4514 & a4508;
assign a4518 = l668 & ~i90;
assign a4520 = ~l668 & i90;
assign a4522 = ~a4520 & ~a4518;
assign a4524 = a4522 & a4516;
assign a4526 = l670 & ~i92;
assign a4528 = ~l670 & i92;
assign a4530 = ~a4528 & ~a4526;
assign a4532 = a4530 & a4524;
assign a4534 = l672 & ~i94;
assign a4536 = ~l672 & i94;
assign a4538 = ~a4536 & ~a4534;
assign a4540 = a4538 & a4532;
assign a4542 = l674 & ~i96;
assign a4544 = ~l674 & i96;
assign a4546 = ~a4544 & ~a4542;
assign a4548 = a4546 & a4540;
assign a4550 = l676 & ~i98;
assign a4552 = ~l676 & i98;
assign a4554 = ~a4552 & ~a4550;
assign a4556 = a4554 & a4548;
assign a4558 = l678 & ~i100;
assign a4560 = ~l678 & i100;
assign a4562 = ~a4560 & ~a4558;
assign a4564 = a4562 & a4556;
assign a4566 = l680 & ~i102;
assign a4568 = ~l680 & i102;
assign a4570 = ~a4568 & ~a4566;
assign a4572 = a4570 & a4564;
assign a4574 = l682 & ~i104;
assign a4576 = ~l682 & i104;
assign a4578 = ~a4576 & ~a4574;
assign a4580 = a4578 & a4572;
assign a4582 = l684 & ~i106;
assign a4584 = ~l684 & i106;
assign a4586 = ~a4584 & ~a4582;
assign a4588 = a4586 & a4580;
assign a4590 = l686 & ~i108;
assign a4592 = ~l686 & i108;
assign a4594 = ~a4592 & ~a4590;
assign a4596 = a4594 & a4588;
assign a4598 = l688 & ~i110;
assign a4600 = ~l688 & i110;
assign a4602 = ~a4600 & ~a4598;
assign a4604 = a4602 & a4596;
assign a4606 = l690 & ~i112;
assign a4608 = ~l690 & i112;
assign a4610 = ~a4608 & ~a4606;
assign a4612 = a4610 & a4604;
assign a4614 = l692 & ~i114;
assign a4616 = ~l692 & i114;
assign a4618 = ~a4616 & ~a4614;
assign a4620 = a4618 & a4612;
assign a4622 = l694 & ~i116;
assign a4624 = ~l694 & i116;
assign a4626 = ~a4624 & ~a4622;
assign a4628 = a4626 & a4620;
assign a4630 = l696 & ~i118;
assign a4632 = ~l696 & i118;
assign a4634 = ~a4632 & ~a4630;
assign a4636 = a4634 & a4628;
assign a4638 = l698 & ~i120;
assign a4640 = ~l698 & i120;
assign a4642 = ~a4640 & ~a4638;
assign a4644 = a4642 & a4636;
assign a4646 = l700 & ~i122;
assign a4648 = ~l700 & i122;
assign a4650 = ~a4648 & ~a4646;
assign a4652 = a4650 & a4644;
assign a4654 = l702 & ~i124;
assign a4656 = ~l702 & i124;
assign a4658 = ~a4656 & ~a4654;
assign a4660 = a4658 & a4652;
assign a4662 = l704 & ~i126;
assign a4664 = ~l704 & i126;
assign a4666 = ~a4664 & ~a4662;
assign a4668 = a4666 & a4660;
assign a4670 = l706 & ~i128;
assign a4672 = ~l706 & i128;
assign a4674 = ~a4672 & ~a4670;
assign a4676 = a4674 & a4668;
assign a4678 = l708 & ~i130;
assign a4680 = ~l708 & i130;
assign a4682 = ~a4680 & ~a4678;
assign a4684 = a4682 & a4676;
assign a4686 = l710 & ~i132;
assign a4688 = ~l710 & i132;
assign a4690 = ~a4688 & ~a4686;
assign a4692 = a4690 & a4684;
assign a4694 = l712 & ~i134;
assign a4696 = ~l712 & i134;
assign a4698 = ~a4696 & ~a4694;
assign a4700 = a4698 & a4692;
assign a4702 = l714 & ~i136;
assign a4704 = ~l714 & i136;
assign a4706 = ~a4704 & ~a4702;
assign a4708 = a4706 & a4700;
assign a4710 = l716 & ~i138;
assign a4712 = ~l716 & i138;
assign a4714 = ~a4712 & ~a4710;
assign a4716 = a4714 & a4708;
assign a4718 = l718 & ~i140;
assign a4720 = ~l718 & i140;
assign a4722 = ~a4720 & ~a4718;
assign a4724 = a4722 & a4716;
assign a4726 = l720 & ~i142;
assign a4728 = ~l720 & i142;
assign a4730 = ~a4728 & ~a4726;
assign a4732 = a4730 & a4724;
assign a4734 = l722 & ~i144;
assign a4736 = ~l722 & i144;
assign a4738 = ~a4736 & ~a4734;
assign a4740 = a4738 & a4732;
assign a4742 = l724 & ~i146;
assign a4744 = ~l724 & i146;
assign a4746 = ~a4744 & ~a4742;
assign a4748 = a4746 & a4740;
assign a4750 = l726 & ~i148;
assign a4752 = ~l726 & i148;
assign a4754 = ~a4752 & ~a4750;
assign a4756 = a4754 & a4748;
assign a4758 = l728 & ~i150;
assign a4760 = ~l728 & i150;
assign a4762 = ~a4760 & ~a4758;
assign a4764 = a4762 & a4756;
assign a4766 = l730 & ~i152;
assign a4768 = ~l730 & i152;
assign a4770 = ~a4768 & ~a4766;
assign a4772 = a4770 & a4764;
assign a4774 = l732 & ~i154;
assign a4776 = ~l732 & i154;
assign a4778 = ~a4776 & ~a4774;
assign a4780 = a4778 & a4772;
assign a4782 = l734 & ~i156;
assign a4784 = ~l734 & i156;
assign a4786 = ~a4784 & ~a4782;
assign a4788 = a4786 & a4780;
assign a4790 = l736 & ~i158;
assign a4792 = ~l736 & i158;
assign a4794 = ~a4792 & ~a4790;
assign a4796 = a4794 & a4788;
assign a4798 = l738 & ~i160;
assign a4800 = ~l738 & i160;
assign a4802 = ~a4800 & ~a4798;
assign a4804 = a4802 & a4796;
assign a4806 = l748 & ~i166;
assign a4808 = ~l748 & i166;
assign a4810 = ~a4808 & ~a4806;
assign a4812 = a4810 & a4804;
assign a4814 = a1416 & ~l752;
assign a4816 = a4814 & a1356;
assign a4818 = ~a4816 & a1422;
assign a4820 = ~a4818 & l750;
assign a4822 = a4820 & ~a1412;
assign a4824 = a4822 & ~i168;
assign a4826 = ~a4822 & i168;
assign a4828 = ~a4826 & ~a4824;
assign a4830 = a4828 & a4812;
assign a4832 = l762 & ~i174;
assign a4834 = ~l762 & i174;
assign a4836 = ~a4834 & ~a4832;
assign a4838 = a4836 & a4830;
assign a4840 = a1416 & ~l766;
assign a4842 = a4840 & a1448;
assign a4844 = ~a4842 & a1502;
assign a4846 = ~a4844 & l764;
assign a4848 = a4846 & ~a1496;
assign a4850 = a4848 & ~i176;
assign a4852 = ~a4848 & i176;
assign a4854 = ~a4852 & ~a4850;
assign a4856 = a4854 & a4838;
assign a4858 = l776 & ~i182;
assign a4860 = ~l776 & i182;
assign a4862 = ~a4860 & ~a4858;
assign a4864 = a4862 & a4856;
assign a4866 = a1416 & ~l780;
assign a4868 = a4866 & a1528;
assign a4870 = ~a4868 & a1582;
assign a4872 = ~a4870 & l778;
assign a4874 = a4872 & ~a1576;
assign a4876 = a4874 & ~i184;
assign a4878 = ~a4874 & i184;
assign a4880 = ~a4878 & ~a4876;
assign a4882 = a4880 & a4864;
assign a4884 = l790 & ~i190;
assign a4886 = ~l790 & i190;
assign a4888 = ~a4886 & ~a4884;
assign a4890 = a4888 & a4882;
assign a4892 = a1416 & ~l794;
assign a4894 = a4892 & a1608;
assign a4896 = ~a4894 & a1662;
assign a4898 = ~a4896 & l792;
assign a4900 = a4898 & ~a1656;
assign a4902 = a4900 & ~i192;
assign a4904 = ~a4900 & i192;
assign a4906 = ~a4904 & ~a4902;
assign a4908 = a4906 & a4890;
assign a4910 = a1676 & ~a1596;
assign a4912 = ~a4910 & a1334;
assign a4914 = ~a1334 & ~l802;
assign a4916 = ~a4914 & ~a4912;
assign a4918 = a4916 & ~i194;
assign a4920 = ~a4916 & i194;
assign a4922 = ~a4920 & ~a4918;
assign a4924 = a4922 & a4908;
assign a4926 = ~a1598 & ~l804;
assign a4928 = a4926 & ~a1518;
assign a4930 = ~a4928 & ~a1438;
assign a4932 = a4930 & ~a1340;
assign a4934 = a4932 & ~i196;
assign a4936 = ~a4932 & i196;
assign a4938 = ~a4936 & ~a4934;
assign a4940 = a4938 & a4924;
assign a4942 = ~a1598 & ~l806;
assign a4944 = ~a4942 & ~a1518;
assign a4946 = ~a4944 & ~a1438;
assign a4948 = ~a4946 & ~a1340;
assign a4950 = a4948 & ~i198;
assign a4952 = ~a4948 & i198;
assign a4954 = ~a4952 & ~a4950;
assign a4956 = a4954 & a4940;
assign a4958 = l808 & ~i200;
assign a4960 = ~l808 & i200;
assign a4962 = ~a4960 & ~a4958;
assign a4964 = a4962 & a4956;
assign a4966 = a1416 & l1318;
assign a4968 = ~a1416 & ~l810;
assign a4970 = ~a4968 & ~a4966;
assign a4972 = a4970 & ~i202;
assign a4974 = ~a4970 & i202;
assign a4976 = ~a4974 & ~a4972;
assign a4978 = a4976 & a4964;
assign a4980 = l830 & ~i208;
assign a4982 = ~l830 & i208;
assign a4984 = ~a4982 & ~a4980;
assign a4986 = a4984 & a4978;
assign a4988 = a2114 & ~l834;
assign a4990 = a4988 & a2054;
assign a4992 = ~a4990 & a2120;
assign a4994 = ~a4992 & l832;
assign a4996 = a4994 & ~a2110;
assign a4998 = a4996 & ~i210;
assign a5000 = ~a4996 & i210;
assign a5002 = ~a5000 & ~a4998;
assign a5004 = a5002 & a4986;
assign a5006 = l844 & ~i216;
assign a5008 = ~l844 & i216;
assign a5010 = ~a5008 & ~a5006;
assign a5012 = a5010 & a5004;
assign a5014 = a2114 & ~l848;
assign a5016 = a5014 & a2146;
assign a5018 = ~a5016 & a2200;
assign a5020 = ~a5018 & l846;
assign a5022 = a5020 & ~a2194;
assign a5024 = a5022 & ~i218;
assign a5026 = ~a5022 & i218;
assign a5028 = ~a5026 & ~a5024;
assign a5030 = a5028 & a5012;
assign a5032 = l858 & ~i224;
assign a5034 = ~l858 & i224;
assign a5036 = ~a5034 & ~a5032;
assign a5038 = a5036 & a5030;
assign a5040 = a2114 & ~l862;
assign a5042 = a5040 & a2226;
assign a5044 = ~a5042 & a2280;
assign a5046 = ~a5044 & l860;
assign a5048 = a5046 & ~a2274;
assign a5050 = a5048 & ~i226;
assign a5052 = ~a5048 & i226;
assign a5054 = ~a5052 & ~a5050;
assign a5056 = a5054 & a5038;
assign a5058 = l872 & ~i232;
assign a5060 = ~l872 & i232;
assign a5062 = ~a5060 & ~a5058;
assign a5064 = a5062 & a5056;
assign a5066 = a2114 & ~l876;
assign a5068 = a5066 & a2306;
assign a5070 = ~a5068 & a2360;
assign a5072 = ~a5070 & l874;
assign a5074 = a5072 & ~a2354;
assign a5076 = a5074 & ~i234;
assign a5078 = ~a5074 & i234;
assign a5080 = ~a5078 & ~a5076;
assign a5082 = a5080 & a5064;
assign a5084 = a2374 & ~a2294;
assign a5086 = ~a5084 & a2032;
assign a5088 = ~a2032 & ~l884;
assign a5090 = ~a5088 & ~a5086;
assign a5092 = a5090 & ~i236;
assign a5094 = ~a5090 & i236;
assign a5096 = ~a5094 & ~a5092;
assign a5098 = a5096 & a5082;
assign a5100 = ~a2296 & ~l886;
assign a5102 = a5100 & ~a2216;
assign a5104 = ~a5102 & ~a2136;
assign a5106 = a5104 & ~a2038;
assign a5108 = a5106 & ~i238;
assign a5110 = ~a5106 & i238;
assign a5112 = ~a5110 & ~a5108;
assign a5114 = a5112 & a5098;
assign a5116 = ~a2296 & ~l888;
assign a5118 = ~a5116 & ~a2216;
assign a5120 = ~a5118 & ~a2136;
assign a5122 = ~a5120 & ~a2038;
assign a5124 = a5122 & ~i240;
assign a5126 = ~a5122 & i240;
assign a5128 = ~a5126 & ~a5124;
assign a5130 = a5128 & a5114;
assign a5132 = l890 & ~i242;
assign a5134 = ~l890 & i242;
assign a5136 = ~a5134 & ~a5132;
assign a5138 = a5136 & a5130;
assign a5140 = a2114 & l1320;
assign a5142 = ~a2114 & ~l892;
assign a5144 = ~a5142 & ~a5140;
assign a5146 = a5144 & ~i244;
assign a5148 = ~a5144 & i244;
assign a5150 = ~a5148 & ~a5146;
assign a5152 = a5150 & a5138;
assign a5154 = l912 & ~i250;
assign a5156 = ~l912 & i250;
assign a5158 = ~a5156 & ~a5154;
assign a5160 = a5158 & a5152;
assign a5162 = a2812 & ~l916;
assign a5164 = a5162 & a2752;
assign a5166 = ~a5164 & a2818;
assign a5168 = ~a5166 & l914;
assign a5170 = a5168 & ~a2808;
assign a5172 = a5170 & ~i252;
assign a5174 = ~a5170 & i252;
assign a5176 = ~a5174 & ~a5172;
assign a5178 = a5176 & a5160;
assign a5180 = l926 & ~i258;
assign a5182 = ~l926 & i258;
assign a5184 = ~a5182 & ~a5180;
assign a5186 = a5184 & a5178;
assign a5188 = a2812 & ~l930;
assign a5190 = a5188 & a2844;
assign a5192 = ~a5190 & a2898;
assign a5194 = ~a5192 & l928;
assign a5196 = a5194 & ~a2892;
assign a5198 = a5196 & ~i260;
assign a5200 = ~a5196 & i260;
assign a5202 = ~a5200 & ~a5198;
assign a5204 = a5202 & a5186;
assign a5206 = l940 & ~i266;
assign a5208 = ~l940 & i266;
assign a5210 = ~a5208 & ~a5206;
assign a5212 = a5210 & a5204;
assign a5214 = a2812 & ~l944;
assign a5216 = a5214 & a2924;
assign a5218 = ~a5216 & a2978;
assign a5220 = ~a5218 & l942;
assign a5222 = a5220 & ~a2972;
assign a5224 = a5222 & ~i268;
assign a5226 = ~a5222 & i268;
assign a5228 = ~a5226 & ~a5224;
assign a5230 = a5228 & a5212;
assign a5232 = l954 & ~i274;
assign a5234 = ~l954 & i274;
assign a5236 = ~a5234 & ~a5232;
assign a5238 = a5236 & a5230;
assign a5240 = a2812 & ~l958;
assign a5242 = a5240 & a3004;
assign a5244 = ~a5242 & a3058;
assign a5246 = ~a5244 & l956;
assign a5248 = a5246 & ~a3052;
assign a5250 = a5248 & ~i276;
assign a5252 = ~a5248 & i276;
assign a5254 = ~a5252 & ~a5250;
assign a5256 = a5254 & a5238;
assign a5258 = a3072 & ~a2992;
assign a5260 = ~a5258 & a2730;
assign a5262 = ~a2730 & ~l966;
assign a5264 = ~a5262 & ~a5260;
assign a5266 = a5264 & ~i278;
assign a5268 = ~a5264 & i278;
assign a5270 = ~a5268 & ~a5266;
assign a5272 = a5270 & a5256;
assign a5274 = ~a2994 & ~l968;
assign a5276 = a5274 & ~a2914;
assign a5278 = ~a5276 & ~a2834;
assign a5280 = a5278 & ~a2736;
assign a5282 = a5280 & ~i280;
assign a5284 = ~a5280 & i280;
assign a5286 = ~a5284 & ~a5282;
assign a5288 = a5286 & a5272;
assign a5290 = ~a2994 & ~l970;
assign a5292 = ~a5290 & ~a2914;
assign a5294 = ~a5292 & ~a2834;
assign a5296 = ~a5294 & ~a2736;
assign a5298 = a5296 & ~i282;
assign a5300 = ~a5296 & i282;
assign a5302 = ~a5300 & ~a5298;
assign a5304 = a5302 & a5288;
assign a5306 = l972 & ~i284;
assign a5308 = ~l972 & i284;
assign a5310 = ~a5308 & ~a5306;
assign a5312 = a5310 & a5304;
assign a5314 = a2812 & l1322;
assign a5316 = ~a2812 & ~l974;
assign a5318 = ~a5316 & ~a5314;
assign a5320 = a5318 & ~i286;
assign a5322 = ~a5318 & i286;
assign a5324 = ~a5322 & ~a5320;
assign a5326 = a5324 & a5312;
assign a5328 = l994 & ~i292;
assign a5330 = ~l994 & i292;
assign a5332 = ~a5330 & ~a5328;
assign a5334 = a5332 & a5326;
assign a5336 = a3510 & ~l998;
assign a5338 = a5336 & a3450;
assign a5340 = ~a5338 & a3516;
assign a5342 = ~a5340 & l996;
assign a5344 = a5342 & ~a3506;
assign a5346 = a5344 & ~i294;
assign a5348 = ~a5344 & i294;
assign a5350 = ~a5348 & ~a5346;
assign a5352 = a5350 & a5334;
assign a5354 = l1008 & ~i300;
assign a5356 = ~l1008 & i300;
assign a5358 = ~a5356 & ~a5354;
assign a5360 = a5358 & a5352;
assign a5362 = a3510 & ~l1012;
assign a5364 = a5362 & a3542;
assign a5366 = ~a5364 & a3596;
assign a5368 = ~a5366 & l1010;
assign a5370 = a5368 & ~a3590;
assign a5372 = a5370 & ~i302;
assign a5374 = ~a5370 & i302;
assign a5376 = ~a5374 & ~a5372;
assign a5378 = a5376 & a5360;
assign a5380 = l1022 & ~i308;
assign a5382 = ~l1022 & i308;
assign a5384 = ~a5382 & ~a5380;
assign a5386 = a5384 & a5378;
assign a5388 = a3510 & ~l1026;
assign a5390 = a5388 & a3622;
assign a5392 = ~a5390 & a3676;
assign a5394 = ~a5392 & l1024;
assign a5396 = a5394 & ~a3670;
assign a5398 = a5396 & ~i310;
assign a5400 = ~a5396 & i310;
assign a5402 = ~a5400 & ~a5398;
assign a5404 = a5402 & a5386;
assign a5406 = l1036 & ~i316;
assign a5408 = ~l1036 & i316;
assign a5410 = ~a5408 & ~a5406;
assign a5412 = a5410 & a5404;
assign a5414 = a3510 & ~l1040;
assign a5416 = a5414 & a3702;
assign a5418 = ~a5416 & a3756;
assign a5420 = ~a5418 & l1038;
assign a5422 = a5420 & ~a3750;
assign a5424 = a5422 & ~i318;
assign a5426 = ~a5422 & i318;
assign a5428 = ~a5426 & ~a5424;
assign a5430 = a5428 & a5412;
assign a5432 = a3770 & ~a3690;
assign a5434 = ~a5432 & a3428;
assign a5436 = ~a3428 & ~l1048;
assign a5438 = ~a5436 & ~a5434;
assign a5440 = a5438 & ~i320;
assign a5442 = ~a5438 & i320;
assign a5444 = ~a5442 & ~a5440;
assign a5446 = a5444 & a5430;
assign a5448 = ~a3692 & ~l1050;
assign a5450 = a5448 & ~a3612;
assign a5452 = ~a5450 & ~a3532;
assign a5454 = a5452 & ~a3434;
assign a5456 = a5454 & ~i322;
assign a5458 = ~a5454 & i322;
assign a5460 = ~a5458 & ~a5456;
assign a5462 = a5460 & a5446;
assign a5464 = ~a3692 & ~l1052;
assign a5466 = ~a5464 & ~a3612;
assign a5468 = ~a5466 & ~a3532;
assign a5470 = ~a5468 & ~a3434;
assign a5472 = a5470 & ~i324;
assign a5474 = ~a5470 & i324;
assign a5476 = ~a5474 & ~a5472;
assign a5478 = a5476 & a5462;
assign a5480 = l1054 & ~i326;
assign a5482 = ~l1054 & i326;
assign a5484 = ~a5482 & ~a5480;
assign a5486 = a5484 & a5478;
assign a5488 = a3510 & l1324;
assign a5490 = ~a3510 & ~l1056;
assign a5492 = ~a5490 & ~a5488;
assign a5494 = a5492 & ~i328;
assign a5496 = ~a5492 & i328;
assign a5498 = ~a5496 & ~a5494;
assign a5500 = a5498 & a5486;
assign a5502 = ~l1316 & l1314;
assign a5504 = a5502 & ~l744;
assign a5506 = ~a5502 & ~l1076;
assign a5508 = ~a5506 & ~a5504;
assign a5510 = a5508 & ~i336;
assign a5512 = ~a5508 & i336;
assign a5514 = ~a5512 & ~a5510;
assign a5516 = a5514 & a5500;
assign a5518 = ~a5502 & ~l1078;
assign a5520 = a5502 & l746;
assign a5522 = ~a5520 & ~a5518;
assign a5524 = a5522 & ~i338;
assign a5526 = ~a5522 & i338;
assign a5528 = ~a5526 & ~a5524;
assign a5530 = a5528 & a5516;
assign a5532 = a5502 & ~l750;
assign a5534 = ~a5502 & ~l1080;
assign a5536 = ~a5534 & ~a5532;
assign a5538 = a5536 & ~i340;
assign a5540 = ~a5536 & i340;
assign a5542 = ~a5540 & ~a5538;
assign a5544 = a5542 & a5530;
assign a5546 = ~a5502 & ~l1082;
assign a5548 = a5502 & l752;
assign a5550 = ~a5548 & ~a5546;
assign a5552 = a5550 & ~i342;
assign a5554 = ~a5550 & i342;
assign a5556 = ~a5554 & ~a5552;
assign a5558 = a5556 & a5544;
assign a5560 = a5502 & ~l758;
assign a5562 = ~a5502 & ~l1084;
assign a5564 = ~a5562 & ~a5560;
assign a5566 = a5564 & ~i344;
assign a5568 = ~a5564 & i344;
assign a5570 = ~a5568 & ~a5566;
assign a5572 = a5570 & a5558;
assign a5574 = ~a5502 & ~l1086;
assign a5576 = a5502 & l760;
assign a5578 = ~a5576 & ~a5574;
assign a5580 = a5578 & ~i346;
assign a5582 = ~a5578 & i346;
assign a5584 = ~a5582 & ~a5580;
assign a5586 = a5584 & a5572;
assign a5588 = a5502 & ~l764;
assign a5590 = ~a5502 & ~l1088;
assign a5592 = ~a5590 & ~a5588;
assign a5594 = a5592 & ~i348;
assign a5596 = ~a5592 & i348;
assign a5598 = ~a5596 & ~a5594;
assign a5600 = a5598 & a5586;
assign a5602 = ~a5502 & ~l1090;
assign a5604 = a5502 & l766;
assign a5606 = ~a5604 & ~a5602;
assign a5608 = a5606 & ~i350;
assign a5610 = ~a5606 & i350;
assign a5612 = ~a5610 & ~a5608;
assign a5614 = a5612 & a5600;
assign a5616 = a5502 & ~l772;
assign a5618 = ~a5502 & ~l1092;
assign a5620 = ~a5618 & ~a5616;
assign a5622 = a5620 & ~i352;
assign a5624 = ~a5620 & i352;
assign a5626 = ~a5624 & ~a5622;
assign a5628 = a5626 & a5614;
assign a5630 = ~a5502 & ~l1094;
assign a5632 = a5502 & l774;
assign a5634 = ~a5632 & ~a5630;
assign a5636 = a5634 & ~i354;
assign a5638 = ~a5634 & i354;
assign a5640 = ~a5638 & ~a5636;
assign a5642 = a5640 & a5628;
assign a5644 = a5502 & ~l778;
assign a5646 = ~a5502 & ~l1096;
assign a5648 = ~a5646 & ~a5644;
assign a5650 = a5648 & ~i356;
assign a5652 = ~a5648 & i356;
assign a5654 = ~a5652 & ~a5650;
assign a5656 = a5654 & a5642;
assign a5658 = ~a5502 & ~l1098;
assign a5660 = a5502 & l780;
assign a5662 = ~a5660 & ~a5658;
assign a5664 = a5662 & ~i358;
assign a5666 = ~a5662 & i358;
assign a5668 = ~a5666 & ~a5664;
assign a5670 = a5668 & a5656;
assign a5672 = a5502 & ~l786;
assign a5674 = ~a5502 & ~l1100;
assign a5676 = ~a5674 & ~a5672;
assign a5678 = a5676 & ~i360;
assign a5680 = ~a5676 & i360;
assign a5682 = ~a5680 & ~a5678;
assign a5684 = a5682 & a5670;
assign a5686 = ~a5502 & ~l1102;
assign a5688 = a5502 & l788;
assign a5690 = ~a5688 & ~a5686;
assign a5692 = a5690 & ~i362;
assign a5694 = ~a5690 & i362;
assign a5696 = ~a5694 & ~a5692;
assign a5698 = a5696 & a5684;
assign a5700 = a5502 & ~l792;
assign a5702 = ~a5502 & ~l1104;
assign a5704 = ~a5702 & ~a5700;
assign a5706 = a5704 & ~i364;
assign a5708 = ~a5704 & i364;
assign a5710 = ~a5708 & ~a5706;
assign a5712 = a5710 & a5698;
assign a5714 = ~a5502 & ~l1106;
assign a5716 = a5502 & l794;
assign a5718 = ~a5716 & ~a5714;
assign a5720 = a5718 & ~i366;
assign a5722 = ~a5718 & i366;
assign a5724 = ~a5722 & ~a5720;
assign a5726 = a5724 & a5712;
assign a5728 = a5502 & ~l796;
assign a5730 = ~a5502 & ~l1108;
assign a5732 = ~a5730 & ~a5728;
assign a5734 = a5732 & ~i368;
assign a5736 = ~a5732 & i368;
assign a5738 = ~a5736 & ~a5734;
assign a5740 = a5738 & a5726;
assign a5742 = a5502 & ~l798;
assign a5744 = ~a5502 & ~l1110;
assign a5746 = ~a5744 & ~a5742;
assign a5748 = a5746 & ~i370;
assign a5750 = ~a5746 & i370;
assign a5752 = ~a5750 & ~a5748;
assign a5754 = a5752 & a5740;
assign a5756 = ~a5502 & ~l1112;
assign a5758 = a5502 & l800;
assign a5760 = ~a5758 & ~a5756;
assign a5762 = a5760 & ~i372;
assign a5764 = ~a5760 & i372;
assign a5766 = ~a5764 & ~a5762;
assign a5768 = a5766 & a5754;
assign a5770 = a5502 & ~l802;
assign a5772 = ~a5502 & ~l1114;
assign a5774 = ~a5772 & ~a5770;
assign a5776 = a5774 & ~i374;
assign a5778 = ~a5774 & i374;
assign a5780 = ~a5778 & ~a5776;
assign a5782 = a5780 & a5768;
assign a5784 = a5502 & ~l804;
assign a5786 = ~a5502 & ~l1116;
assign a5788 = ~a5786 & ~a5784;
assign a5790 = a5788 & ~i376;
assign a5792 = ~a5788 & i376;
assign a5794 = ~a5792 & ~a5790;
assign a5796 = a5794 & a5782;
assign a5798 = a5502 & ~l806;
assign a5800 = ~a5502 & ~l1118;
assign a5802 = ~a5800 & ~a5798;
assign a5804 = a5802 & ~i378;
assign a5806 = ~a5802 & i378;
assign a5808 = ~a5806 & ~a5804;
assign a5810 = a5808 & a5796;
assign a5812 = a5502 & ~l810;
assign a5814 = ~a5502 & ~l1120;
assign a5816 = ~a5814 & ~a5812;
assign a5818 = a5816 & ~i380;
assign a5820 = ~a5816 & i380;
assign a5822 = ~a5820 & ~a5818;
assign a5824 = a5822 & a5810;
assign a5826 = a5502 & ~l812;
assign a5828 = ~a5502 & ~l1122;
assign a5830 = ~a5828 & ~a5826;
assign a5832 = a5830 & ~i382;
assign a5834 = ~a5830 & i382;
assign a5836 = ~a5834 & ~a5832;
assign a5838 = a5836 & a5824;
assign a5840 = a5502 & ~l814;
assign a5842 = ~a5502 & ~l1124;
assign a5844 = ~a5842 & ~a5840;
assign a5846 = a5844 & ~i384;
assign a5848 = ~a5844 & i384;
assign a5850 = ~a5848 & ~a5846;
assign a5852 = a5850 & a5838;
assign a5854 = a5502 & ~l816;
assign a5856 = ~a5502 & ~l1126;
assign a5858 = ~a5856 & ~a5854;
assign a5860 = a5858 & ~i386;
assign a5862 = ~a5858 & i386;
assign a5864 = ~a5862 & ~a5860;
assign a5866 = a5864 & a5852;
assign a5868 = a5502 & ~l818;
assign a5870 = ~a5502 & ~l1128;
assign a5872 = ~a5870 & ~a5868;
assign a5874 = a5872 & ~i388;
assign a5876 = ~a5872 & i388;
assign a5878 = ~a5876 & ~a5874;
assign a5880 = a5878 & a5866;
assign a5882 = a5502 & ~l820;
assign a5884 = ~a5502 & ~l1130;
assign a5886 = ~a5884 & ~a5882;
assign a5888 = a5886 & ~i390;
assign a5890 = ~a5886 & i390;
assign a5892 = ~a5890 & ~a5888;
assign a5894 = a5892 & a5880;
assign a5896 = a5502 & ~l826;
assign a5898 = ~a5502 & ~l1132;
assign a5900 = ~a5898 & ~a5896;
assign a5902 = a5900 & ~i392;
assign a5904 = ~a5900 & i392;
assign a5906 = ~a5904 & ~a5902;
assign a5908 = a5906 & a5894;
assign a5910 = ~a5502 & ~l1134;
assign a5912 = a5502 & l828;
assign a5914 = ~a5912 & ~a5910;
assign a5916 = a5914 & ~i394;
assign a5918 = ~a5914 & i394;
assign a5920 = ~a5918 & ~a5916;
assign a5922 = a5920 & a5908;
assign a5924 = a5502 & ~l832;
assign a5926 = ~a5502 & ~l1136;
assign a5928 = ~a5926 & ~a5924;
assign a5930 = a5928 & ~i396;
assign a5932 = ~a5928 & i396;
assign a5934 = ~a5932 & ~a5930;
assign a5936 = a5934 & a5922;
assign a5938 = ~a5502 & ~l1138;
assign a5940 = a5502 & l834;
assign a5942 = ~a5940 & ~a5938;
assign a5944 = a5942 & ~i398;
assign a5946 = ~a5942 & i398;
assign a5948 = ~a5946 & ~a5944;
assign a5950 = a5948 & a5936;
assign a5952 = a5502 & ~l840;
assign a5954 = ~a5502 & ~l1140;
assign a5956 = ~a5954 & ~a5952;
assign a5958 = a5956 & ~i400;
assign a5960 = ~a5956 & i400;
assign a5962 = ~a5960 & ~a5958;
assign a5964 = a5962 & a5950;
assign a5966 = ~a5502 & ~l1142;
assign a5968 = a5502 & l842;
assign a5970 = ~a5968 & ~a5966;
assign a5972 = a5970 & ~i402;
assign a5974 = ~a5970 & i402;
assign a5976 = ~a5974 & ~a5972;
assign a5978 = a5976 & a5964;
assign a5980 = a5502 & ~l846;
assign a5982 = ~a5502 & ~l1144;
assign a5984 = ~a5982 & ~a5980;
assign a5986 = a5984 & ~i404;
assign a5988 = ~a5984 & i404;
assign a5990 = ~a5988 & ~a5986;
assign a5992 = a5990 & a5978;
assign a5994 = ~a5502 & ~l1146;
assign a5996 = a5502 & l848;
assign a5998 = ~a5996 & ~a5994;
assign a6000 = a5998 & ~i406;
assign a6002 = ~a5998 & i406;
assign a6004 = ~a6002 & ~a6000;
assign a6006 = a6004 & a5992;
assign a6008 = a5502 & ~l854;
assign a6010 = ~a5502 & ~l1148;
assign a6012 = ~a6010 & ~a6008;
assign a6014 = a6012 & ~i408;
assign a6016 = ~a6012 & i408;
assign a6018 = ~a6016 & ~a6014;
assign a6020 = a6018 & a6006;
assign a6022 = ~a5502 & ~l1150;
assign a6024 = a5502 & l856;
assign a6026 = ~a6024 & ~a6022;
assign a6028 = a6026 & ~i410;
assign a6030 = ~a6026 & i410;
assign a6032 = ~a6030 & ~a6028;
assign a6034 = a6032 & a6020;
assign a6036 = a5502 & ~l860;
assign a6038 = ~a5502 & ~l1152;
assign a6040 = ~a6038 & ~a6036;
assign a6042 = a6040 & ~i412;
assign a6044 = ~a6040 & i412;
assign a6046 = ~a6044 & ~a6042;
assign a6048 = a6046 & a6034;
assign a6050 = ~a5502 & ~l1154;
assign a6052 = a5502 & l862;
assign a6054 = ~a6052 & ~a6050;
assign a6056 = a6054 & ~i414;
assign a6058 = ~a6054 & i414;
assign a6060 = ~a6058 & ~a6056;
assign a6062 = a6060 & a6048;
assign a6064 = a5502 & ~l868;
assign a6066 = ~a5502 & ~l1156;
assign a6068 = ~a6066 & ~a6064;
assign a6070 = a6068 & ~i416;
assign a6072 = ~a6068 & i416;
assign a6074 = ~a6072 & ~a6070;
assign a6076 = a6074 & a6062;
assign a6078 = ~a5502 & ~l1158;
assign a6080 = a5502 & l870;
assign a6082 = ~a6080 & ~a6078;
assign a6084 = a6082 & ~i418;
assign a6086 = ~a6082 & i418;
assign a6088 = ~a6086 & ~a6084;
assign a6090 = a6088 & a6076;
assign a6092 = a5502 & ~l874;
assign a6094 = ~a5502 & ~l1160;
assign a6096 = ~a6094 & ~a6092;
assign a6098 = a6096 & ~i420;
assign a6100 = ~a6096 & i420;
assign a6102 = ~a6100 & ~a6098;
assign a6104 = a6102 & a6090;
assign a6106 = ~a5502 & ~l1162;
assign a6108 = a5502 & l876;
assign a6110 = ~a6108 & ~a6106;
assign a6112 = a6110 & ~i422;
assign a6114 = ~a6110 & i422;
assign a6116 = ~a6114 & ~a6112;
assign a6118 = a6116 & a6104;
assign a6120 = a5502 & ~l878;
assign a6122 = ~a5502 & ~l1164;
assign a6124 = ~a6122 & ~a6120;
assign a6126 = a6124 & ~i424;
assign a6128 = ~a6124 & i424;
assign a6130 = ~a6128 & ~a6126;
assign a6132 = a6130 & a6118;
assign a6134 = a5502 & ~l880;
assign a6136 = ~a5502 & ~l1166;
assign a6138 = ~a6136 & ~a6134;
assign a6140 = a6138 & ~i426;
assign a6142 = ~a6138 & i426;
assign a6144 = ~a6142 & ~a6140;
assign a6146 = a6144 & a6132;
assign a6148 = ~a5502 & ~l1168;
assign a6150 = a5502 & l882;
assign a6152 = ~a6150 & ~a6148;
assign a6154 = a6152 & ~i428;
assign a6156 = ~a6152 & i428;
assign a6158 = ~a6156 & ~a6154;
assign a6160 = a6158 & a6146;
assign a6162 = a5502 & ~l884;
assign a6164 = ~a5502 & ~l1170;
assign a6166 = ~a6164 & ~a6162;
assign a6168 = a6166 & ~i430;
assign a6170 = ~a6166 & i430;
assign a6172 = ~a6170 & ~a6168;
assign a6174 = a6172 & a6160;
assign a6176 = a5502 & ~l886;
assign a6178 = ~a5502 & ~l1172;
assign a6180 = ~a6178 & ~a6176;
assign a6182 = a6180 & ~i432;
assign a6184 = ~a6180 & i432;
assign a6186 = ~a6184 & ~a6182;
assign a6188 = a6186 & a6174;
assign a6190 = a5502 & ~l888;
assign a6192 = ~a5502 & ~l1174;
assign a6194 = ~a6192 & ~a6190;
assign a6196 = a6194 & ~i434;
assign a6198 = ~a6194 & i434;
assign a6200 = ~a6198 & ~a6196;
assign a6202 = a6200 & a6188;
assign a6204 = a5502 & ~l892;
assign a6206 = ~a5502 & ~l1176;
assign a6208 = ~a6206 & ~a6204;
assign a6210 = a6208 & ~i436;
assign a6212 = ~a6208 & i436;
assign a6214 = ~a6212 & ~a6210;
assign a6216 = a6214 & a6202;
assign a6218 = a5502 & ~l894;
assign a6220 = ~a5502 & ~l1178;
assign a6222 = ~a6220 & ~a6218;
assign a6224 = a6222 & ~i438;
assign a6226 = ~a6222 & i438;
assign a6228 = ~a6226 & ~a6224;
assign a6230 = a6228 & a6216;
assign a6232 = a5502 & ~l896;
assign a6234 = ~a5502 & ~l1180;
assign a6236 = ~a6234 & ~a6232;
assign a6238 = a6236 & ~i440;
assign a6240 = ~a6236 & i440;
assign a6242 = ~a6240 & ~a6238;
assign a6244 = a6242 & a6230;
assign a6246 = a5502 & ~l898;
assign a6248 = ~a5502 & ~l1182;
assign a6250 = ~a6248 & ~a6246;
assign a6252 = a6250 & ~i442;
assign a6254 = ~a6250 & i442;
assign a6256 = ~a6254 & ~a6252;
assign a6258 = a6256 & a6244;
assign a6260 = a5502 & ~l900;
assign a6262 = ~a5502 & ~l1184;
assign a6264 = ~a6262 & ~a6260;
assign a6266 = a6264 & ~i444;
assign a6268 = ~a6264 & i444;
assign a6270 = ~a6268 & ~a6266;
assign a6272 = a6270 & a6258;
assign a6274 = a5502 & ~l902;
assign a6276 = ~a5502 & ~l1186;
assign a6278 = ~a6276 & ~a6274;
assign a6280 = a6278 & ~i446;
assign a6282 = ~a6278 & i446;
assign a6284 = ~a6282 & ~a6280;
assign a6286 = a6284 & a6272;
assign a6288 = a5502 & ~l908;
assign a6290 = ~a5502 & ~l1188;
assign a6292 = ~a6290 & ~a6288;
assign a6294 = a6292 & ~i448;
assign a6296 = ~a6292 & i448;
assign a6298 = ~a6296 & ~a6294;
assign a6300 = a6298 & a6286;
assign a6302 = ~a5502 & ~l1190;
assign a6304 = a5502 & l910;
assign a6306 = ~a6304 & ~a6302;
assign a6308 = a6306 & ~i450;
assign a6310 = ~a6306 & i450;
assign a6312 = ~a6310 & ~a6308;
assign a6314 = a6312 & a6300;
assign a6316 = a5502 & ~l914;
assign a6318 = ~a5502 & ~l1192;
assign a6320 = ~a6318 & ~a6316;
assign a6322 = a6320 & ~i452;
assign a6324 = ~a6320 & i452;
assign a6326 = ~a6324 & ~a6322;
assign a6328 = a6326 & a6314;
assign a6330 = ~a5502 & ~l1194;
assign a6332 = a5502 & l916;
assign a6334 = ~a6332 & ~a6330;
assign a6336 = a6334 & ~i454;
assign a6338 = ~a6334 & i454;
assign a6340 = ~a6338 & ~a6336;
assign a6342 = a6340 & a6328;
assign a6344 = a5502 & ~l922;
assign a6346 = ~a5502 & ~l1196;
assign a6348 = ~a6346 & ~a6344;
assign a6350 = a6348 & ~i456;
assign a6352 = ~a6348 & i456;
assign a6354 = ~a6352 & ~a6350;
assign a6356 = a6354 & a6342;
assign a6358 = ~a5502 & ~l1198;
assign a6360 = a5502 & l924;
assign a6362 = ~a6360 & ~a6358;
assign a6364 = a6362 & ~i458;
assign a6366 = ~a6362 & i458;
assign a6368 = ~a6366 & ~a6364;
assign a6370 = a6368 & a6356;
assign a6372 = a5502 & ~l928;
assign a6374 = ~a5502 & ~l1200;
assign a6376 = ~a6374 & ~a6372;
assign a6378 = a6376 & ~i460;
assign a6380 = ~a6376 & i460;
assign a6382 = ~a6380 & ~a6378;
assign a6384 = a6382 & a6370;
assign a6386 = ~a5502 & ~l1202;
assign a6388 = a5502 & l930;
assign a6390 = ~a6388 & ~a6386;
assign a6392 = a6390 & ~i462;
assign a6394 = ~a6390 & i462;
assign a6396 = ~a6394 & ~a6392;
assign a6398 = a6396 & a6384;
assign a6400 = a5502 & ~l936;
assign a6402 = ~a5502 & ~l1204;
assign a6404 = ~a6402 & ~a6400;
assign a6406 = a6404 & ~i464;
assign a6408 = ~a6404 & i464;
assign a6410 = ~a6408 & ~a6406;
assign a6412 = a6410 & a6398;
assign a6414 = ~a5502 & ~l1206;
assign a6416 = a5502 & l938;
assign a6418 = ~a6416 & ~a6414;
assign a6420 = a6418 & ~i466;
assign a6422 = ~a6418 & i466;
assign a6424 = ~a6422 & ~a6420;
assign a6426 = a6424 & a6412;
assign a6428 = a5502 & ~l942;
assign a6430 = ~a5502 & ~l1208;
assign a6432 = ~a6430 & ~a6428;
assign a6434 = a6432 & ~i468;
assign a6436 = ~a6432 & i468;
assign a6438 = ~a6436 & ~a6434;
assign a6440 = a6438 & a6426;
assign a6442 = ~a5502 & ~l1210;
assign a6444 = a5502 & l944;
assign a6446 = ~a6444 & ~a6442;
assign a6448 = a6446 & ~i470;
assign a6450 = ~a6446 & i470;
assign a6452 = ~a6450 & ~a6448;
assign a6454 = a6452 & a6440;
assign a6456 = a5502 & ~l950;
assign a6458 = ~a5502 & ~l1212;
assign a6460 = ~a6458 & ~a6456;
assign a6462 = a6460 & ~i472;
assign a6464 = ~a6460 & i472;
assign a6466 = ~a6464 & ~a6462;
assign a6468 = a6466 & a6454;
assign a6470 = ~a5502 & ~l1214;
assign a6472 = a5502 & l952;
assign a6474 = ~a6472 & ~a6470;
assign a6476 = a6474 & ~i474;
assign a6478 = ~a6474 & i474;
assign a6480 = ~a6478 & ~a6476;
assign a6482 = a6480 & a6468;
assign a6484 = a5502 & ~l956;
assign a6486 = ~a5502 & ~l1216;
assign a6488 = ~a6486 & ~a6484;
assign a6490 = a6488 & ~i476;
assign a6492 = ~a6488 & i476;
assign a6494 = ~a6492 & ~a6490;
assign a6496 = a6494 & a6482;
assign a6498 = ~a5502 & ~l1218;
assign a6500 = a5502 & l958;
assign a6502 = ~a6500 & ~a6498;
assign a6504 = a6502 & ~i478;
assign a6506 = ~a6502 & i478;
assign a6508 = ~a6506 & ~a6504;
assign a6510 = a6508 & a6496;
assign a6512 = a5502 & ~l960;
assign a6514 = ~a5502 & ~l1220;
assign a6516 = ~a6514 & ~a6512;
assign a6518 = a6516 & ~i480;
assign a6520 = ~a6516 & i480;
assign a6522 = ~a6520 & ~a6518;
assign a6524 = a6522 & a6510;
assign a6526 = a5502 & ~l962;
assign a6528 = ~a5502 & ~l1222;
assign a6530 = ~a6528 & ~a6526;
assign a6532 = a6530 & ~i482;
assign a6534 = ~a6530 & i482;
assign a6536 = ~a6534 & ~a6532;
assign a6538 = a6536 & a6524;
assign a6540 = ~a5502 & ~l1224;
assign a6542 = a5502 & l964;
assign a6544 = ~a6542 & ~a6540;
assign a6546 = a6544 & ~i484;
assign a6548 = ~a6544 & i484;
assign a6550 = ~a6548 & ~a6546;
assign a6552 = a6550 & a6538;
assign a6554 = a5502 & ~l966;
assign a6556 = ~a5502 & ~l1226;
assign a6558 = ~a6556 & ~a6554;
assign a6560 = a6558 & ~i486;
assign a6562 = ~a6558 & i486;
assign a6564 = ~a6562 & ~a6560;
assign a6566 = a6564 & a6552;
assign a6568 = a5502 & ~l968;
assign a6570 = ~a5502 & ~l1228;
assign a6572 = ~a6570 & ~a6568;
assign a6574 = a6572 & ~i488;
assign a6576 = ~a6572 & i488;
assign a6578 = ~a6576 & ~a6574;
assign a6580 = a6578 & a6566;
assign a6582 = a5502 & ~l970;
assign a6584 = ~a5502 & ~l1230;
assign a6586 = ~a6584 & ~a6582;
assign a6588 = a6586 & ~i490;
assign a6590 = ~a6586 & i490;
assign a6592 = ~a6590 & ~a6588;
assign a6594 = a6592 & a6580;
assign a6596 = a5502 & ~l974;
assign a6598 = ~a5502 & ~l1232;
assign a6600 = ~a6598 & ~a6596;
assign a6602 = a6600 & ~i492;
assign a6604 = ~a6600 & i492;
assign a6606 = ~a6604 & ~a6602;
assign a6608 = a6606 & a6594;
assign a6610 = a5502 & ~l976;
assign a6612 = ~a5502 & ~l1234;
assign a6614 = ~a6612 & ~a6610;
assign a6616 = a6614 & ~i494;
assign a6618 = ~a6614 & i494;
assign a6620 = ~a6618 & ~a6616;
assign a6622 = a6620 & a6608;
assign a6624 = a5502 & ~l978;
assign a6626 = ~a5502 & ~l1236;
assign a6628 = ~a6626 & ~a6624;
assign a6630 = a6628 & ~i496;
assign a6632 = ~a6628 & i496;
assign a6634 = ~a6632 & ~a6630;
assign a6636 = a6634 & a6622;
assign a6638 = a5502 & ~l980;
assign a6640 = ~a5502 & ~l1238;
assign a6642 = ~a6640 & ~a6638;
assign a6644 = a6642 & ~i498;
assign a6646 = ~a6642 & i498;
assign a6648 = ~a6646 & ~a6644;
assign a6650 = a6648 & a6636;
assign a6652 = a5502 & ~l982;
assign a6654 = ~a5502 & ~l1240;
assign a6656 = ~a6654 & ~a6652;
assign a6658 = a6656 & ~i500;
assign a6660 = ~a6656 & i500;
assign a6662 = ~a6660 & ~a6658;
assign a6664 = a6662 & a6650;
assign a6666 = a5502 & ~l984;
assign a6668 = ~a5502 & ~l1242;
assign a6670 = ~a6668 & ~a6666;
assign a6672 = a6670 & ~i502;
assign a6674 = ~a6670 & i502;
assign a6676 = ~a6674 & ~a6672;
assign a6678 = a6676 & a6664;
assign a6680 = a5502 & ~l990;
assign a6682 = ~a5502 & ~l1244;
assign a6684 = ~a6682 & ~a6680;
assign a6686 = a6684 & ~i504;
assign a6688 = ~a6684 & i504;
assign a6690 = ~a6688 & ~a6686;
assign a6692 = a6690 & a6678;
assign a6694 = ~a5502 & ~l1246;
assign a6696 = a5502 & l992;
assign a6698 = ~a6696 & ~a6694;
assign a6700 = a6698 & ~i506;
assign a6702 = ~a6698 & i506;
assign a6704 = ~a6702 & ~a6700;
assign a6706 = a6704 & a6692;
assign a6708 = a5502 & ~l996;
assign a6710 = ~a5502 & ~l1248;
assign a6712 = ~a6710 & ~a6708;
assign a6714 = a6712 & ~i508;
assign a6716 = ~a6712 & i508;
assign a6718 = ~a6716 & ~a6714;
assign a6720 = a6718 & a6706;
assign a6722 = ~a5502 & ~l1250;
assign a6724 = a5502 & l998;
assign a6726 = ~a6724 & ~a6722;
assign a6728 = a6726 & ~i510;
assign a6730 = ~a6726 & i510;
assign a6732 = ~a6730 & ~a6728;
assign a6734 = a6732 & a6720;
assign a6736 = a5502 & ~l1004;
assign a6738 = ~a5502 & ~l1252;
assign a6740 = ~a6738 & ~a6736;
assign a6742 = a6740 & ~i512;
assign a6744 = ~a6740 & i512;
assign a6746 = ~a6744 & ~a6742;
assign a6748 = a6746 & a6734;
assign a6750 = ~a5502 & ~l1254;
assign a6752 = a5502 & l1006;
assign a6754 = ~a6752 & ~a6750;
assign a6756 = a6754 & ~i514;
assign a6758 = ~a6754 & i514;
assign a6760 = ~a6758 & ~a6756;
assign a6762 = a6760 & a6748;
assign a6764 = a5502 & ~l1010;
assign a6766 = ~a5502 & ~l1256;
assign a6768 = ~a6766 & ~a6764;
assign a6770 = a6768 & ~i516;
assign a6772 = ~a6768 & i516;
assign a6774 = ~a6772 & ~a6770;
assign a6776 = a6774 & a6762;
assign a6778 = ~a5502 & ~l1258;
assign a6780 = a5502 & l1012;
assign a6782 = ~a6780 & ~a6778;
assign a6784 = a6782 & ~i518;
assign a6786 = ~a6782 & i518;
assign a6788 = ~a6786 & ~a6784;
assign a6790 = a6788 & a6776;
assign a6792 = a5502 & ~l1018;
assign a6794 = ~a5502 & ~l1260;
assign a6796 = ~a6794 & ~a6792;
assign a6798 = a6796 & ~i520;
assign a6800 = ~a6796 & i520;
assign a6802 = ~a6800 & ~a6798;
assign a6804 = a6802 & a6790;
assign a6806 = ~a5502 & ~l1262;
assign a6808 = a5502 & l1020;
assign a6810 = ~a6808 & ~a6806;
assign a6812 = a6810 & ~i522;
assign a6814 = ~a6810 & i522;
assign a6816 = ~a6814 & ~a6812;
assign a6818 = a6816 & a6804;
assign a6820 = a5502 & ~l1024;
assign a6822 = ~a5502 & ~l1264;
assign a6824 = ~a6822 & ~a6820;
assign a6826 = a6824 & ~i524;
assign a6828 = ~a6824 & i524;
assign a6830 = ~a6828 & ~a6826;
assign a6832 = a6830 & a6818;
assign a6834 = ~a5502 & ~l1266;
assign a6836 = a5502 & l1026;
assign a6838 = ~a6836 & ~a6834;
assign a6840 = a6838 & ~i526;
assign a6842 = ~a6838 & i526;
assign a6844 = ~a6842 & ~a6840;
assign a6846 = a6844 & a6832;
assign a6848 = a5502 & ~l1032;
assign a6850 = ~a5502 & ~l1268;
assign a6852 = ~a6850 & ~a6848;
assign a6854 = a6852 & ~i528;
assign a6856 = ~a6852 & i528;
assign a6858 = ~a6856 & ~a6854;
assign a6860 = a6858 & a6846;
assign a6862 = ~a5502 & ~l1270;
assign a6864 = a5502 & l1034;
assign a6866 = ~a6864 & ~a6862;
assign a6868 = a6866 & ~i530;
assign a6870 = ~a6866 & i530;
assign a6872 = ~a6870 & ~a6868;
assign a6874 = a6872 & a6860;
assign a6876 = a5502 & ~l1038;
assign a6878 = ~a5502 & ~l1272;
assign a6880 = ~a6878 & ~a6876;
assign a6882 = a6880 & ~i532;
assign a6884 = ~a6880 & i532;
assign a6886 = ~a6884 & ~a6882;
assign a6888 = a6886 & a6874;
assign a6890 = ~a5502 & ~l1274;
assign a6892 = a5502 & l1040;
assign a6894 = ~a6892 & ~a6890;
assign a6896 = a6894 & ~i534;
assign a6898 = ~a6894 & i534;
assign a6900 = ~a6898 & ~a6896;
assign a6902 = a6900 & a6888;
assign a6904 = a5502 & ~l1042;
assign a6906 = ~a5502 & ~l1276;
assign a6908 = ~a6906 & ~a6904;
assign a6910 = a6908 & ~i536;
assign a6912 = ~a6908 & i536;
assign a6914 = ~a6912 & ~a6910;
assign a6916 = a6914 & a6902;
assign a6918 = a5502 & ~l1044;
assign a6920 = ~a5502 & ~l1278;
assign a6922 = ~a6920 & ~a6918;
assign a6924 = a6922 & ~i538;
assign a6926 = ~a6922 & i538;
assign a6928 = ~a6926 & ~a6924;
assign a6930 = a6928 & a6916;
assign a6932 = ~a5502 & ~l1280;
assign a6934 = a5502 & l1046;
assign a6936 = ~a6934 & ~a6932;
assign a6938 = a6936 & ~i540;
assign a6940 = ~a6936 & i540;
assign a6942 = ~a6940 & ~a6938;
assign a6944 = a6942 & a6930;
assign a6946 = a5502 & ~l1048;
assign a6948 = ~a5502 & ~l1282;
assign a6950 = ~a6948 & ~a6946;
assign a6952 = a6950 & ~i542;
assign a6954 = ~a6950 & i542;
assign a6956 = ~a6954 & ~a6952;
assign a6958 = a6956 & a6944;
assign a6960 = a5502 & ~l1050;
assign a6962 = ~a5502 & ~l1284;
assign a6964 = ~a6962 & ~a6960;
assign a6966 = a6964 & ~i544;
assign a6968 = ~a6964 & i544;
assign a6970 = ~a6968 & ~a6966;
assign a6972 = a6970 & a6958;
assign a6974 = a5502 & ~l1052;
assign a6976 = ~a5502 & ~l1286;
assign a6978 = ~a6976 & ~a6974;
assign a6980 = a6978 & ~i546;
assign a6982 = ~a6978 & i546;
assign a6984 = ~a6982 & ~a6980;
assign a6986 = a6984 & a6972;
assign a6988 = a5502 & ~l1056;
assign a6990 = ~a5502 & ~l1288;
assign a6992 = ~a6990 & ~a6988;
assign a6994 = a6992 & ~i548;
assign a6996 = ~a6992 & i548;
assign a6998 = ~a6996 & ~a6994;
assign a7000 = a6998 & a6986;
assign a7002 = a5502 & ~l1058;
assign a7004 = ~a5502 & ~l1290;
assign a7006 = ~a7004 & ~a7002;
assign a7008 = a7006 & ~i550;
assign a7010 = ~a7006 & i550;
assign a7012 = ~a7010 & ~a7008;
assign a7014 = a7012 & a7000;
assign a7016 = a5502 & ~l1060;
assign a7018 = ~a5502 & ~l1292;
assign a7020 = ~a7018 & ~a7016;
assign a7022 = a7020 & ~i552;
assign a7024 = ~a7020 & i552;
assign a7026 = ~a7024 & ~a7022;
assign a7028 = a7026 & a7014;
assign a7030 = a5502 & ~l1062;
assign a7032 = ~a5502 & ~l1294;
assign a7034 = ~a7032 & ~a7030;
assign a7036 = a7034 & ~i554;
assign a7038 = ~a7034 & i554;
assign a7040 = ~a7038 & ~a7036;
assign a7042 = a7040 & a7028;
assign a7044 = a5502 & ~l1064;
assign a7046 = ~a5502 & ~l1296;
assign a7048 = ~a7046 & ~a7044;
assign a7050 = a7048 & ~i556;
assign a7052 = ~a7048 & i556;
assign a7054 = ~a7052 & ~a7050;
assign a7056 = a7054 & a7042;
assign a7058 = a5502 & ~l1066;
assign a7060 = ~a5502 & ~l1298;
assign a7062 = ~a7060 & ~a7058;
assign a7064 = a7062 & ~i558;
assign a7066 = ~a7062 & i558;
assign a7068 = ~a7066 & ~a7064;
assign a7070 = a7068 & a7056;
assign a7072 = a5502 & ~l1068;
assign a7074 = ~a5502 & ~l1300;
assign a7076 = ~a7074 & ~a7072;
assign a7078 = a7076 & ~i560;
assign a7080 = ~a7076 & i560;
assign a7082 = ~a7080 & ~a7078;
assign a7084 = a7082 & a7070;
assign a7086 = a5502 & ~l1070;
assign a7088 = ~a5502 & ~l1302;
assign a7090 = ~a7088 & ~a7086;
assign a7092 = a7090 & ~i562;
assign a7094 = ~a7090 & i562;
assign a7096 = ~a7094 & ~a7092;
assign a7098 = a7096 & a7084;
assign a7100 = a5502 & ~l1072;
assign a7102 = ~a5502 & ~l1304;
assign a7104 = ~a7102 & ~a7100;
assign a7106 = a7104 & ~i564;
assign a7108 = ~a7104 & i564;
assign a7110 = ~a7108 & ~a7106;
assign a7112 = a7110 & a7098;
assign a7114 = a5502 & ~l1074;
assign a7116 = ~a5502 & ~l1306;
assign a7118 = ~a7116 & ~a7114;
assign a7120 = a7118 & ~i566;
assign a7122 = ~a7118 & i566;
assign a7124 = ~a7122 & ~a7120;
assign a7126 = a7124 & a7112;
assign a7128 = ~l584 & ~l582;
assign a7130 = ~a7128 & l580;
assign a7132 = ~l594 & ~l592;
assign a7134 = ~a7132 & l590;
assign a7136 = ~l604 & ~l602;
assign a7138 = ~a7136 & l600;
assign a7140 = ~l614 & ~l612;
assign a7142 = ~a7140 & l610;
assign a7144 = ~l624 & ~l622;
assign a7146 = ~a7144 & l620;
assign a7148 = ~l634 & ~l632;
assign a7150 = ~a7148 & l630;
assign a7152 = ~l644 & ~l642;
assign a7154 = ~a7152 & l640;
assign a7156 = ~l654 & ~l652;
assign a7158 = ~a7156 & l650;
assign a7160 = ~l664 & ~l662;
assign a7162 = ~a7160 & l660;
assign a7164 = ~l674 & ~l672;
assign a7166 = ~a7164 & l670;
assign a7168 = ~l684 & ~l682;
assign a7170 = ~a7168 & l680;
assign a7172 = ~l694 & ~l692;
assign a7174 = ~a7172 & l690;
assign a7176 = ~l704 & ~l702;
assign a7178 = ~a7176 & l700;
assign a7180 = ~l714 & ~l712;
assign a7182 = ~a7180 & l710;
assign a7184 = ~l724 & ~l722;
assign a7186 = ~a7184 & l720;
assign a7188 = ~l734 & ~l732;
assign a7190 = ~a7188 & l730;
assign a7192 = l742 & l740;
assign a7194 = ~l746 & l744;
assign a7196 = l756 & l754;
assign a7198 = ~l760 & l758;
assign a7200 = l770 & l768;
assign a7202 = ~l774 & l772;
assign a7204 = l784 & l782;
assign a7206 = ~l788 & l786;
assign a7208 = a1414 & l796;
assign a7210 = a1872 & l814;
assign a7212 = l824 & l822;
assign a7214 = ~l828 & l826;
assign a7216 = l838 & l836;
assign a7218 = ~l842 & l840;
assign a7220 = l852 & l850;
assign a7222 = ~l856 & l854;
assign a7224 = l866 & l864;
assign a7226 = ~l870 & l868;
assign a7228 = a2112 & l878;
assign a7230 = a2570 & l896;
assign a7232 = l906 & l904;
assign a7234 = ~l910 & l908;
assign a7236 = l920 & l918;
assign a7238 = ~l924 & l922;
assign a7240 = l934 & l932;
assign a7242 = ~l938 & l936;
assign a7244 = l948 & l946;
assign a7246 = ~l952 & l950;
assign a7248 = a2810 & l960;
assign a7250 = a3268 & l978;
assign a7252 = l988 & l986;
assign a7254 = ~l992 & l990;
assign a7256 = l1002 & l1000;
assign a7258 = ~l1006 & l1004;
assign a7260 = l1016 & l1014;
assign a7262 = ~l1020 & l1018;
assign a7264 = l1030 & l1028;
assign a7266 = ~l1034 & l1032;
assign a7268 = a3508 & l1042;
assign a7270 = a3966 & l1060;
assign a7272 = l1078 & l1076;
assign a7274 = l1086 & l1084;
assign a7276 = l1094 & l1092;
assign a7278 = l1102 & l1100;
assign a7280 = l1112 & l1110;
assign a7282 = a7280 & l1108;
assign a7284 = l1128 & l1126;
assign a7286 = a7284 & l1124;
assign a7288 = l1134 & l1132;
assign a7290 = l1142 & l1140;
assign a7292 = l1150 & l1148;
assign a7294 = l1158 & l1156;
assign a7296 = l1168 & l1166;
assign a7298 = a7296 & l1164;
assign a7300 = l1184 & l1182;
assign a7302 = a7300 & l1180;
assign a7304 = l1190 & l1188;
assign a7306 = l1198 & l1196;
assign a7308 = l1206 & l1204;
assign a7310 = l1214 & l1212;
assign a7312 = l1224 & l1222;
assign a7314 = a7312 & l1220;
assign a7316 = l1240 & l1238;
assign a7318 = a7316 & l1236;
assign a7320 = l1246 & l1244;
assign a7322 = l1254 & l1252;
assign a7324 = l1262 & l1260;
assign a7326 = l1270 & l1268;
assign a7328 = l1280 & l1278;
assign a7330 = a7328 & l1276;
assign a7332 = l1296 & l1294;
assign a7334 = a7332 & l1292;
assign a7336 = ~l974 & ~l892;
assign a7338 = l974 & l892;
assign a7340 = ~a7338 & ~a7336;
assign a7342 = a2740 & a2042;
assign a7344 = a7342 & ~a7340;
assign a7346 = ~l892 & ~l810;
assign a7348 = l892 & l810;
assign a7350 = ~a7348 & ~a7346;
assign a7352 = ~a7350 & a2042;
assign a7354 = ~l974 & ~l810;
assign a7356 = l974 & l810;
assign a7358 = ~a7356 & ~a7354;
assign a7360 = ~a7358 & a2740;
assign a7362 = ~l1056 & ~l810;
assign a7364 = l1056 & l810;
assign a7366 = ~a7364 & ~a7362;
assign a7368 = ~a7366 & a3438;
assign a7370 = ~a7368 & ~a7360;
assign a7372 = a7370 & ~a7352;
assign a7374 = ~a7372 & a1344;
assign a7376 = ~l1056 & ~l892;
assign a7378 = l1056 & l892;
assign a7380 = ~a7378 & ~a7376;
assign a7382 = a3438 & a2042;
assign a7384 = a7382 & ~a7380;
assign a7386 = ~l1056 & ~l974;
assign a7388 = l1056 & l974;
assign a7390 = ~a7388 & ~a7386;
assign a7392 = a3438 & a2740;
assign a7394 = a7392 & ~a7390;
assign a7396 = ~a7394 & ~a7384;
assign a7398 = a7396 & ~a7374;
assign a7400 = a7398 & ~a7344;
assign a7402 = ~a7400 & l1068;
assign a7404 = a7128 & ~l580;
assign a7406 = l584 & ~l582;
assign a7408 = a7406 & ~l580;
assign a7410 = ~l584 & l582;
assign a7412 = a7410 & ~l580;
assign a7414 = l584 & l582;
assign a7416 = a7414 & ~l580;
assign a7418 = a7128 & l580;
assign a7420 = ~l588 & ~l586;
assign a7422 = l588 & ~l586;
assign a7424 = ~l588 & l586;
assign a7426 = l588 & l586;
assign a7428 = a7426 & ~l1032;
assign a7430 = a7428 & ~a7424;
assign a7432 = a7424 & ~l1018;
assign a7434 = ~a7432 & ~a7430;
assign a7436 = ~a7434 & ~a7422;
assign a7438 = a7422 & ~l1004;
assign a7440 = ~a7438 & ~a7436;
assign a7442 = ~a7440 & ~a7420;
assign a7444 = a7420 & ~l990;
assign a7446 = ~a7444 & ~a7442;
assign a7448 = ~a7446 & a7418;
assign a7450 = a7448 & ~a7416;
assign a7452 = a7426 & ~l950;
assign a7454 = a7452 & ~a7424;
assign a7456 = a7424 & ~l936;
assign a7458 = ~a7456 & ~a7454;
assign a7460 = ~a7458 & ~a7422;
assign a7462 = a7422 & ~l922;
assign a7464 = ~a7462 & ~a7460;
assign a7466 = ~a7464 & ~a7420;
assign a7468 = a7420 & ~l908;
assign a7470 = ~a7468 & ~a7466;
assign a7472 = ~a7470 & a7416;
assign a7474 = ~a7472 & ~a7450;
assign a7476 = ~a7474 & ~a7412;
assign a7478 = a7426 & ~l868;
assign a7480 = a7478 & ~a7424;
assign a7482 = a7424 & ~l854;
assign a7484 = ~a7482 & ~a7480;
assign a7486 = ~a7484 & ~a7422;
assign a7488 = a7422 & ~l840;
assign a7490 = ~a7488 & ~a7486;
assign a7492 = ~a7490 & ~a7420;
assign a7494 = a7420 & ~l826;
assign a7496 = ~a7494 & ~a7492;
assign a7498 = ~a7496 & a7412;
assign a7500 = ~a7498 & ~a7476;
assign a7502 = ~a7500 & ~a7408;
assign a7504 = a7426 & ~l786;
assign a7506 = a7504 & ~a7424;
assign a7508 = a7424 & ~l772;
assign a7510 = ~a7508 & ~a7506;
assign a7512 = ~a7510 & ~a7422;
assign a7514 = a7422 & ~l758;
assign a7516 = ~a7514 & ~a7512;
assign a7518 = ~a7516 & ~a7420;
assign a7520 = a7420 & ~l744;
assign a7522 = ~a7520 & ~a7518;
assign a7524 = ~a7522 & a7408;
assign a7526 = ~a7524 & ~a7502;
assign a7528 = a7526 & ~l740;
assign a7530 = ~a7526 & l740;
assign a7532 = ~a7530 & ~a7528;
assign a7534 = a7426 & l1034;
assign a7536 = a7534 & ~a7424;
assign a7538 = a7424 & l1020;
assign a7540 = ~a7538 & ~a7536;
assign a7542 = ~a7540 & ~a7422;
assign a7544 = a7422 & l1006;
assign a7546 = ~a7544 & ~a7542;
assign a7548 = ~a7546 & ~a7420;
assign a7550 = a7420 & l992;
assign a7552 = ~a7550 & ~a7548;
assign a7554 = ~a7552 & a7418;
assign a7556 = a7554 & ~a7416;
assign a7558 = a7426 & l952;
assign a7560 = a7558 & ~a7424;
assign a7562 = a7424 & l938;
assign a7564 = ~a7562 & ~a7560;
assign a7566 = ~a7564 & ~a7422;
assign a7568 = a7422 & l924;
assign a7570 = ~a7568 & ~a7566;
assign a7572 = ~a7570 & ~a7420;
assign a7574 = a7420 & l910;
assign a7576 = ~a7574 & ~a7572;
assign a7578 = ~a7576 & a7416;
assign a7580 = ~a7578 & ~a7556;
assign a7582 = ~a7580 & ~a7412;
assign a7584 = a7426 & l870;
assign a7586 = a7584 & ~a7424;
assign a7588 = a7424 & l856;
assign a7590 = ~a7588 & ~a7586;
assign a7592 = ~a7590 & ~a7422;
assign a7594 = a7422 & l842;
assign a7596 = ~a7594 & ~a7592;
assign a7598 = ~a7596 & ~a7420;
assign a7600 = a7420 & l828;
assign a7602 = ~a7600 & ~a7598;
assign a7604 = ~a7602 & a7412;
assign a7606 = ~a7604 & ~a7582;
assign a7608 = ~a7606 & ~a7408;
assign a7610 = a7426 & l788;
assign a7612 = a7610 & ~a7424;
assign a7614 = a7424 & l774;
assign a7616 = ~a7614 & ~a7612;
assign a7618 = ~a7616 & ~a7422;
assign a7620 = a7422 & l760;
assign a7622 = ~a7620 & ~a7618;
assign a7624 = ~a7622 & ~a7420;
assign a7626 = a7420 & l746;
assign a7628 = ~a7626 & ~a7624;
assign a7630 = ~a7628 & a7408;
assign a7632 = ~a7630 & ~a7608;
assign a7634 = a7632 & ~l742;
assign a7636 = ~a7632 & l742;
assign a7638 = ~a7636 & ~a7634;
assign a7640 = a7638 & a7532;
assign a7642 = ~a7640 & ~a7404;
assign a7644 = a7132 & ~l590;
assign a7646 = l594 & ~l592;
assign a7648 = a7646 & ~l590;
assign a7650 = ~l594 & l592;
assign a7652 = a7650 & ~l590;
assign a7654 = l594 & l592;
assign a7656 = a7654 & ~l590;
assign a7658 = a7132 & l590;
assign a7660 = ~l598 & ~l596;
assign a7662 = l598 & ~l596;
assign a7664 = ~l598 & l596;
assign a7666 = l598 & l596;
assign a7668 = a7666 & ~l1032;
assign a7670 = a7668 & ~a7664;
assign a7672 = a7664 & ~l1018;
assign a7674 = ~a7672 & ~a7670;
assign a7676 = ~a7674 & ~a7662;
assign a7678 = a7662 & ~l1004;
assign a7680 = ~a7678 & ~a7676;
assign a7682 = ~a7680 & ~a7660;
assign a7684 = a7660 & ~l990;
assign a7686 = ~a7684 & ~a7682;
assign a7688 = ~a7686 & a7658;
assign a7690 = a7688 & ~a7656;
assign a7692 = a7666 & ~l950;
assign a7694 = a7692 & ~a7664;
assign a7696 = a7664 & ~l936;
assign a7698 = ~a7696 & ~a7694;
assign a7700 = ~a7698 & ~a7662;
assign a7702 = a7662 & ~l922;
assign a7704 = ~a7702 & ~a7700;
assign a7706 = ~a7704 & ~a7660;
assign a7708 = a7660 & ~l908;
assign a7710 = ~a7708 & ~a7706;
assign a7712 = ~a7710 & a7656;
assign a7714 = ~a7712 & ~a7690;
assign a7716 = ~a7714 & ~a7652;
assign a7718 = a7666 & ~l868;
assign a7720 = a7718 & ~a7664;
assign a7722 = a7664 & ~l854;
assign a7724 = ~a7722 & ~a7720;
assign a7726 = ~a7724 & ~a7662;
assign a7728 = a7662 & ~l840;
assign a7730 = ~a7728 & ~a7726;
assign a7732 = ~a7730 & ~a7660;
assign a7734 = a7660 & ~l826;
assign a7736 = ~a7734 & ~a7732;
assign a7738 = ~a7736 & a7652;
assign a7740 = ~a7738 & ~a7716;
assign a7742 = ~a7740 & ~a7648;
assign a7744 = a7666 & ~l786;
assign a7746 = a7744 & ~a7664;
assign a7748 = a7664 & ~l772;
assign a7750 = ~a7748 & ~a7746;
assign a7752 = ~a7750 & ~a7662;
assign a7754 = a7662 & ~l758;
assign a7756 = ~a7754 & ~a7752;
assign a7758 = ~a7756 & ~a7660;
assign a7760 = a7660 & ~l744;
assign a7762 = ~a7760 & ~a7758;
assign a7764 = ~a7762 & a7648;
assign a7766 = ~a7764 & ~a7742;
assign a7768 = a7766 & ~l754;
assign a7770 = ~a7766 & l754;
assign a7772 = ~a7770 & ~a7768;
assign a7774 = a7666 & l1034;
assign a7776 = a7774 & ~a7664;
assign a7778 = a7664 & l1020;
assign a7780 = ~a7778 & ~a7776;
assign a7782 = ~a7780 & ~a7662;
assign a7784 = a7662 & l1006;
assign a7786 = ~a7784 & ~a7782;
assign a7788 = ~a7786 & ~a7660;
assign a7790 = a7660 & l992;
assign a7792 = ~a7790 & ~a7788;
assign a7794 = ~a7792 & a7658;
assign a7796 = a7794 & ~a7656;
assign a7798 = a7666 & l952;
assign a7800 = a7798 & ~a7664;
assign a7802 = a7664 & l938;
assign a7804 = ~a7802 & ~a7800;
assign a7806 = ~a7804 & ~a7662;
assign a7808 = a7662 & l924;
assign a7810 = ~a7808 & ~a7806;
assign a7812 = ~a7810 & ~a7660;
assign a7814 = a7660 & l910;
assign a7816 = ~a7814 & ~a7812;
assign a7818 = ~a7816 & a7656;
assign a7820 = ~a7818 & ~a7796;
assign a7822 = ~a7820 & ~a7652;
assign a7824 = a7666 & l870;
assign a7826 = a7824 & ~a7664;
assign a7828 = a7664 & l856;
assign a7830 = ~a7828 & ~a7826;
assign a7832 = ~a7830 & ~a7662;
assign a7834 = a7662 & l842;
assign a7836 = ~a7834 & ~a7832;
assign a7838 = ~a7836 & ~a7660;
assign a7840 = a7660 & l828;
assign a7842 = ~a7840 & ~a7838;
assign a7844 = ~a7842 & a7652;
assign a7846 = ~a7844 & ~a7822;
assign a7848 = ~a7846 & ~a7648;
assign a7850 = a7666 & l788;
assign a7852 = a7850 & ~a7664;
assign a7854 = a7664 & l774;
assign a7856 = ~a7854 & ~a7852;
assign a7858 = ~a7856 & ~a7662;
assign a7860 = a7662 & l760;
assign a7862 = ~a7860 & ~a7858;
assign a7864 = ~a7862 & ~a7660;
assign a7866 = a7660 & l746;
assign a7868 = ~a7866 & ~a7864;
assign a7870 = ~a7868 & a7648;
assign a7872 = ~a7870 & ~a7848;
assign a7874 = a7872 & ~l756;
assign a7876 = ~a7872 & l756;
assign a7878 = ~a7876 & ~a7874;
assign a7880 = a7878 & a7772;
assign a7882 = ~a7880 & ~a7644;
assign a7884 = a7136 & ~l600;
assign a7886 = l604 & ~l602;
assign a7888 = a7886 & ~l600;
assign a7890 = ~l604 & l602;
assign a7892 = a7890 & ~l600;
assign a7894 = l604 & l602;
assign a7896 = a7894 & ~l600;
assign a7898 = a7136 & l600;
assign a7900 = ~l608 & ~l606;
assign a7902 = l608 & ~l606;
assign a7904 = ~l608 & l606;
assign a7906 = l608 & l606;
assign a7908 = a7906 & ~l1032;
assign a7910 = a7908 & ~a7904;
assign a7912 = a7904 & ~l1018;
assign a7914 = ~a7912 & ~a7910;
assign a7916 = ~a7914 & ~a7902;
assign a7918 = a7902 & ~l1004;
assign a7920 = ~a7918 & ~a7916;
assign a7922 = ~a7920 & ~a7900;
assign a7924 = a7900 & ~l990;
assign a7926 = ~a7924 & ~a7922;
assign a7928 = ~a7926 & a7898;
assign a7930 = a7928 & ~a7896;
assign a7932 = a7906 & ~l950;
assign a7934 = a7932 & ~a7904;
assign a7936 = a7904 & ~l936;
assign a7938 = ~a7936 & ~a7934;
assign a7940 = ~a7938 & ~a7902;
assign a7942 = a7902 & ~l922;
assign a7944 = ~a7942 & ~a7940;
assign a7946 = ~a7944 & ~a7900;
assign a7948 = a7900 & ~l908;
assign a7950 = ~a7948 & ~a7946;
assign a7952 = ~a7950 & a7896;
assign a7954 = ~a7952 & ~a7930;
assign a7956 = ~a7954 & ~a7892;
assign a7958 = a7906 & ~l868;
assign a7960 = a7958 & ~a7904;
assign a7962 = a7904 & ~l854;
assign a7964 = ~a7962 & ~a7960;
assign a7966 = ~a7964 & ~a7902;
assign a7968 = a7902 & ~l840;
assign a7970 = ~a7968 & ~a7966;
assign a7972 = ~a7970 & ~a7900;
assign a7974 = a7900 & ~l826;
assign a7976 = ~a7974 & ~a7972;
assign a7978 = ~a7976 & a7892;
assign a7980 = ~a7978 & ~a7956;
assign a7982 = ~a7980 & ~a7888;
assign a7984 = a7906 & ~l786;
assign a7986 = a7984 & ~a7904;
assign a7988 = a7904 & ~l772;
assign a7990 = ~a7988 & ~a7986;
assign a7992 = ~a7990 & ~a7902;
assign a7994 = a7902 & ~l758;
assign a7996 = ~a7994 & ~a7992;
assign a7998 = ~a7996 & ~a7900;
assign a8000 = a7900 & ~l744;
assign a8002 = ~a8000 & ~a7998;
assign a8004 = ~a8002 & a7888;
assign a8006 = ~a8004 & ~a7982;
assign a8008 = a8006 & ~l768;
assign a8010 = ~a8006 & l768;
assign a8012 = ~a8010 & ~a8008;
assign a8014 = a7906 & l1034;
assign a8016 = a8014 & ~a7904;
assign a8018 = a7904 & l1020;
assign a8020 = ~a8018 & ~a8016;
assign a8022 = ~a8020 & ~a7902;
assign a8024 = a7902 & l1006;
assign a8026 = ~a8024 & ~a8022;
assign a8028 = ~a8026 & ~a7900;
assign a8030 = a7900 & l992;
assign a8032 = ~a8030 & ~a8028;
assign a8034 = ~a8032 & a7898;
assign a8036 = a8034 & ~a7896;
assign a8038 = a7906 & l952;
assign a8040 = a8038 & ~a7904;
assign a8042 = a7904 & l938;
assign a8044 = ~a8042 & ~a8040;
assign a8046 = ~a8044 & ~a7902;
assign a8048 = a7902 & l924;
assign a8050 = ~a8048 & ~a8046;
assign a8052 = ~a8050 & ~a7900;
assign a8054 = a7900 & l910;
assign a8056 = ~a8054 & ~a8052;
assign a8058 = ~a8056 & a7896;
assign a8060 = ~a8058 & ~a8036;
assign a8062 = ~a8060 & ~a7892;
assign a8064 = a7906 & l870;
assign a8066 = a8064 & ~a7904;
assign a8068 = a7904 & l856;
assign a8070 = ~a8068 & ~a8066;
assign a8072 = ~a8070 & ~a7902;
assign a8074 = a7902 & l842;
assign a8076 = ~a8074 & ~a8072;
assign a8078 = ~a8076 & ~a7900;
assign a8080 = a7900 & l828;
assign a8082 = ~a8080 & ~a8078;
assign a8084 = ~a8082 & a7892;
assign a8086 = ~a8084 & ~a8062;
assign a8088 = ~a8086 & ~a7888;
assign a8090 = a7906 & l788;
assign a8092 = a8090 & ~a7904;
assign a8094 = a7904 & l774;
assign a8096 = ~a8094 & ~a8092;
assign a8098 = ~a8096 & ~a7902;
assign a8100 = a7902 & l760;
assign a8102 = ~a8100 & ~a8098;
assign a8104 = ~a8102 & ~a7900;
assign a8106 = a7900 & l746;
assign a8108 = ~a8106 & ~a8104;
assign a8110 = ~a8108 & a7888;
assign a8112 = ~a8110 & ~a8088;
assign a8114 = a8112 & ~l770;
assign a8116 = ~a8112 & l770;
assign a8118 = ~a8116 & ~a8114;
assign a8120 = a8118 & a8012;
assign a8122 = ~a8120 & ~a7884;
assign a8124 = a7140 & ~l610;
assign a8126 = l614 & ~l612;
assign a8128 = a8126 & ~l610;
assign a8130 = ~l614 & l612;
assign a8132 = a8130 & ~l610;
assign a8134 = l614 & l612;
assign a8136 = a8134 & ~l610;
assign a8138 = a7140 & l610;
assign a8140 = ~l618 & ~l616;
assign a8142 = l618 & ~l616;
assign a8144 = ~l618 & l616;
assign a8146 = l618 & l616;
assign a8148 = a8146 & ~l1032;
assign a8150 = a8148 & ~a8144;
assign a8152 = a8144 & ~l1018;
assign a8154 = ~a8152 & ~a8150;
assign a8156 = ~a8154 & ~a8142;
assign a8158 = a8142 & ~l1004;
assign a8160 = ~a8158 & ~a8156;
assign a8162 = ~a8160 & ~a8140;
assign a8164 = a8140 & ~l990;
assign a8166 = ~a8164 & ~a8162;
assign a8168 = ~a8166 & a8138;
assign a8170 = a8168 & ~a8136;
assign a8172 = a8146 & ~l950;
assign a8174 = a8172 & ~a8144;
assign a8176 = a8144 & ~l936;
assign a8178 = ~a8176 & ~a8174;
assign a8180 = ~a8178 & ~a8142;
assign a8182 = a8142 & ~l922;
assign a8184 = ~a8182 & ~a8180;
assign a8186 = ~a8184 & ~a8140;
assign a8188 = a8140 & ~l908;
assign a8190 = ~a8188 & ~a8186;
assign a8192 = ~a8190 & a8136;
assign a8194 = ~a8192 & ~a8170;
assign a8196 = ~a8194 & ~a8132;
assign a8198 = a8146 & ~l868;
assign a8200 = a8198 & ~a8144;
assign a8202 = a8144 & ~l854;
assign a8204 = ~a8202 & ~a8200;
assign a8206 = ~a8204 & ~a8142;
assign a8208 = a8142 & ~l840;
assign a8210 = ~a8208 & ~a8206;
assign a8212 = ~a8210 & ~a8140;
assign a8214 = a8140 & ~l826;
assign a8216 = ~a8214 & ~a8212;
assign a8218 = ~a8216 & a8132;
assign a8220 = ~a8218 & ~a8196;
assign a8222 = ~a8220 & ~a8128;
assign a8224 = a8146 & ~l786;
assign a8226 = a8224 & ~a8144;
assign a8228 = a8144 & ~l772;
assign a8230 = ~a8228 & ~a8226;
assign a8232 = ~a8230 & ~a8142;
assign a8234 = a8142 & ~l758;
assign a8236 = ~a8234 & ~a8232;
assign a8238 = ~a8236 & ~a8140;
assign a8240 = a8140 & ~l744;
assign a8242 = ~a8240 & ~a8238;
assign a8244 = ~a8242 & a8128;
assign a8246 = ~a8244 & ~a8222;
assign a8248 = a8246 & ~l782;
assign a8250 = ~a8246 & l782;
assign a8252 = ~a8250 & ~a8248;
assign a8254 = a8146 & l1034;
assign a8256 = a8254 & ~a8144;
assign a8258 = a8144 & l1020;
assign a8260 = ~a8258 & ~a8256;
assign a8262 = ~a8260 & ~a8142;
assign a8264 = a8142 & l1006;
assign a8266 = ~a8264 & ~a8262;
assign a8268 = ~a8266 & ~a8140;
assign a8270 = a8140 & l992;
assign a8272 = ~a8270 & ~a8268;
assign a8274 = ~a8272 & a8138;
assign a8276 = a8274 & ~a8136;
assign a8278 = a8146 & l952;
assign a8280 = a8278 & ~a8144;
assign a8282 = a8144 & l938;
assign a8284 = ~a8282 & ~a8280;
assign a8286 = ~a8284 & ~a8142;
assign a8288 = a8142 & l924;
assign a8290 = ~a8288 & ~a8286;
assign a8292 = ~a8290 & ~a8140;
assign a8294 = a8140 & l910;
assign a8296 = ~a8294 & ~a8292;
assign a8298 = ~a8296 & a8136;
assign a8300 = ~a8298 & ~a8276;
assign a8302 = ~a8300 & ~a8132;
assign a8304 = a8146 & l870;
assign a8306 = a8304 & ~a8144;
assign a8308 = a8144 & l856;
assign a8310 = ~a8308 & ~a8306;
assign a8312 = ~a8310 & ~a8142;
assign a8314 = a8142 & l842;
assign a8316 = ~a8314 & ~a8312;
assign a8318 = ~a8316 & ~a8140;
assign a8320 = a8140 & l828;
assign a8322 = ~a8320 & ~a8318;
assign a8324 = ~a8322 & a8132;
assign a8326 = ~a8324 & ~a8302;
assign a8328 = ~a8326 & ~a8128;
assign a8330 = a8146 & l788;
assign a8332 = a8330 & ~a8144;
assign a8334 = a8144 & l774;
assign a8336 = ~a8334 & ~a8332;
assign a8338 = ~a8336 & ~a8142;
assign a8340 = a8142 & l760;
assign a8342 = ~a8340 & ~a8338;
assign a8344 = ~a8342 & ~a8140;
assign a8346 = a8140 & l746;
assign a8348 = ~a8346 & ~a8344;
assign a8350 = ~a8348 & a8128;
assign a8352 = ~a8350 & ~a8328;
assign a8354 = a8352 & ~l784;
assign a8356 = ~a8352 & l784;
assign a8358 = ~a8356 & ~a8354;
assign a8360 = a8358 & a8252;
assign a8362 = ~a8360 & ~a8124;
assign a8364 = a7144 & ~l620;
assign a8366 = l624 & ~l622;
assign a8368 = a8366 & ~l620;
assign a8370 = ~l624 & l622;
assign a8372 = a8370 & ~l620;
assign a8374 = l624 & l622;
assign a8376 = a8374 & ~l620;
assign a8378 = a7144 & l620;
assign a8380 = ~l628 & ~l626;
assign a8382 = l628 & ~l626;
assign a8384 = ~l628 & l626;
assign a8386 = l628 & l626;
assign a8388 = a8386 & ~l1032;
assign a8390 = a8388 & ~a8384;
assign a8392 = a8384 & ~l1018;
assign a8394 = ~a8392 & ~a8390;
assign a8396 = ~a8394 & ~a8382;
assign a8398 = a8382 & ~l1004;
assign a8400 = ~a8398 & ~a8396;
assign a8402 = ~a8400 & ~a8380;
assign a8404 = a8380 & ~l990;
assign a8406 = ~a8404 & ~a8402;
assign a8408 = ~a8406 & a8378;
assign a8410 = a8408 & ~a8376;
assign a8412 = a8386 & ~l950;
assign a8414 = a8412 & ~a8384;
assign a8416 = a8384 & ~l936;
assign a8418 = ~a8416 & ~a8414;
assign a8420 = ~a8418 & ~a8382;
assign a8422 = a8382 & ~l922;
assign a8424 = ~a8422 & ~a8420;
assign a8426 = ~a8424 & ~a8380;
assign a8428 = a8380 & ~l908;
assign a8430 = ~a8428 & ~a8426;
assign a8432 = ~a8430 & a8376;
assign a8434 = ~a8432 & ~a8410;
assign a8436 = ~a8434 & ~a8372;
assign a8438 = a8386 & ~l868;
assign a8440 = a8438 & ~a8384;
assign a8442 = a8384 & ~l854;
assign a8444 = ~a8442 & ~a8440;
assign a8446 = ~a8444 & ~a8382;
assign a8448 = a8382 & ~l840;
assign a8450 = ~a8448 & ~a8446;
assign a8452 = ~a8450 & ~a8380;
assign a8454 = a8380 & ~l826;
assign a8456 = ~a8454 & ~a8452;
assign a8458 = ~a8456 & a8372;
assign a8460 = ~a8458 & ~a8436;
assign a8462 = ~a8460 & ~a8368;
assign a8464 = a8386 & ~l786;
assign a8466 = a8464 & ~a8384;
assign a8468 = a8384 & ~l772;
assign a8470 = ~a8468 & ~a8466;
assign a8472 = ~a8470 & ~a8382;
assign a8474 = a8382 & ~l758;
assign a8476 = ~a8474 & ~a8472;
assign a8478 = ~a8476 & ~a8380;
assign a8480 = a8380 & ~l744;
assign a8482 = ~a8480 & ~a8478;
assign a8484 = ~a8482 & a8368;
assign a8486 = ~a8484 & ~a8462;
assign a8488 = a8486 & ~l822;
assign a8490 = ~a8486 & l822;
assign a8492 = ~a8490 & ~a8488;
assign a8494 = a8386 & l1034;
assign a8496 = a8494 & ~a8384;
assign a8498 = a8384 & l1020;
assign a8500 = ~a8498 & ~a8496;
assign a8502 = ~a8500 & ~a8382;
assign a8504 = a8382 & l1006;
assign a8506 = ~a8504 & ~a8502;
assign a8508 = ~a8506 & ~a8380;
assign a8510 = a8380 & l992;
assign a8512 = ~a8510 & ~a8508;
assign a8514 = ~a8512 & a8378;
assign a8516 = a8514 & ~a8376;
assign a8518 = a8386 & l952;
assign a8520 = a8518 & ~a8384;
assign a8522 = a8384 & l938;
assign a8524 = ~a8522 & ~a8520;
assign a8526 = ~a8524 & ~a8382;
assign a8528 = a8382 & l924;
assign a8530 = ~a8528 & ~a8526;
assign a8532 = ~a8530 & ~a8380;
assign a8534 = a8380 & l910;
assign a8536 = ~a8534 & ~a8532;
assign a8538 = ~a8536 & a8376;
assign a8540 = ~a8538 & ~a8516;
assign a8542 = ~a8540 & ~a8372;
assign a8544 = a8386 & l870;
assign a8546 = a8544 & ~a8384;
assign a8548 = a8384 & l856;
assign a8550 = ~a8548 & ~a8546;
assign a8552 = ~a8550 & ~a8382;
assign a8554 = a8382 & l842;
assign a8556 = ~a8554 & ~a8552;
assign a8558 = ~a8556 & ~a8380;
assign a8560 = a8380 & l828;
assign a8562 = ~a8560 & ~a8558;
assign a8564 = ~a8562 & a8372;
assign a8566 = ~a8564 & ~a8542;
assign a8568 = ~a8566 & ~a8368;
assign a8570 = a8386 & l788;
assign a8572 = a8570 & ~a8384;
assign a8574 = a8384 & l774;
assign a8576 = ~a8574 & ~a8572;
assign a8578 = ~a8576 & ~a8382;
assign a8580 = a8382 & l760;
assign a8582 = ~a8580 & ~a8578;
assign a8584 = ~a8582 & ~a8380;
assign a8586 = a8380 & l746;
assign a8588 = ~a8586 & ~a8584;
assign a8590 = ~a8588 & a8368;
assign a8592 = ~a8590 & ~a8568;
assign a8594 = a8592 & ~l824;
assign a8596 = ~a8592 & l824;
assign a8598 = ~a8596 & ~a8594;
assign a8600 = a8598 & a8492;
assign a8602 = ~a8600 & ~a8364;
assign a8604 = a7148 & ~l630;
assign a8606 = l634 & ~l632;
assign a8608 = a8606 & ~l630;
assign a8610 = ~l634 & l632;
assign a8612 = a8610 & ~l630;
assign a8614 = l634 & l632;
assign a8616 = a8614 & ~l630;
assign a8618 = a7148 & l630;
assign a8620 = ~l638 & ~l636;
assign a8622 = l638 & ~l636;
assign a8624 = ~l638 & l636;
assign a8626 = l638 & l636;
assign a8628 = a8626 & ~l1032;
assign a8630 = a8628 & ~a8624;
assign a8632 = a8624 & ~l1018;
assign a8634 = ~a8632 & ~a8630;
assign a8636 = ~a8634 & ~a8622;
assign a8638 = a8622 & ~l1004;
assign a8640 = ~a8638 & ~a8636;
assign a8642 = ~a8640 & ~a8620;
assign a8644 = a8620 & ~l990;
assign a8646 = ~a8644 & ~a8642;
assign a8648 = ~a8646 & a8618;
assign a8650 = a8648 & ~a8616;
assign a8652 = a8626 & ~l950;
assign a8654 = a8652 & ~a8624;
assign a8656 = a8624 & ~l936;
assign a8658 = ~a8656 & ~a8654;
assign a8660 = ~a8658 & ~a8622;
assign a8662 = a8622 & ~l922;
assign a8664 = ~a8662 & ~a8660;
assign a8666 = ~a8664 & ~a8620;
assign a8668 = a8620 & ~l908;
assign a8670 = ~a8668 & ~a8666;
assign a8672 = ~a8670 & a8616;
assign a8674 = ~a8672 & ~a8650;
assign a8676 = ~a8674 & ~a8612;
assign a8678 = a8626 & ~l868;
assign a8680 = a8678 & ~a8624;
assign a8682 = a8624 & ~l854;
assign a8684 = ~a8682 & ~a8680;
assign a8686 = ~a8684 & ~a8622;
assign a8688 = a8622 & ~l840;
assign a8690 = ~a8688 & ~a8686;
assign a8692 = ~a8690 & ~a8620;
assign a8694 = a8620 & ~l826;
assign a8696 = ~a8694 & ~a8692;
assign a8698 = ~a8696 & a8612;
assign a8700 = ~a8698 & ~a8676;
assign a8702 = ~a8700 & ~a8608;
assign a8704 = a8626 & ~l786;
assign a8706 = a8704 & ~a8624;
assign a8708 = a8624 & ~l772;
assign a8710 = ~a8708 & ~a8706;
assign a8712 = ~a8710 & ~a8622;
assign a8714 = a8622 & ~l758;
assign a8716 = ~a8714 & ~a8712;
assign a8718 = ~a8716 & ~a8620;
assign a8720 = a8620 & ~l744;
assign a8722 = ~a8720 & ~a8718;
assign a8724 = ~a8722 & a8608;
assign a8726 = ~a8724 & ~a8702;
assign a8728 = a8726 & ~l836;
assign a8730 = ~a8726 & l836;
assign a8732 = ~a8730 & ~a8728;
assign a8734 = a8626 & l1034;
assign a8736 = a8734 & ~a8624;
assign a8738 = a8624 & l1020;
assign a8740 = ~a8738 & ~a8736;
assign a8742 = ~a8740 & ~a8622;
assign a8744 = a8622 & l1006;
assign a8746 = ~a8744 & ~a8742;
assign a8748 = ~a8746 & ~a8620;
assign a8750 = a8620 & l992;
assign a8752 = ~a8750 & ~a8748;
assign a8754 = ~a8752 & a8618;
assign a8756 = a8754 & ~a8616;
assign a8758 = a8626 & l952;
assign a8760 = a8758 & ~a8624;
assign a8762 = a8624 & l938;
assign a8764 = ~a8762 & ~a8760;
assign a8766 = ~a8764 & ~a8622;
assign a8768 = a8622 & l924;
assign a8770 = ~a8768 & ~a8766;
assign a8772 = ~a8770 & ~a8620;
assign a8774 = a8620 & l910;
assign a8776 = ~a8774 & ~a8772;
assign a8778 = ~a8776 & a8616;
assign a8780 = ~a8778 & ~a8756;
assign a8782 = ~a8780 & ~a8612;
assign a8784 = a8626 & l870;
assign a8786 = a8784 & ~a8624;
assign a8788 = a8624 & l856;
assign a8790 = ~a8788 & ~a8786;
assign a8792 = ~a8790 & ~a8622;
assign a8794 = a8622 & l842;
assign a8796 = ~a8794 & ~a8792;
assign a8798 = ~a8796 & ~a8620;
assign a8800 = a8620 & l828;
assign a8802 = ~a8800 & ~a8798;
assign a8804 = ~a8802 & a8612;
assign a8806 = ~a8804 & ~a8782;
assign a8808 = ~a8806 & ~a8608;
assign a8810 = a8626 & l788;
assign a8812 = a8810 & ~a8624;
assign a8814 = a8624 & l774;
assign a8816 = ~a8814 & ~a8812;
assign a8818 = ~a8816 & ~a8622;
assign a8820 = a8622 & l760;
assign a8822 = ~a8820 & ~a8818;
assign a8824 = ~a8822 & ~a8620;
assign a8826 = a8620 & l746;
assign a8828 = ~a8826 & ~a8824;
assign a8830 = ~a8828 & a8608;
assign a8832 = ~a8830 & ~a8808;
assign a8834 = a8832 & ~l838;
assign a8836 = ~a8832 & l838;
assign a8838 = ~a8836 & ~a8834;
assign a8840 = a8838 & a8732;
assign a8842 = ~a8840 & ~a8604;
assign a8844 = a7152 & ~l640;
assign a8846 = l644 & ~l642;
assign a8848 = a8846 & ~l640;
assign a8850 = ~l644 & l642;
assign a8852 = a8850 & ~l640;
assign a8854 = l644 & l642;
assign a8856 = a8854 & ~l640;
assign a8858 = a7152 & l640;
assign a8860 = ~l648 & ~l646;
assign a8862 = l648 & ~l646;
assign a8864 = ~l648 & l646;
assign a8866 = l648 & l646;
assign a8868 = a8866 & ~l1032;
assign a8870 = a8868 & ~a8864;
assign a8872 = a8864 & ~l1018;
assign a8874 = ~a8872 & ~a8870;
assign a8876 = ~a8874 & ~a8862;
assign a8878 = a8862 & ~l1004;
assign a8880 = ~a8878 & ~a8876;
assign a8882 = ~a8880 & ~a8860;
assign a8884 = a8860 & ~l990;
assign a8886 = ~a8884 & ~a8882;
assign a8888 = ~a8886 & a8858;
assign a8890 = a8888 & ~a8856;
assign a8892 = a8866 & ~l950;
assign a8894 = a8892 & ~a8864;
assign a8896 = a8864 & ~l936;
assign a8898 = ~a8896 & ~a8894;
assign a8900 = ~a8898 & ~a8862;
assign a8902 = a8862 & ~l922;
assign a8904 = ~a8902 & ~a8900;
assign a8906 = ~a8904 & ~a8860;
assign a8908 = a8860 & ~l908;
assign a8910 = ~a8908 & ~a8906;
assign a8912 = ~a8910 & a8856;
assign a8914 = ~a8912 & ~a8890;
assign a8916 = ~a8914 & ~a8852;
assign a8918 = a8866 & ~l868;
assign a8920 = a8918 & ~a8864;
assign a8922 = a8864 & ~l854;
assign a8924 = ~a8922 & ~a8920;
assign a8926 = ~a8924 & ~a8862;
assign a8928 = a8862 & ~l840;
assign a8930 = ~a8928 & ~a8926;
assign a8932 = ~a8930 & ~a8860;
assign a8934 = a8860 & ~l826;
assign a8936 = ~a8934 & ~a8932;
assign a8938 = ~a8936 & a8852;
assign a8940 = ~a8938 & ~a8916;
assign a8942 = ~a8940 & ~a8848;
assign a8944 = a8866 & ~l786;
assign a8946 = a8944 & ~a8864;
assign a8948 = a8864 & ~l772;
assign a8950 = ~a8948 & ~a8946;
assign a8952 = ~a8950 & ~a8862;
assign a8954 = a8862 & ~l758;
assign a8956 = ~a8954 & ~a8952;
assign a8958 = ~a8956 & ~a8860;
assign a8960 = a8860 & ~l744;
assign a8962 = ~a8960 & ~a8958;
assign a8964 = ~a8962 & a8848;
assign a8966 = ~a8964 & ~a8942;
assign a8968 = a8966 & ~l850;
assign a8970 = ~a8966 & l850;
assign a8972 = ~a8970 & ~a8968;
assign a8974 = a8866 & l1034;
assign a8976 = a8974 & ~a8864;
assign a8978 = a8864 & l1020;
assign a8980 = ~a8978 & ~a8976;
assign a8982 = ~a8980 & ~a8862;
assign a8984 = a8862 & l1006;
assign a8986 = ~a8984 & ~a8982;
assign a8988 = ~a8986 & ~a8860;
assign a8990 = a8860 & l992;
assign a8992 = ~a8990 & ~a8988;
assign a8994 = ~a8992 & a8858;
assign a8996 = a8994 & ~a8856;
assign a8998 = a8866 & l952;
assign a9000 = a8998 & ~a8864;
assign a9002 = a8864 & l938;
assign a9004 = ~a9002 & ~a9000;
assign a9006 = ~a9004 & ~a8862;
assign a9008 = a8862 & l924;
assign a9010 = ~a9008 & ~a9006;
assign a9012 = ~a9010 & ~a8860;
assign a9014 = a8860 & l910;
assign a9016 = ~a9014 & ~a9012;
assign a9018 = ~a9016 & a8856;
assign a9020 = ~a9018 & ~a8996;
assign a9022 = ~a9020 & ~a8852;
assign a9024 = a8866 & l870;
assign a9026 = a9024 & ~a8864;
assign a9028 = a8864 & l856;
assign a9030 = ~a9028 & ~a9026;
assign a9032 = ~a9030 & ~a8862;
assign a9034 = a8862 & l842;
assign a9036 = ~a9034 & ~a9032;
assign a9038 = ~a9036 & ~a8860;
assign a9040 = a8860 & l828;
assign a9042 = ~a9040 & ~a9038;
assign a9044 = ~a9042 & a8852;
assign a9046 = ~a9044 & ~a9022;
assign a9048 = ~a9046 & ~a8848;
assign a9050 = a8866 & l788;
assign a9052 = a9050 & ~a8864;
assign a9054 = a8864 & l774;
assign a9056 = ~a9054 & ~a9052;
assign a9058 = ~a9056 & ~a8862;
assign a9060 = a8862 & l760;
assign a9062 = ~a9060 & ~a9058;
assign a9064 = ~a9062 & ~a8860;
assign a9066 = a8860 & l746;
assign a9068 = ~a9066 & ~a9064;
assign a9070 = ~a9068 & a8848;
assign a9072 = ~a9070 & ~a9048;
assign a9074 = a9072 & ~l852;
assign a9076 = ~a9072 & l852;
assign a9078 = ~a9076 & ~a9074;
assign a9080 = a9078 & a8972;
assign a9082 = ~a9080 & ~a8844;
assign a9084 = a7156 & ~l650;
assign a9086 = l654 & ~l652;
assign a9088 = a9086 & ~l650;
assign a9090 = ~l654 & l652;
assign a9092 = a9090 & ~l650;
assign a9094 = l654 & l652;
assign a9096 = a9094 & ~l650;
assign a9098 = a7156 & l650;
assign a9100 = ~l658 & ~l656;
assign a9102 = l658 & ~l656;
assign a9104 = ~l658 & l656;
assign a9106 = l658 & l656;
assign a9108 = a9106 & ~l1032;
assign a9110 = a9108 & ~a9104;
assign a9112 = a9104 & ~l1018;
assign a9114 = ~a9112 & ~a9110;
assign a9116 = ~a9114 & ~a9102;
assign a9118 = a9102 & ~l1004;
assign a9120 = ~a9118 & ~a9116;
assign a9122 = ~a9120 & ~a9100;
assign a9124 = a9100 & ~l990;
assign a9126 = ~a9124 & ~a9122;
assign a9128 = ~a9126 & a9098;
assign a9130 = a9128 & ~a9096;
assign a9132 = a9106 & ~l950;
assign a9134 = a9132 & ~a9104;
assign a9136 = a9104 & ~l936;
assign a9138 = ~a9136 & ~a9134;
assign a9140 = ~a9138 & ~a9102;
assign a9142 = a9102 & ~l922;
assign a9144 = ~a9142 & ~a9140;
assign a9146 = ~a9144 & ~a9100;
assign a9148 = a9100 & ~l908;
assign a9150 = ~a9148 & ~a9146;
assign a9152 = ~a9150 & a9096;
assign a9154 = ~a9152 & ~a9130;
assign a9156 = ~a9154 & ~a9092;
assign a9158 = a9106 & ~l868;
assign a9160 = a9158 & ~a9104;
assign a9162 = a9104 & ~l854;
assign a9164 = ~a9162 & ~a9160;
assign a9166 = ~a9164 & ~a9102;
assign a9168 = a9102 & ~l840;
assign a9170 = ~a9168 & ~a9166;
assign a9172 = ~a9170 & ~a9100;
assign a9174 = a9100 & ~l826;
assign a9176 = ~a9174 & ~a9172;
assign a9178 = ~a9176 & a9092;
assign a9180 = ~a9178 & ~a9156;
assign a9182 = ~a9180 & ~a9088;
assign a9184 = a9106 & ~l786;
assign a9186 = a9184 & ~a9104;
assign a9188 = a9104 & ~l772;
assign a9190 = ~a9188 & ~a9186;
assign a9192 = ~a9190 & ~a9102;
assign a9194 = a9102 & ~l758;
assign a9196 = ~a9194 & ~a9192;
assign a9198 = ~a9196 & ~a9100;
assign a9200 = a9100 & ~l744;
assign a9202 = ~a9200 & ~a9198;
assign a9204 = ~a9202 & a9088;
assign a9206 = ~a9204 & ~a9182;
assign a9208 = a9206 & ~l864;
assign a9210 = ~a9206 & l864;
assign a9212 = ~a9210 & ~a9208;
assign a9214 = a9106 & l1034;
assign a9216 = a9214 & ~a9104;
assign a9218 = a9104 & l1020;
assign a9220 = ~a9218 & ~a9216;
assign a9222 = ~a9220 & ~a9102;
assign a9224 = a9102 & l1006;
assign a9226 = ~a9224 & ~a9222;
assign a9228 = ~a9226 & ~a9100;
assign a9230 = a9100 & l992;
assign a9232 = ~a9230 & ~a9228;
assign a9234 = ~a9232 & a9098;
assign a9236 = a9234 & ~a9096;
assign a9238 = a9106 & l952;
assign a9240 = a9238 & ~a9104;
assign a9242 = a9104 & l938;
assign a9244 = ~a9242 & ~a9240;
assign a9246 = ~a9244 & ~a9102;
assign a9248 = a9102 & l924;
assign a9250 = ~a9248 & ~a9246;
assign a9252 = ~a9250 & ~a9100;
assign a9254 = a9100 & l910;
assign a9256 = ~a9254 & ~a9252;
assign a9258 = ~a9256 & a9096;
assign a9260 = ~a9258 & ~a9236;
assign a9262 = ~a9260 & ~a9092;
assign a9264 = a9106 & l870;
assign a9266 = a9264 & ~a9104;
assign a9268 = a9104 & l856;
assign a9270 = ~a9268 & ~a9266;
assign a9272 = ~a9270 & ~a9102;
assign a9274 = a9102 & l842;
assign a9276 = ~a9274 & ~a9272;
assign a9278 = ~a9276 & ~a9100;
assign a9280 = a9100 & l828;
assign a9282 = ~a9280 & ~a9278;
assign a9284 = ~a9282 & a9092;
assign a9286 = ~a9284 & ~a9262;
assign a9288 = ~a9286 & ~a9088;
assign a9290 = a9106 & l788;
assign a9292 = a9290 & ~a9104;
assign a9294 = a9104 & l774;
assign a9296 = ~a9294 & ~a9292;
assign a9298 = ~a9296 & ~a9102;
assign a9300 = a9102 & l760;
assign a9302 = ~a9300 & ~a9298;
assign a9304 = ~a9302 & ~a9100;
assign a9306 = a9100 & l746;
assign a9308 = ~a9306 & ~a9304;
assign a9310 = ~a9308 & a9088;
assign a9312 = ~a9310 & ~a9288;
assign a9314 = a9312 & ~l866;
assign a9316 = ~a9312 & l866;
assign a9318 = ~a9316 & ~a9314;
assign a9320 = a9318 & a9212;
assign a9322 = ~a9320 & ~a9084;
assign a9324 = a7160 & ~l660;
assign a9326 = l664 & ~l662;
assign a9328 = a9326 & ~l660;
assign a9330 = ~l664 & l662;
assign a9332 = a9330 & ~l660;
assign a9334 = l664 & l662;
assign a9336 = a9334 & ~l660;
assign a9338 = a7160 & l660;
assign a9340 = ~l668 & ~l666;
assign a9342 = l668 & ~l666;
assign a9344 = ~l668 & l666;
assign a9346 = l668 & l666;
assign a9348 = a9346 & ~l1032;
assign a9350 = a9348 & ~a9344;
assign a9352 = a9344 & ~l1018;
assign a9354 = ~a9352 & ~a9350;
assign a9356 = ~a9354 & ~a9342;
assign a9358 = a9342 & ~l1004;
assign a9360 = ~a9358 & ~a9356;
assign a9362 = ~a9360 & ~a9340;
assign a9364 = a9340 & ~l990;
assign a9366 = ~a9364 & ~a9362;
assign a9368 = ~a9366 & a9338;
assign a9370 = a9368 & ~a9336;
assign a9372 = a9346 & ~l950;
assign a9374 = a9372 & ~a9344;
assign a9376 = a9344 & ~l936;
assign a9378 = ~a9376 & ~a9374;
assign a9380 = ~a9378 & ~a9342;
assign a9382 = a9342 & ~l922;
assign a9384 = ~a9382 & ~a9380;
assign a9386 = ~a9384 & ~a9340;
assign a9388 = a9340 & ~l908;
assign a9390 = ~a9388 & ~a9386;
assign a9392 = ~a9390 & a9336;
assign a9394 = ~a9392 & ~a9370;
assign a9396 = ~a9394 & ~a9332;
assign a9398 = a9346 & ~l868;
assign a9400 = a9398 & ~a9344;
assign a9402 = a9344 & ~l854;
assign a9404 = ~a9402 & ~a9400;
assign a9406 = ~a9404 & ~a9342;
assign a9408 = a9342 & ~l840;
assign a9410 = ~a9408 & ~a9406;
assign a9412 = ~a9410 & ~a9340;
assign a9414 = a9340 & ~l826;
assign a9416 = ~a9414 & ~a9412;
assign a9418 = ~a9416 & a9332;
assign a9420 = ~a9418 & ~a9396;
assign a9422 = ~a9420 & ~a9328;
assign a9424 = a9346 & ~l786;
assign a9426 = a9424 & ~a9344;
assign a9428 = a9344 & ~l772;
assign a9430 = ~a9428 & ~a9426;
assign a9432 = ~a9430 & ~a9342;
assign a9434 = a9342 & ~l758;
assign a9436 = ~a9434 & ~a9432;
assign a9438 = ~a9436 & ~a9340;
assign a9440 = a9340 & ~l744;
assign a9442 = ~a9440 & ~a9438;
assign a9444 = ~a9442 & a9328;
assign a9446 = ~a9444 & ~a9422;
assign a9448 = a9446 & ~l904;
assign a9450 = ~a9446 & l904;
assign a9452 = ~a9450 & ~a9448;
assign a9454 = a9346 & l1034;
assign a9456 = a9454 & ~a9344;
assign a9458 = a9344 & l1020;
assign a9460 = ~a9458 & ~a9456;
assign a9462 = ~a9460 & ~a9342;
assign a9464 = a9342 & l1006;
assign a9466 = ~a9464 & ~a9462;
assign a9468 = ~a9466 & ~a9340;
assign a9470 = a9340 & l992;
assign a9472 = ~a9470 & ~a9468;
assign a9474 = ~a9472 & a9338;
assign a9476 = a9474 & ~a9336;
assign a9478 = a9346 & l952;
assign a9480 = a9478 & ~a9344;
assign a9482 = a9344 & l938;
assign a9484 = ~a9482 & ~a9480;
assign a9486 = ~a9484 & ~a9342;
assign a9488 = a9342 & l924;
assign a9490 = ~a9488 & ~a9486;
assign a9492 = ~a9490 & ~a9340;
assign a9494 = a9340 & l910;
assign a9496 = ~a9494 & ~a9492;
assign a9498 = ~a9496 & a9336;
assign a9500 = ~a9498 & ~a9476;
assign a9502 = ~a9500 & ~a9332;
assign a9504 = a9346 & l870;
assign a9506 = a9504 & ~a9344;
assign a9508 = a9344 & l856;
assign a9510 = ~a9508 & ~a9506;
assign a9512 = ~a9510 & ~a9342;
assign a9514 = a9342 & l842;
assign a9516 = ~a9514 & ~a9512;
assign a9518 = ~a9516 & ~a9340;
assign a9520 = a9340 & l828;
assign a9522 = ~a9520 & ~a9518;
assign a9524 = ~a9522 & a9332;
assign a9526 = ~a9524 & ~a9502;
assign a9528 = ~a9526 & ~a9328;
assign a9530 = a9346 & l788;
assign a9532 = a9530 & ~a9344;
assign a9534 = a9344 & l774;
assign a9536 = ~a9534 & ~a9532;
assign a9538 = ~a9536 & ~a9342;
assign a9540 = a9342 & l760;
assign a9542 = ~a9540 & ~a9538;
assign a9544 = ~a9542 & ~a9340;
assign a9546 = a9340 & l746;
assign a9548 = ~a9546 & ~a9544;
assign a9550 = ~a9548 & a9328;
assign a9552 = ~a9550 & ~a9528;
assign a9554 = a9552 & ~l906;
assign a9556 = ~a9552 & l906;
assign a9558 = ~a9556 & ~a9554;
assign a9560 = a9558 & a9452;
assign a9562 = ~a9560 & ~a9324;
assign a9564 = a7164 & ~l670;
assign a9566 = l674 & ~l672;
assign a9568 = a9566 & ~l670;
assign a9570 = ~l674 & l672;
assign a9572 = a9570 & ~l670;
assign a9574 = l674 & l672;
assign a9576 = a9574 & ~l670;
assign a9578 = a7164 & l670;
assign a9580 = ~l678 & ~l676;
assign a9582 = l678 & ~l676;
assign a9584 = ~l678 & l676;
assign a9586 = l678 & l676;
assign a9588 = a9586 & ~l1032;
assign a9590 = a9588 & ~a9584;
assign a9592 = a9584 & ~l1018;
assign a9594 = ~a9592 & ~a9590;
assign a9596 = ~a9594 & ~a9582;
assign a9598 = a9582 & ~l1004;
assign a9600 = ~a9598 & ~a9596;
assign a9602 = ~a9600 & ~a9580;
assign a9604 = a9580 & ~l990;
assign a9606 = ~a9604 & ~a9602;
assign a9608 = ~a9606 & a9578;
assign a9610 = a9608 & ~a9576;
assign a9612 = a9586 & ~l950;
assign a9614 = a9612 & ~a9584;
assign a9616 = a9584 & ~l936;
assign a9618 = ~a9616 & ~a9614;
assign a9620 = ~a9618 & ~a9582;
assign a9622 = a9582 & ~l922;
assign a9624 = ~a9622 & ~a9620;
assign a9626 = ~a9624 & ~a9580;
assign a9628 = a9580 & ~l908;
assign a9630 = ~a9628 & ~a9626;
assign a9632 = ~a9630 & a9576;
assign a9634 = ~a9632 & ~a9610;
assign a9636 = ~a9634 & ~a9572;
assign a9638 = a9586 & ~l868;
assign a9640 = a9638 & ~a9584;
assign a9642 = a9584 & ~l854;
assign a9644 = ~a9642 & ~a9640;
assign a9646 = ~a9644 & ~a9582;
assign a9648 = a9582 & ~l840;
assign a9650 = ~a9648 & ~a9646;
assign a9652 = ~a9650 & ~a9580;
assign a9654 = a9580 & ~l826;
assign a9656 = ~a9654 & ~a9652;
assign a9658 = ~a9656 & a9572;
assign a9660 = ~a9658 & ~a9636;
assign a9662 = ~a9660 & ~a9568;
assign a9664 = a9586 & ~l786;
assign a9666 = a9664 & ~a9584;
assign a9668 = a9584 & ~l772;
assign a9670 = ~a9668 & ~a9666;
assign a9672 = ~a9670 & ~a9582;
assign a9674 = a9582 & ~l758;
assign a9676 = ~a9674 & ~a9672;
assign a9678 = ~a9676 & ~a9580;
assign a9680 = a9580 & ~l744;
assign a9682 = ~a9680 & ~a9678;
assign a9684 = ~a9682 & a9568;
assign a9686 = ~a9684 & ~a9662;
assign a9688 = a9686 & ~l918;
assign a9690 = ~a9686 & l918;
assign a9692 = ~a9690 & ~a9688;
assign a9694 = a9586 & l1034;
assign a9696 = a9694 & ~a9584;
assign a9698 = a9584 & l1020;
assign a9700 = ~a9698 & ~a9696;
assign a9702 = ~a9700 & ~a9582;
assign a9704 = a9582 & l1006;
assign a9706 = ~a9704 & ~a9702;
assign a9708 = ~a9706 & ~a9580;
assign a9710 = a9580 & l992;
assign a9712 = ~a9710 & ~a9708;
assign a9714 = ~a9712 & a9578;
assign a9716 = a9714 & ~a9576;
assign a9718 = a9586 & l952;
assign a9720 = a9718 & ~a9584;
assign a9722 = a9584 & l938;
assign a9724 = ~a9722 & ~a9720;
assign a9726 = ~a9724 & ~a9582;
assign a9728 = a9582 & l924;
assign a9730 = ~a9728 & ~a9726;
assign a9732 = ~a9730 & ~a9580;
assign a9734 = a9580 & l910;
assign a9736 = ~a9734 & ~a9732;
assign a9738 = ~a9736 & a9576;
assign a9740 = ~a9738 & ~a9716;
assign a9742 = ~a9740 & ~a9572;
assign a9744 = a9586 & l870;
assign a9746 = a9744 & ~a9584;
assign a9748 = a9584 & l856;
assign a9750 = ~a9748 & ~a9746;
assign a9752 = ~a9750 & ~a9582;
assign a9754 = a9582 & l842;
assign a9756 = ~a9754 & ~a9752;
assign a9758 = ~a9756 & ~a9580;
assign a9760 = a9580 & l828;
assign a9762 = ~a9760 & ~a9758;
assign a9764 = ~a9762 & a9572;
assign a9766 = ~a9764 & ~a9742;
assign a9768 = ~a9766 & ~a9568;
assign a9770 = a9586 & l788;
assign a9772 = a9770 & ~a9584;
assign a9774 = a9584 & l774;
assign a9776 = ~a9774 & ~a9772;
assign a9778 = ~a9776 & ~a9582;
assign a9780 = a9582 & l760;
assign a9782 = ~a9780 & ~a9778;
assign a9784 = ~a9782 & ~a9580;
assign a9786 = a9580 & l746;
assign a9788 = ~a9786 & ~a9784;
assign a9790 = ~a9788 & a9568;
assign a9792 = ~a9790 & ~a9768;
assign a9794 = a9792 & ~l920;
assign a9796 = ~a9792 & l920;
assign a9798 = ~a9796 & ~a9794;
assign a9800 = a9798 & a9692;
assign a9802 = ~a9800 & ~a9564;
assign a9804 = a7168 & ~l680;
assign a9806 = l684 & ~l682;
assign a9808 = a9806 & ~l680;
assign a9810 = ~l684 & l682;
assign a9812 = a9810 & ~l680;
assign a9814 = l684 & l682;
assign a9816 = a9814 & ~l680;
assign a9818 = a7168 & l680;
assign a9820 = ~l688 & ~l686;
assign a9822 = l688 & ~l686;
assign a9824 = ~l688 & l686;
assign a9826 = l688 & l686;
assign a9828 = a9826 & ~l1032;
assign a9830 = a9828 & ~a9824;
assign a9832 = a9824 & ~l1018;
assign a9834 = ~a9832 & ~a9830;
assign a9836 = ~a9834 & ~a9822;
assign a9838 = a9822 & ~l1004;
assign a9840 = ~a9838 & ~a9836;
assign a9842 = ~a9840 & ~a9820;
assign a9844 = a9820 & ~l990;
assign a9846 = ~a9844 & ~a9842;
assign a9848 = ~a9846 & a9818;
assign a9850 = a9848 & ~a9816;
assign a9852 = a9826 & ~l950;
assign a9854 = a9852 & ~a9824;
assign a9856 = a9824 & ~l936;
assign a9858 = ~a9856 & ~a9854;
assign a9860 = ~a9858 & ~a9822;
assign a9862 = a9822 & ~l922;
assign a9864 = ~a9862 & ~a9860;
assign a9866 = ~a9864 & ~a9820;
assign a9868 = a9820 & ~l908;
assign a9870 = ~a9868 & ~a9866;
assign a9872 = ~a9870 & a9816;
assign a9874 = ~a9872 & ~a9850;
assign a9876 = ~a9874 & ~a9812;
assign a9878 = a9826 & ~l868;
assign a9880 = a9878 & ~a9824;
assign a9882 = a9824 & ~l854;
assign a9884 = ~a9882 & ~a9880;
assign a9886 = ~a9884 & ~a9822;
assign a9888 = a9822 & ~l840;
assign a9890 = ~a9888 & ~a9886;
assign a9892 = ~a9890 & ~a9820;
assign a9894 = a9820 & ~l826;
assign a9896 = ~a9894 & ~a9892;
assign a9898 = ~a9896 & a9812;
assign a9900 = ~a9898 & ~a9876;
assign a9902 = ~a9900 & ~a9808;
assign a9904 = a9826 & ~l786;
assign a9906 = a9904 & ~a9824;
assign a9908 = a9824 & ~l772;
assign a9910 = ~a9908 & ~a9906;
assign a9912 = ~a9910 & ~a9822;
assign a9914 = a9822 & ~l758;
assign a9916 = ~a9914 & ~a9912;
assign a9918 = ~a9916 & ~a9820;
assign a9920 = a9820 & ~l744;
assign a9922 = ~a9920 & ~a9918;
assign a9924 = ~a9922 & a9808;
assign a9926 = ~a9924 & ~a9902;
assign a9928 = a9926 & ~l932;
assign a9930 = ~a9926 & l932;
assign a9932 = ~a9930 & ~a9928;
assign a9934 = a9826 & l1034;
assign a9936 = a9934 & ~a9824;
assign a9938 = a9824 & l1020;
assign a9940 = ~a9938 & ~a9936;
assign a9942 = ~a9940 & ~a9822;
assign a9944 = a9822 & l1006;
assign a9946 = ~a9944 & ~a9942;
assign a9948 = ~a9946 & ~a9820;
assign a9950 = a9820 & l992;
assign a9952 = ~a9950 & ~a9948;
assign a9954 = ~a9952 & a9818;
assign a9956 = a9954 & ~a9816;
assign a9958 = a9826 & l952;
assign a9960 = a9958 & ~a9824;
assign a9962 = a9824 & l938;
assign a9964 = ~a9962 & ~a9960;
assign a9966 = ~a9964 & ~a9822;
assign a9968 = a9822 & l924;
assign a9970 = ~a9968 & ~a9966;
assign a9972 = ~a9970 & ~a9820;
assign a9974 = a9820 & l910;
assign a9976 = ~a9974 & ~a9972;
assign a9978 = ~a9976 & a9816;
assign a9980 = ~a9978 & ~a9956;
assign a9982 = ~a9980 & ~a9812;
assign a9984 = a9826 & l870;
assign a9986 = a9984 & ~a9824;
assign a9988 = a9824 & l856;
assign a9990 = ~a9988 & ~a9986;
assign a9992 = ~a9990 & ~a9822;
assign a9994 = a9822 & l842;
assign a9996 = ~a9994 & ~a9992;
assign a9998 = ~a9996 & ~a9820;
assign a10000 = a9820 & l828;
assign a10002 = ~a10000 & ~a9998;
assign a10004 = ~a10002 & a9812;
assign a10006 = ~a10004 & ~a9982;
assign a10008 = ~a10006 & ~a9808;
assign a10010 = a9826 & l788;
assign a10012 = a10010 & ~a9824;
assign a10014 = a9824 & l774;
assign a10016 = ~a10014 & ~a10012;
assign a10018 = ~a10016 & ~a9822;
assign a10020 = a9822 & l760;
assign a10022 = ~a10020 & ~a10018;
assign a10024 = ~a10022 & ~a9820;
assign a10026 = a9820 & l746;
assign a10028 = ~a10026 & ~a10024;
assign a10030 = ~a10028 & a9808;
assign a10032 = ~a10030 & ~a10008;
assign a10034 = a10032 & ~l934;
assign a10036 = ~a10032 & l934;
assign a10038 = ~a10036 & ~a10034;
assign a10040 = a10038 & a9932;
assign a10042 = ~a10040 & ~a9804;
assign a10044 = a7172 & ~l690;
assign a10046 = l694 & ~l692;
assign a10048 = a10046 & ~l690;
assign a10050 = ~l694 & l692;
assign a10052 = a10050 & ~l690;
assign a10054 = l694 & l692;
assign a10056 = a10054 & ~l690;
assign a10058 = a7172 & l690;
assign a10060 = ~l698 & ~l696;
assign a10062 = l698 & ~l696;
assign a10064 = ~l698 & l696;
assign a10066 = l698 & l696;
assign a10068 = a10066 & ~l1032;
assign a10070 = a10068 & ~a10064;
assign a10072 = a10064 & ~l1018;
assign a10074 = ~a10072 & ~a10070;
assign a10076 = ~a10074 & ~a10062;
assign a10078 = a10062 & ~l1004;
assign a10080 = ~a10078 & ~a10076;
assign a10082 = ~a10080 & ~a10060;
assign a10084 = a10060 & ~l990;
assign a10086 = ~a10084 & ~a10082;
assign a10088 = ~a10086 & a10058;
assign a10090 = a10088 & ~a10056;
assign a10092 = a10066 & ~l950;
assign a10094 = a10092 & ~a10064;
assign a10096 = a10064 & ~l936;
assign a10098 = ~a10096 & ~a10094;
assign a10100 = ~a10098 & ~a10062;
assign a10102 = a10062 & ~l922;
assign a10104 = ~a10102 & ~a10100;
assign a10106 = ~a10104 & ~a10060;
assign a10108 = a10060 & ~l908;
assign a10110 = ~a10108 & ~a10106;
assign a10112 = ~a10110 & a10056;
assign a10114 = ~a10112 & ~a10090;
assign a10116 = ~a10114 & ~a10052;
assign a10118 = a10066 & ~l868;
assign a10120 = a10118 & ~a10064;
assign a10122 = a10064 & ~l854;
assign a10124 = ~a10122 & ~a10120;
assign a10126 = ~a10124 & ~a10062;
assign a10128 = a10062 & ~l840;
assign a10130 = ~a10128 & ~a10126;
assign a10132 = ~a10130 & ~a10060;
assign a10134 = a10060 & ~l826;
assign a10136 = ~a10134 & ~a10132;
assign a10138 = ~a10136 & a10052;
assign a10140 = ~a10138 & ~a10116;
assign a10142 = ~a10140 & ~a10048;
assign a10144 = a10066 & ~l786;
assign a10146 = a10144 & ~a10064;
assign a10148 = a10064 & ~l772;
assign a10150 = ~a10148 & ~a10146;
assign a10152 = ~a10150 & ~a10062;
assign a10154 = a10062 & ~l758;
assign a10156 = ~a10154 & ~a10152;
assign a10158 = ~a10156 & ~a10060;
assign a10160 = a10060 & ~l744;
assign a10162 = ~a10160 & ~a10158;
assign a10164 = ~a10162 & a10048;
assign a10166 = ~a10164 & ~a10142;
assign a10168 = a10166 & ~l946;
assign a10170 = ~a10166 & l946;
assign a10172 = ~a10170 & ~a10168;
assign a10174 = a10066 & l1034;
assign a10176 = a10174 & ~a10064;
assign a10178 = a10064 & l1020;
assign a10180 = ~a10178 & ~a10176;
assign a10182 = ~a10180 & ~a10062;
assign a10184 = a10062 & l1006;
assign a10186 = ~a10184 & ~a10182;
assign a10188 = ~a10186 & ~a10060;
assign a10190 = a10060 & l992;
assign a10192 = ~a10190 & ~a10188;
assign a10194 = ~a10192 & a10058;
assign a10196 = a10194 & ~a10056;
assign a10198 = a10066 & l952;
assign a10200 = a10198 & ~a10064;
assign a10202 = a10064 & l938;
assign a10204 = ~a10202 & ~a10200;
assign a10206 = ~a10204 & ~a10062;
assign a10208 = a10062 & l924;
assign a10210 = ~a10208 & ~a10206;
assign a10212 = ~a10210 & ~a10060;
assign a10214 = a10060 & l910;
assign a10216 = ~a10214 & ~a10212;
assign a10218 = ~a10216 & a10056;
assign a10220 = ~a10218 & ~a10196;
assign a10222 = ~a10220 & ~a10052;
assign a10224 = a10066 & l870;
assign a10226 = a10224 & ~a10064;
assign a10228 = a10064 & l856;
assign a10230 = ~a10228 & ~a10226;
assign a10232 = ~a10230 & ~a10062;
assign a10234 = a10062 & l842;
assign a10236 = ~a10234 & ~a10232;
assign a10238 = ~a10236 & ~a10060;
assign a10240 = a10060 & l828;
assign a10242 = ~a10240 & ~a10238;
assign a10244 = ~a10242 & a10052;
assign a10246 = ~a10244 & ~a10222;
assign a10248 = ~a10246 & ~a10048;
assign a10250 = a10066 & l788;
assign a10252 = a10250 & ~a10064;
assign a10254 = a10064 & l774;
assign a10256 = ~a10254 & ~a10252;
assign a10258 = ~a10256 & ~a10062;
assign a10260 = a10062 & l760;
assign a10262 = ~a10260 & ~a10258;
assign a10264 = ~a10262 & ~a10060;
assign a10266 = a10060 & l746;
assign a10268 = ~a10266 & ~a10264;
assign a10270 = ~a10268 & a10048;
assign a10272 = ~a10270 & ~a10248;
assign a10274 = a10272 & ~l948;
assign a10276 = ~a10272 & l948;
assign a10278 = ~a10276 & ~a10274;
assign a10280 = a10278 & a10172;
assign a10282 = ~a10280 & ~a10044;
assign a10284 = a7176 & ~l700;
assign a10286 = l704 & ~l702;
assign a10288 = a10286 & ~l700;
assign a10290 = ~l704 & l702;
assign a10292 = a10290 & ~l700;
assign a10294 = l704 & l702;
assign a10296 = a10294 & ~l700;
assign a10298 = a7176 & l700;
assign a10300 = ~l708 & ~l706;
assign a10302 = l708 & ~l706;
assign a10304 = ~l708 & l706;
assign a10306 = l708 & l706;
assign a10308 = a10306 & ~l1032;
assign a10310 = a10308 & ~a10304;
assign a10312 = a10304 & ~l1018;
assign a10314 = ~a10312 & ~a10310;
assign a10316 = ~a10314 & ~a10302;
assign a10318 = a10302 & ~l1004;
assign a10320 = ~a10318 & ~a10316;
assign a10322 = ~a10320 & ~a10300;
assign a10324 = a10300 & ~l990;
assign a10326 = ~a10324 & ~a10322;
assign a10328 = ~a10326 & a10298;
assign a10330 = a10328 & ~a10296;
assign a10332 = a10306 & ~l950;
assign a10334 = a10332 & ~a10304;
assign a10336 = a10304 & ~l936;
assign a10338 = ~a10336 & ~a10334;
assign a10340 = ~a10338 & ~a10302;
assign a10342 = a10302 & ~l922;
assign a10344 = ~a10342 & ~a10340;
assign a10346 = ~a10344 & ~a10300;
assign a10348 = a10300 & ~l908;
assign a10350 = ~a10348 & ~a10346;
assign a10352 = ~a10350 & a10296;
assign a10354 = ~a10352 & ~a10330;
assign a10356 = ~a10354 & ~a10292;
assign a10358 = a10306 & ~l868;
assign a10360 = a10358 & ~a10304;
assign a10362 = a10304 & ~l854;
assign a10364 = ~a10362 & ~a10360;
assign a10366 = ~a10364 & ~a10302;
assign a10368 = a10302 & ~l840;
assign a10370 = ~a10368 & ~a10366;
assign a10372 = ~a10370 & ~a10300;
assign a10374 = a10300 & ~l826;
assign a10376 = ~a10374 & ~a10372;
assign a10378 = ~a10376 & a10292;
assign a10380 = ~a10378 & ~a10356;
assign a10382 = ~a10380 & ~a10288;
assign a10384 = a10306 & ~l786;
assign a10386 = a10384 & ~a10304;
assign a10388 = a10304 & ~l772;
assign a10390 = ~a10388 & ~a10386;
assign a10392 = ~a10390 & ~a10302;
assign a10394 = a10302 & ~l758;
assign a10396 = ~a10394 & ~a10392;
assign a10398 = ~a10396 & ~a10300;
assign a10400 = a10300 & ~l744;
assign a10402 = ~a10400 & ~a10398;
assign a10404 = ~a10402 & a10288;
assign a10406 = ~a10404 & ~a10382;
assign a10408 = a10406 & ~l986;
assign a10410 = ~a10406 & l986;
assign a10412 = ~a10410 & ~a10408;
assign a10414 = a10306 & l1034;
assign a10416 = a10414 & ~a10304;
assign a10418 = a10304 & l1020;
assign a10420 = ~a10418 & ~a10416;
assign a10422 = ~a10420 & ~a10302;
assign a10424 = a10302 & l1006;
assign a10426 = ~a10424 & ~a10422;
assign a10428 = ~a10426 & ~a10300;
assign a10430 = a10300 & l992;
assign a10432 = ~a10430 & ~a10428;
assign a10434 = ~a10432 & a10298;
assign a10436 = a10434 & ~a10296;
assign a10438 = a10306 & l952;
assign a10440 = a10438 & ~a10304;
assign a10442 = a10304 & l938;
assign a10444 = ~a10442 & ~a10440;
assign a10446 = ~a10444 & ~a10302;
assign a10448 = a10302 & l924;
assign a10450 = ~a10448 & ~a10446;
assign a10452 = ~a10450 & ~a10300;
assign a10454 = a10300 & l910;
assign a10456 = ~a10454 & ~a10452;
assign a10458 = ~a10456 & a10296;
assign a10460 = ~a10458 & ~a10436;
assign a10462 = ~a10460 & ~a10292;
assign a10464 = a10306 & l870;
assign a10466 = a10464 & ~a10304;
assign a10468 = a10304 & l856;
assign a10470 = ~a10468 & ~a10466;
assign a10472 = ~a10470 & ~a10302;
assign a10474 = a10302 & l842;
assign a10476 = ~a10474 & ~a10472;
assign a10478 = ~a10476 & ~a10300;
assign a10480 = a10300 & l828;
assign a10482 = ~a10480 & ~a10478;
assign a10484 = ~a10482 & a10292;
assign a10486 = ~a10484 & ~a10462;
assign a10488 = ~a10486 & ~a10288;
assign a10490 = a10306 & l788;
assign a10492 = a10490 & ~a10304;
assign a10494 = a10304 & l774;
assign a10496 = ~a10494 & ~a10492;
assign a10498 = ~a10496 & ~a10302;
assign a10500 = a10302 & l760;
assign a10502 = ~a10500 & ~a10498;
assign a10504 = ~a10502 & ~a10300;
assign a10506 = a10300 & l746;
assign a10508 = ~a10506 & ~a10504;
assign a10510 = ~a10508 & a10288;
assign a10512 = ~a10510 & ~a10488;
assign a10514 = a10512 & ~l988;
assign a10516 = ~a10512 & l988;
assign a10518 = ~a10516 & ~a10514;
assign a10520 = a10518 & a10412;
assign a10522 = ~a10520 & ~a10284;
assign a10524 = a7180 & ~l710;
assign a10526 = l714 & ~l712;
assign a10528 = a10526 & ~l710;
assign a10530 = ~l714 & l712;
assign a10532 = a10530 & ~l710;
assign a10534 = l714 & l712;
assign a10536 = a10534 & ~l710;
assign a10538 = a7180 & l710;
assign a10540 = ~l718 & ~l716;
assign a10542 = l718 & ~l716;
assign a10544 = ~l718 & l716;
assign a10546 = l718 & l716;
assign a10548 = a10546 & ~l1032;
assign a10550 = a10548 & ~a10544;
assign a10552 = a10544 & ~l1018;
assign a10554 = ~a10552 & ~a10550;
assign a10556 = ~a10554 & ~a10542;
assign a10558 = a10542 & ~l1004;
assign a10560 = ~a10558 & ~a10556;
assign a10562 = ~a10560 & ~a10540;
assign a10564 = a10540 & ~l990;
assign a10566 = ~a10564 & ~a10562;
assign a10568 = ~a10566 & a10538;
assign a10570 = a10568 & ~a10536;
assign a10572 = a10546 & ~l950;
assign a10574 = a10572 & ~a10544;
assign a10576 = a10544 & ~l936;
assign a10578 = ~a10576 & ~a10574;
assign a10580 = ~a10578 & ~a10542;
assign a10582 = a10542 & ~l922;
assign a10584 = ~a10582 & ~a10580;
assign a10586 = ~a10584 & ~a10540;
assign a10588 = a10540 & ~l908;
assign a10590 = ~a10588 & ~a10586;
assign a10592 = ~a10590 & a10536;
assign a10594 = ~a10592 & ~a10570;
assign a10596 = ~a10594 & ~a10532;
assign a10598 = a10546 & ~l868;
assign a10600 = a10598 & ~a10544;
assign a10602 = a10544 & ~l854;
assign a10604 = ~a10602 & ~a10600;
assign a10606 = ~a10604 & ~a10542;
assign a10608 = a10542 & ~l840;
assign a10610 = ~a10608 & ~a10606;
assign a10612 = ~a10610 & ~a10540;
assign a10614 = a10540 & ~l826;
assign a10616 = ~a10614 & ~a10612;
assign a10618 = ~a10616 & a10532;
assign a10620 = ~a10618 & ~a10596;
assign a10622 = ~a10620 & ~a10528;
assign a10624 = a10546 & ~l786;
assign a10626 = a10624 & ~a10544;
assign a10628 = a10544 & ~l772;
assign a10630 = ~a10628 & ~a10626;
assign a10632 = ~a10630 & ~a10542;
assign a10634 = a10542 & ~l758;
assign a10636 = ~a10634 & ~a10632;
assign a10638 = ~a10636 & ~a10540;
assign a10640 = a10540 & ~l744;
assign a10642 = ~a10640 & ~a10638;
assign a10644 = ~a10642 & a10528;
assign a10646 = ~a10644 & ~a10622;
assign a10648 = a10646 & ~l1000;
assign a10650 = ~a10646 & l1000;
assign a10652 = ~a10650 & ~a10648;
assign a10654 = a10546 & l1034;
assign a10656 = a10654 & ~a10544;
assign a10658 = a10544 & l1020;
assign a10660 = ~a10658 & ~a10656;
assign a10662 = ~a10660 & ~a10542;
assign a10664 = a10542 & l1006;
assign a10666 = ~a10664 & ~a10662;
assign a10668 = ~a10666 & ~a10540;
assign a10670 = a10540 & l992;
assign a10672 = ~a10670 & ~a10668;
assign a10674 = ~a10672 & a10538;
assign a10676 = a10674 & ~a10536;
assign a10678 = a10546 & l952;
assign a10680 = a10678 & ~a10544;
assign a10682 = a10544 & l938;
assign a10684 = ~a10682 & ~a10680;
assign a10686 = ~a10684 & ~a10542;
assign a10688 = a10542 & l924;
assign a10690 = ~a10688 & ~a10686;
assign a10692 = ~a10690 & ~a10540;
assign a10694 = a10540 & l910;
assign a10696 = ~a10694 & ~a10692;
assign a10698 = ~a10696 & a10536;
assign a10700 = ~a10698 & ~a10676;
assign a10702 = ~a10700 & ~a10532;
assign a10704 = a10546 & l870;
assign a10706 = a10704 & ~a10544;
assign a10708 = a10544 & l856;
assign a10710 = ~a10708 & ~a10706;
assign a10712 = ~a10710 & ~a10542;
assign a10714 = a10542 & l842;
assign a10716 = ~a10714 & ~a10712;
assign a10718 = ~a10716 & ~a10540;
assign a10720 = a10540 & l828;
assign a10722 = ~a10720 & ~a10718;
assign a10724 = ~a10722 & a10532;
assign a10726 = ~a10724 & ~a10702;
assign a10728 = ~a10726 & ~a10528;
assign a10730 = a10546 & l788;
assign a10732 = a10730 & ~a10544;
assign a10734 = a10544 & l774;
assign a10736 = ~a10734 & ~a10732;
assign a10738 = ~a10736 & ~a10542;
assign a10740 = a10542 & l760;
assign a10742 = ~a10740 & ~a10738;
assign a10744 = ~a10742 & ~a10540;
assign a10746 = a10540 & l746;
assign a10748 = ~a10746 & ~a10744;
assign a10750 = ~a10748 & a10528;
assign a10752 = ~a10750 & ~a10728;
assign a10754 = a10752 & ~l1002;
assign a10756 = ~a10752 & l1002;
assign a10758 = ~a10756 & ~a10754;
assign a10760 = a10758 & a10652;
assign a10762 = ~a10760 & ~a10524;
assign a10764 = a7184 & ~l720;
assign a10766 = l724 & ~l722;
assign a10768 = a10766 & ~l720;
assign a10770 = ~l724 & l722;
assign a10772 = a10770 & ~l720;
assign a10774 = l724 & l722;
assign a10776 = a10774 & ~l720;
assign a10778 = a7184 & l720;
assign a10780 = ~l728 & ~l726;
assign a10782 = l728 & ~l726;
assign a10784 = ~l728 & l726;
assign a10786 = l728 & l726;
assign a10788 = a10786 & ~l1032;
assign a10790 = a10788 & ~a10784;
assign a10792 = a10784 & ~l1018;
assign a10794 = ~a10792 & ~a10790;
assign a10796 = ~a10794 & ~a10782;
assign a10798 = a10782 & ~l1004;
assign a10800 = ~a10798 & ~a10796;
assign a10802 = ~a10800 & ~a10780;
assign a10804 = a10780 & ~l990;
assign a10806 = ~a10804 & ~a10802;
assign a10808 = ~a10806 & a10778;
assign a10810 = a10808 & ~a10776;
assign a10812 = a10786 & ~l950;
assign a10814 = a10812 & ~a10784;
assign a10816 = a10784 & ~l936;
assign a10818 = ~a10816 & ~a10814;
assign a10820 = ~a10818 & ~a10782;
assign a10822 = a10782 & ~l922;
assign a10824 = ~a10822 & ~a10820;
assign a10826 = ~a10824 & ~a10780;
assign a10828 = a10780 & ~l908;
assign a10830 = ~a10828 & ~a10826;
assign a10832 = ~a10830 & a10776;
assign a10834 = ~a10832 & ~a10810;
assign a10836 = ~a10834 & ~a10772;
assign a10838 = a10786 & ~l868;
assign a10840 = a10838 & ~a10784;
assign a10842 = a10784 & ~l854;
assign a10844 = ~a10842 & ~a10840;
assign a10846 = ~a10844 & ~a10782;
assign a10848 = a10782 & ~l840;
assign a10850 = ~a10848 & ~a10846;
assign a10852 = ~a10850 & ~a10780;
assign a10854 = a10780 & ~l826;
assign a10856 = ~a10854 & ~a10852;
assign a10858 = ~a10856 & a10772;
assign a10860 = ~a10858 & ~a10836;
assign a10862 = ~a10860 & ~a10768;
assign a10864 = a10786 & ~l786;
assign a10866 = a10864 & ~a10784;
assign a10868 = a10784 & ~l772;
assign a10870 = ~a10868 & ~a10866;
assign a10872 = ~a10870 & ~a10782;
assign a10874 = a10782 & ~l758;
assign a10876 = ~a10874 & ~a10872;
assign a10878 = ~a10876 & ~a10780;
assign a10880 = a10780 & ~l744;
assign a10882 = ~a10880 & ~a10878;
assign a10884 = ~a10882 & a10768;
assign a10886 = ~a10884 & ~a10862;
assign a10888 = a10886 & ~l1014;
assign a10890 = ~a10886 & l1014;
assign a10892 = ~a10890 & ~a10888;
assign a10894 = a10786 & l1034;
assign a10896 = a10894 & ~a10784;
assign a10898 = a10784 & l1020;
assign a10900 = ~a10898 & ~a10896;
assign a10902 = ~a10900 & ~a10782;
assign a10904 = a10782 & l1006;
assign a10906 = ~a10904 & ~a10902;
assign a10908 = ~a10906 & ~a10780;
assign a10910 = a10780 & l992;
assign a10912 = ~a10910 & ~a10908;
assign a10914 = ~a10912 & a10778;
assign a10916 = a10914 & ~a10776;
assign a10918 = a10786 & l952;
assign a10920 = a10918 & ~a10784;
assign a10922 = a10784 & l938;
assign a10924 = ~a10922 & ~a10920;
assign a10926 = ~a10924 & ~a10782;
assign a10928 = a10782 & l924;
assign a10930 = ~a10928 & ~a10926;
assign a10932 = ~a10930 & ~a10780;
assign a10934 = a10780 & l910;
assign a10936 = ~a10934 & ~a10932;
assign a10938 = ~a10936 & a10776;
assign a10940 = ~a10938 & ~a10916;
assign a10942 = ~a10940 & ~a10772;
assign a10944 = a10786 & l870;
assign a10946 = a10944 & ~a10784;
assign a10948 = a10784 & l856;
assign a10950 = ~a10948 & ~a10946;
assign a10952 = ~a10950 & ~a10782;
assign a10954 = a10782 & l842;
assign a10956 = ~a10954 & ~a10952;
assign a10958 = ~a10956 & ~a10780;
assign a10960 = a10780 & l828;
assign a10962 = ~a10960 & ~a10958;
assign a10964 = ~a10962 & a10772;
assign a10966 = ~a10964 & ~a10942;
assign a10968 = ~a10966 & ~a10768;
assign a10970 = a10786 & l788;
assign a10972 = a10970 & ~a10784;
assign a10974 = a10784 & l774;
assign a10976 = ~a10974 & ~a10972;
assign a10978 = ~a10976 & ~a10782;
assign a10980 = a10782 & l760;
assign a10982 = ~a10980 & ~a10978;
assign a10984 = ~a10982 & ~a10780;
assign a10986 = a10780 & l746;
assign a10988 = ~a10986 & ~a10984;
assign a10990 = ~a10988 & a10768;
assign a10992 = ~a10990 & ~a10968;
assign a10994 = a10992 & ~l1016;
assign a10996 = ~a10992 & l1016;
assign a10998 = ~a10996 & ~a10994;
assign a11000 = a10998 & a10892;
assign a11002 = ~a11000 & ~a10764;
assign a11004 = a7188 & ~l730;
assign a11006 = l734 & ~l732;
assign a11008 = a11006 & ~l730;
assign a11010 = ~l734 & l732;
assign a11012 = a11010 & ~l730;
assign a11014 = l734 & l732;
assign a11016 = a11014 & ~l730;
assign a11018 = a7188 & l730;
assign a11020 = ~l738 & ~l736;
assign a11022 = l738 & ~l736;
assign a11024 = ~l738 & l736;
assign a11026 = l738 & l736;
assign a11028 = a11026 & ~l1032;
assign a11030 = a11028 & ~a11024;
assign a11032 = a11024 & ~l1018;
assign a11034 = ~a11032 & ~a11030;
assign a11036 = ~a11034 & ~a11022;
assign a11038 = a11022 & ~l1004;
assign a11040 = ~a11038 & ~a11036;
assign a11042 = ~a11040 & ~a11020;
assign a11044 = a11020 & ~l990;
assign a11046 = ~a11044 & ~a11042;
assign a11048 = ~a11046 & a11018;
assign a11050 = a11048 & ~a11016;
assign a11052 = a11026 & ~l950;
assign a11054 = a11052 & ~a11024;
assign a11056 = a11024 & ~l936;
assign a11058 = ~a11056 & ~a11054;
assign a11060 = ~a11058 & ~a11022;
assign a11062 = a11022 & ~l922;
assign a11064 = ~a11062 & ~a11060;
assign a11066 = ~a11064 & ~a11020;
assign a11068 = a11020 & ~l908;
assign a11070 = ~a11068 & ~a11066;
assign a11072 = ~a11070 & a11016;
assign a11074 = ~a11072 & ~a11050;
assign a11076 = ~a11074 & ~a11012;
assign a11078 = a11026 & ~l868;
assign a11080 = a11078 & ~a11024;
assign a11082 = a11024 & ~l854;
assign a11084 = ~a11082 & ~a11080;
assign a11086 = ~a11084 & ~a11022;
assign a11088 = a11022 & ~l840;
assign a11090 = ~a11088 & ~a11086;
assign a11092 = ~a11090 & ~a11020;
assign a11094 = a11020 & ~l826;
assign a11096 = ~a11094 & ~a11092;
assign a11098 = ~a11096 & a11012;
assign a11100 = ~a11098 & ~a11076;
assign a11102 = ~a11100 & ~a11008;
assign a11104 = a11026 & ~l786;
assign a11106 = a11104 & ~a11024;
assign a11108 = a11024 & ~l772;
assign a11110 = ~a11108 & ~a11106;
assign a11112 = ~a11110 & ~a11022;
assign a11114 = a11022 & ~l758;
assign a11116 = ~a11114 & ~a11112;
assign a11118 = ~a11116 & ~a11020;
assign a11120 = a11020 & ~l744;
assign a11122 = ~a11120 & ~a11118;
assign a11124 = ~a11122 & a11008;
assign a11126 = ~a11124 & ~a11102;
assign a11128 = a11126 & ~l1028;
assign a11130 = ~a11126 & l1028;
assign a11132 = ~a11130 & ~a11128;
assign a11134 = a11026 & l1034;
assign a11136 = a11134 & ~a11024;
assign a11138 = a11024 & l1020;
assign a11140 = ~a11138 & ~a11136;
assign a11142 = ~a11140 & ~a11022;
assign a11144 = a11022 & l1006;
assign a11146 = ~a11144 & ~a11142;
assign a11148 = ~a11146 & ~a11020;
assign a11150 = a11020 & l992;
assign a11152 = ~a11150 & ~a11148;
assign a11154 = ~a11152 & a11018;
assign a11156 = a11154 & ~a11016;
assign a11158 = a11026 & l952;
assign a11160 = a11158 & ~a11024;
assign a11162 = a11024 & l938;
assign a11164 = ~a11162 & ~a11160;
assign a11166 = ~a11164 & ~a11022;
assign a11168 = a11022 & l924;
assign a11170 = ~a11168 & ~a11166;
assign a11172 = ~a11170 & ~a11020;
assign a11174 = a11020 & l910;
assign a11176 = ~a11174 & ~a11172;
assign a11178 = ~a11176 & a11016;
assign a11180 = ~a11178 & ~a11156;
assign a11182 = ~a11180 & ~a11012;
assign a11184 = a11026 & l870;
assign a11186 = a11184 & ~a11024;
assign a11188 = a11024 & l856;
assign a11190 = ~a11188 & ~a11186;
assign a11192 = ~a11190 & ~a11022;
assign a11194 = a11022 & l842;
assign a11196 = ~a11194 & ~a11192;
assign a11198 = ~a11196 & ~a11020;
assign a11200 = a11020 & l828;
assign a11202 = ~a11200 & ~a11198;
assign a11204 = ~a11202 & a11012;
assign a11206 = ~a11204 & ~a11182;
assign a11208 = ~a11206 & ~a11008;
assign a11210 = a11026 & l788;
assign a11212 = a11210 & ~a11024;
assign a11214 = a11024 & l774;
assign a11216 = ~a11214 & ~a11212;
assign a11218 = ~a11216 & ~a11022;
assign a11220 = a11022 & l760;
assign a11222 = ~a11220 & ~a11218;
assign a11224 = ~a11222 & ~a11020;
assign a11226 = a11020 & l746;
assign a11228 = ~a11226 & ~a11224;
assign a11230 = ~a11228 & a11008;
assign a11232 = ~a11230 & ~a11208;
assign a11234 = a11232 & ~l1030;
assign a11236 = ~a11232 & l1030;
assign a11238 = ~a11236 & ~a11234;
assign a11240 = a11238 & a11132;
assign a11242 = ~a11240 & ~a11004;
assign a11244 = a11020 & a11008;
assign a11246 = ~a11244 & a7426;
assign a11248 = a11246 & ~a7424;
assign a11250 = a10780 & a10768;
assign a11252 = ~a11250 & a7424;
assign a11254 = ~a11252 & ~a11248;
assign a11256 = ~a11254 & ~a7422;
assign a11258 = a10540 & a10528;
assign a11260 = ~a11258 & a7422;
assign a11262 = ~a11260 & ~a11256;
assign a11264 = ~a11262 & ~a7420;
assign a11266 = a10300 & a10288;
assign a11268 = ~a11266 & a7420;
assign a11270 = ~a11268 & ~a11264;
assign a11272 = ~a11270 & a7418;
assign a11274 = a11272 & ~a7416;
assign a11276 = a10060 & a10048;
assign a11278 = ~a11276 & a7426;
assign a11280 = a11278 & ~a7424;
assign a11282 = a9820 & a9808;
assign a11284 = ~a11282 & a7424;
assign a11286 = ~a11284 & ~a11280;
assign a11288 = ~a11286 & ~a7422;
assign a11290 = a9580 & a9568;
assign a11292 = ~a11290 & a7422;
assign a11294 = ~a11292 & ~a11288;
assign a11296 = ~a11294 & ~a7420;
assign a11298 = a9340 & a9328;
assign a11300 = ~a11298 & a7420;
assign a11302 = ~a11300 & ~a11296;
assign a11304 = ~a11302 & a7416;
assign a11306 = ~a11304 & ~a11274;
assign a11308 = ~a11306 & ~a7412;
assign a11310 = a9100 & a9088;
assign a11312 = ~a11310 & a7426;
assign a11314 = a11312 & ~a7424;
assign a11316 = a8860 & a8848;
assign a11318 = ~a11316 & a7424;
assign a11320 = ~a11318 & ~a11314;
assign a11322 = ~a11320 & ~a7422;
assign a11324 = a8620 & a8608;
assign a11326 = ~a11324 & a7422;
assign a11328 = ~a11326 & ~a11322;
assign a11330 = ~a11328 & ~a7420;
assign a11332 = a8380 & a8368;
assign a11334 = ~a11332 & a7420;
assign a11336 = ~a11334 & ~a11330;
assign a11338 = ~a11336 & a7412;
assign a11340 = ~a11338 & ~a11308;
assign a11342 = ~a11340 & ~a7408;
assign a11344 = a8140 & a8128;
assign a11346 = ~a11344 & a7426;
assign a11348 = a11346 & ~a7424;
assign a11350 = a7900 & a7888;
assign a11352 = ~a11350 & a7424;
assign a11354 = ~a11352 & ~a11348;
assign a11356 = ~a11354 & ~a7422;
assign a11358 = a7660 & a7648;
assign a11360 = ~a11358 & a7422;
assign a11362 = ~a11360 & ~a11356;
assign a11364 = ~a11362 & ~a7420;
assign a11366 = a7420 & ~a7408;
assign a11368 = ~a11366 & ~a11364;
assign a11370 = ~a11368 & a7408;
assign a11372 = ~a11370 & ~a11342;
assign a11374 = a11022 & a11008;
assign a11376 = ~a11374 & a7666;
assign a11378 = a11376 & ~a7664;
assign a11380 = a10782 & a10768;
assign a11382 = ~a11380 & a7664;
assign a11384 = ~a11382 & ~a11378;
assign a11386 = ~a11384 & ~a7662;
assign a11388 = a10542 & a10528;
assign a11390 = ~a11388 & a7662;
assign a11392 = ~a11390 & ~a11386;
assign a11394 = ~a11392 & ~a7660;
assign a11396 = a10302 & a10288;
assign a11398 = ~a11396 & a7660;
assign a11400 = ~a11398 & ~a11394;
assign a11402 = ~a11400 & a7658;
assign a11404 = a11402 & ~a7656;
assign a11406 = a10062 & a10048;
assign a11408 = ~a11406 & a7666;
assign a11410 = a11408 & ~a7664;
assign a11412 = a9822 & a9808;
assign a11414 = ~a11412 & a7664;
assign a11416 = ~a11414 & ~a11410;
assign a11418 = ~a11416 & ~a7662;
assign a11420 = a9582 & a9568;
assign a11422 = ~a11420 & a7662;
assign a11424 = ~a11422 & ~a11418;
assign a11426 = ~a11424 & ~a7660;
assign a11428 = a9342 & a9328;
assign a11430 = ~a11428 & a7660;
assign a11432 = ~a11430 & ~a11426;
assign a11434 = ~a11432 & a7656;
assign a11436 = ~a11434 & ~a11404;
assign a11438 = ~a11436 & ~a7652;
assign a11440 = a9102 & a9088;
assign a11442 = ~a11440 & a7666;
assign a11444 = a11442 & ~a7664;
assign a11446 = a8862 & a8848;
assign a11448 = ~a11446 & a7664;
assign a11450 = ~a11448 & ~a11444;
assign a11452 = ~a11450 & ~a7662;
assign a11454 = a8622 & a8608;
assign a11456 = ~a11454 & a7662;
assign a11458 = ~a11456 & ~a11452;
assign a11460 = ~a11458 & ~a7660;
assign a11462 = a8382 & a8368;
assign a11464 = ~a11462 & a7660;
assign a11466 = ~a11464 & ~a11460;
assign a11468 = ~a11466 & a7652;
assign a11470 = ~a11468 & ~a11438;
assign a11472 = ~a11470 & ~a7648;
assign a11474 = a8142 & a8128;
assign a11476 = ~a11474 & a7666;
assign a11478 = a11476 & ~a7664;
assign a11480 = a7902 & a7888;
assign a11482 = ~a11480 & a7664;
assign a11484 = ~a11482 & ~a11478;
assign a11486 = ~a11484 & ~a7662;
assign a11488 = a7662 & ~a7648;
assign a11490 = ~a11488 & ~a11486;
assign a11492 = ~a11490 & ~a7660;
assign a11494 = a7422 & a7408;
assign a11496 = ~a11494 & a7660;
assign a11498 = ~a11496 & ~a11492;
assign a11500 = ~a11498 & a7648;
assign a11502 = ~a11500 & ~a11472;
assign a11504 = a11024 & a11008;
assign a11506 = ~a11504 & a7906;
assign a11508 = a11506 & ~a7904;
assign a11510 = a10784 & a10768;
assign a11512 = ~a11510 & a7904;
assign a11514 = ~a11512 & ~a11508;
assign a11516 = ~a11514 & ~a7902;
assign a11518 = a10544 & a10528;
assign a11520 = ~a11518 & a7902;
assign a11522 = ~a11520 & ~a11516;
assign a11524 = ~a11522 & ~a7900;
assign a11526 = a10304 & a10288;
assign a11528 = ~a11526 & a7900;
assign a11530 = ~a11528 & ~a11524;
assign a11532 = ~a11530 & a7898;
assign a11534 = a11532 & ~a7896;
assign a11536 = a10064 & a10048;
assign a11538 = ~a11536 & a7906;
assign a11540 = a11538 & ~a7904;
assign a11542 = a9824 & a9808;
assign a11544 = ~a11542 & a7904;
assign a11546 = ~a11544 & ~a11540;
assign a11548 = ~a11546 & ~a7902;
assign a11550 = a9584 & a9568;
assign a11552 = ~a11550 & a7902;
assign a11554 = ~a11552 & ~a11548;
assign a11556 = ~a11554 & ~a7900;
assign a11558 = a9344 & a9328;
assign a11560 = ~a11558 & a7900;
assign a11562 = ~a11560 & ~a11556;
assign a11564 = ~a11562 & a7896;
assign a11566 = ~a11564 & ~a11534;
assign a11568 = ~a11566 & ~a7892;
assign a11570 = a9104 & a9088;
assign a11572 = ~a11570 & a7906;
assign a11574 = a11572 & ~a7904;
assign a11576 = a8864 & a8848;
assign a11578 = ~a11576 & a7904;
assign a11580 = ~a11578 & ~a11574;
assign a11582 = ~a11580 & ~a7902;
assign a11584 = a8624 & a8608;
assign a11586 = ~a11584 & a7902;
assign a11588 = ~a11586 & ~a11582;
assign a11590 = ~a11588 & ~a7900;
assign a11592 = a8384 & a8368;
assign a11594 = ~a11592 & a7900;
assign a11596 = ~a11594 & ~a11590;
assign a11598 = ~a11596 & a7892;
assign a11600 = ~a11598 & ~a11568;
assign a11602 = ~a11600 & ~a7888;
assign a11604 = a8144 & a8128;
assign a11606 = ~a11604 & a7906;
assign a11608 = a11606 & ~a7904;
assign a11610 = a7904 & ~a7888;
assign a11612 = ~a11610 & ~a11608;
assign a11614 = ~a11612 & ~a7902;
assign a11616 = a7664 & a7648;
assign a11618 = ~a11616 & a7902;
assign a11620 = ~a11618 & ~a11614;
assign a11622 = ~a11620 & ~a7900;
assign a11624 = a7424 & a7408;
assign a11626 = ~a11624 & a7900;
assign a11628 = ~a11626 & ~a11622;
assign a11630 = ~a11628 & a7888;
assign a11632 = ~a11630 & ~a11602;
assign a11634 = a11026 & a11008;
assign a11636 = ~a11634 & a8146;
assign a11638 = a11636 & ~a8144;
assign a11640 = a10786 & a10768;
assign a11642 = ~a11640 & a8144;
assign a11644 = ~a11642 & ~a11638;
assign a11646 = ~a11644 & ~a8142;
assign a11648 = a10546 & a10528;
assign a11650 = ~a11648 & a8142;
assign a11652 = ~a11650 & ~a11646;
assign a11654 = ~a11652 & ~a8140;
assign a11656 = a10306 & a10288;
assign a11658 = ~a11656 & a8140;
assign a11660 = ~a11658 & ~a11654;
assign a11662 = ~a11660 & a8138;
assign a11664 = a11662 & ~a8136;
assign a11666 = a10066 & a10048;
assign a11668 = ~a11666 & a8146;
assign a11670 = a11668 & ~a8144;
assign a11672 = a9826 & a9808;
assign a11674 = ~a11672 & a8144;
assign a11676 = ~a11674 & ~a11670;
assign a11678 = ~a11676 & ~a8142;
assign a11680 = a9586 & a9568;
assign a11682 = ~a11680 & a8142;
assign a11684 = ~a11682 & ~a11678;
assign a11686 = ~a11684 & ~a8140;
assign a11688 = a9346 & a9328;
assign a11690 = ~a11688 & a8140;
assign a11692 = ~a11690 & ~a11686;
assign a11694 = ~a11692 & a8136;
assign a11696 = ~a11694 & ~a11664;
assign a11698 = ~a11696 & ~a8132;
assign a11700 = a9106 & a9088;
assign a11702 = ~a11700 & a8146;
assign a11704 = a11702 & ~a8144;
assign a11706 = a8866 & a8848;
assign a11708 = ~a11706 & a8144;
assign a11710 = ~a11708 & ~a11704;
assign a11712 = ~a11710 & ~a8142;
assign a11714 = a8626 & a8608;
assign a11716 = ~a11714 & a8142;
assign a11718 = ~a11716 & ~a11712;
assign a11720 = ~a11718 & ~a8140;
assign a11722 = a8386 & a8368;
assign a11724 = ~a11722 & a8140;
assign a11726 = ~a11724 & ~a11720;
assign a11728 = ~a11726 & a8132;
assign a11730 = ~a11728 & ~a11698;
assign a11732 = ~a11730 & ~a8128;
assign a11734 = a8146 & ~a8128;
assign a11736 = a11734 & ~a8144;
assign a11738 = a7906 & a7888;
assign a11740 = ~a11738 & a8144;
assign a11742 = ~a11740 & ~a11736;
assign a11744 = ~a11742 & ~a8142;
assign a11746 = a7666 & a7648;
assign a11748 = ~a11746 & a8142;
assign a11750 = ~a11748 & ~a11744;
assign a11752 = ~a11750 & ~a8140;
assign a11754 = a7426 & a7408;
assign a11756 = ~a11754 & a8140;
assign a11758 = ~a11756 & ~a11752;
assign a11760 = ~a11758 & a8128;
assign a11762 = ~a11760 & ~a11732;
assign a11764 = a11020 & a11012;
assign a11766 = ~a11764 & a8386;
assign a11768 = a11766 & ~a8384;
assign a11770 = a10780 & a10772;
assign a11772 = ~a11770 & a8384;
assign a11774 = ~a11772 & ~a11768;
assign a11776 = ~a11774 & ~a8382;
assign a11778 = a10540 & a10532;
assign a11780 = ~a11778 & a8382;
assign a11782 = ~a11780 & ~a11776;
assign a11784 = ~a11782 & ~a8380;
assign a11786 = a10300 & a10292;
assign a11788 = ~a11786 & a8380;
assign a11790 = ~a11788 & ~a11784;
assign a11792 = ~a11790 & a8378;
assign a11794 = a11792 & ~a8376;
assign a11796 = a10060 & a10052;
assign a11798 = ~a11796 & a8386;
assign a11800 = a11798 & ~a8384;
assign a11802 = a9820 & a9812;
assign a11804 = ~a11802 & a8384;
assign a11806 = ~a11804 & ~a11800;
assign a11808 = ~a11806 & ~a8382;
assign a11810 = a9580 & a9572;
assign a11812 = ~a11810 & a8382;
assign a11814 = ~a11812 & ~a11808;
assign a11816 = ~a11814 & ~a8380;
assign a11818 = a9340 & a9332;
assign a11820 = ~a11818 & a8380;
assign a11822 = ~a11820 & ~a11816;
assign a11824 = ~a11822 & a8376;
assign a11826 = ~a11824 & ~a11794;
assign a11828 = ~a11826 & ~a8372;
assign a11830 = a9100 & a9092;
assign a11832 = ~a11830 & a8386;
assign a11834 = a11832 & ~a8384;
assign a11836 = a8860 & a8852;
assign a11838 = ~a11836 & a8384;
assign a11840 = ~a11838 & ~a11834;
assign a11842 = ~a11840 & ~a8382;
assign a11844 = a8620 & a8612;
assign a11846 = ~a11844 & a8382;
assign a11848 = ~a11846 & ~a11842;
assign a11850 = ~a11848 & ~a8380;
assign a11852 = a8380 & ~a8372;
assign a11854 = ~a11852 & ~a11850;
assign a11856 = ~a11854 & a8372;
assign a11858 = ~a11856 & ~a11828;
assign a11860 = ~a11858 & ~a8368;
assign a11862 = a8140 & a8132;
assign a11864 = ~a11862 & a8386;
assign a11866 = a11864 & ~a8384;
assign a11868 = a7900 & a7892;
assign a11870 = ~a11868 & a8384;
assign a11872 = ~a11870 & ~a11866;
assign a11874 = ~a11872 & ~a8382;
assign a11876 = a7660 & a7652;
assign a11878 = ~a11876 & a8382;
assign a11880 = ~a11878 & ~a11874;
assign a11882 = ~a11880 & ~a8380;
assign a11884 = a7420 & a7412;
assign a11886 = ~a11884 & a8380;
assign a11888 = ~a11886 & ~a11882;
assign a11890 = ~a11888 & a8368;
assign a11892 = ~a11890 & ~a11860;
assign a11894 = a11022 & a11012;
assign a11896 = ~a11894 & a8626;
assign a11898 = a11896 & ~a8624;
assign a11900 = a10782 & a10772;
assign a11902 = ~a11900 & a8624;
assign a11904 = ~a11902 & ~a11898;
assign a11906 = ~a11904 & ~a8622;
assign a11908 = a10542 & a10532;
assign a11910 = ~a11908 & a8622;
assign a11912 = ~a11910 & ~a11906;
assign a11914 = ~a11912 & ~a8620;
assign a11916 = a10302 & a10292;
assign a11918 = ~a11916 & a8620;
assign a11920 = ~a11918 & ~a11914;
assign a11922 = ~a11920 & a8618;
assign a11924 = a11922 & ~a8616;
assign a11926 = a10062 & a10052;
assign a11928 = ~a11926 & a8626;
assign a11930 = a11928 & ~a8624;
assign a11932 = a9822 & a9812;
assign a11934 = ~a11932 & a8624;
assign a11936 = ~a11934 & ~a11930;
assign a11938 = ~a11936 & ~a8622;
assign a11940 = a9582 & a9572;
assign a11942 = ~a11940 & a8622;
assign a11944 = ~a11942 & ~a11938;
assign a11946 = ~a11944 & ~a8620;
assign a11948 = a9342 & a9332;
assign a11950 = ~a11948 & a8620;
assign a11952 = ~a11950 & ~a11946;
assign a11954 = ~a11952 & a8616;
assign a11956 = ~a11954 & ~a11924;
assign a11958 = ~a11956 & ~a8612;
assign a11960 = a9102 & a9092;
assign a11962 = ~a11960 & a8626;
assign a11964 = a11962 & ~a8624;
assign a11966 = a8862 & a8852;
assign a11968 = ~a11966 & a8624;
assign a11970 = ~a11968 & ~a11964;
assign a11972 = ~a11970 & ~a8622;
assign a11974 = a8622 & ~a8612;
assign a11976 = ~a11974 & ~a11972;
assign a11978 = ~a11976 & ~a8620;
assign a11980 = a8382 & a8372;
assign a11982 = ~a11980 & a8620;
assign a11984 = ~a11982 & ~a11978;
assign a11986 = ~a11984 & a8612;
assign a11988 = ~a11986 & ~a11958;
assign a11990 = ~a11988 & ~a8608;
assign a11992 = a8142 & a8132;
assign a11994 = ~a11992 & a8626;
assign a11996 = a11994 & ~a8624;
assign a11998 = a7902 & a7892;
assign a12000 = ~a11998 & a8624;
assign a12002 = ~a12000 & ~a11996;
assign a12004 = ~a12002 & ~a8622;
assign a12006 = a7662 & a7652;
assign a12008 = ~a12006 & a8622;
assign a12010 = ~a12008 & ~a12004;
assign a12012 = ~a12010 & ~a8620;
assign a12014 = a7422 & a7412;
assign a12016 = ~a12014 & a8620;
assign a12018 = ~a12016 & ~a12012;
assign a12020 = ~a12018 & a8608;
assign a12022 = ~a12020 & ~a11990;
assign a12024 = a11024 & a11012;
assign a12026 = ~a12024 & a8866;
assign a12028 = a12026 & ~a8864;
assign a12030 = a10784 & a10772;
assign a12032 = ~a12030 & a8864;
assign a12034 = ~a12032 & ~a12028;
assign a12036 = ~a12034 & ~a8862;
assign a12038 = a10544 & a10532;
assign a12040 = ~a12038 & a8862;
assign a12042 = ~a12040 & ~a12036;
assign a12044 = ~a12042 & ~a8860;
assign a12046 = a10304 & a10292;
assign a12048 = ~a12046 & a8860;
assign a12050 = ~a12048 & ~a12044;
assign a12052 = ~a12050 & a8858;
assign a12054 = a12052 & ~a8856;
assign a12056 = a10064 & a10052;
assign a12058 = ~a12056 & a8866;
assign a12060 = a12058 & ~a8864;
assign a12062 = a9824 & a9812;
assign a12064 = ~a12062 & a8864;
assign a12066 = ~a12064 & ~a12060;
assign a12068 = ~a12066 & ~a8862;
assign a12070 = a9584 & a9572;
assign a12072 = ~a12070 & a8862;
assign a12074 = ~a12072 & ~a12068;
assign a12076 = ~a12074 & ~a8860;
assign a12078 = a9344 & a9332;
assign a12080 = ~a12078 & a8860;
assign a12082 = ~a12080 & ~a12076;
assign a12084 = ~a12082 & a8856;
assign a12086 = ~a12084 & ~a12054;
assign a12088 = ~a12086 & ~a8852;
assign a12090 = a9104 & a9092;
assign a12092 = ~a12090 & a8866;
assign a12094 = a12092 & ~a8864;
assign a12096 = a8864 & ~a8852;
assign a12098 = ~a12096 & ~a12094;
assign a12100 = ~a12098 & ~a8862;
assign a12102 = a8624 & a8612;
assign a12104 = ~a12102 & a8862;
assign a12106 = ~a12104 & ~a12100;
assign a12108 = ~a12106 & ~a8860;
assign a12110 = a8384 & a8372;
assign a12112 = ~a12110 & a8860;
assign a12114 = ~a12112 & ~a12108;
assign a12116 = ~a12114 & a8852;
assign a12118 = ~a12116 & ~a12088;
assign a12120 = ~a12118 & ~a8848;
assign a12122 = a8144 & a8132;
assign a12124 = ~a12122 & a8866;
assign a12126 = a12124 & ~a8864;
assign a12128 = a7904 & a7892;
assign a12130 = ~a12128 & a8864;
assign a12132 = ~a12130 & ~a12126;
assign a12134 = ~a12132 & ~a8862;
assign a12136 = a7664 & a7652;
assign a12138 = ~a12136 & a8862;
assign a12140 = ~a12138 & ~a12134;
assign a12142 = ~a12140 & ~a8860;
assign a12144 = a7424 & a7412;
assign a12146 = ~a12144 & a8860;
assign a12148 = ~a12146 & ~a12142;
assign a12150 = ~a12148 & a8848;
assign a12152 = ~a12150 & ~a12120;
assign a12154 = a11026 & a11012;
assign a12156 = ~a12154 & a9106;
assign a12158 = a12156 & ~a9104;
assign a12160 = a10786 & a10772;
assign a12162 = ~a12160 & a9104;
assign a12164 = ~a12162 & ~a12158;
assign a12166 = ~a12164 & ~a9102;
assign a12168 = a10546 & a10532;
assign a12170 = ~a12168 & a9102;
assign a12172 = ~a12170 & ~a12166;
assign a12174 = ~a12172 & ~a9100;
assign a12176 = a10306 & a10292;
assign a12178 = ~a12176 & a9100;
assign a12180 = ~a12178 & ~a12174;
assign a12182 = ~a12180 & a9098;
assign a12184 = a12182 & ~a9096;
assign a12186 = a10066 & a10052;
assign a12188 = ~a12186 & a9106;
assign a12190 = a12188 & ~a9104;
assign a12192 = a9826 & a9812;
assign a12194 = ~a12192 & a9104;
assign a12196 = ~a12194 & ~a12190;
assign a12198 = ~a12196 & ~a9102;
assign a12200 = a9586 & a9572;
assign a12202 = ~a12200 & a9102;
assign a12204 = ~a12202 & ~a12198;
assign a12206 = ~a12204 & ~a9100;
assign a12208 = a9346 & a9332;
assign a12210 = ~a12208 & a9100;
assign a12212 = ~a12210 & ~a12206;
assign a12214 = ~a12212 & a9096;
assign a12216 = ~a12214 & ~a12184;
assign a12218 = ~a12216 & ~a9092;
assign a12220 = a9106 & ~a9092;
assign a12222 = a12220 & ~a9104;
assign a12224 = a8866 & a8852;
assign a12226 = ~a12224 & a9104;
assign a12228 = ~a12226 & ~a12222;
assign a12230 = ~a12228 & ~a9102;
assign a12232 = a8626 & a8612;
assign a12234 = ~a12232 & a9102;
assign a12236 = ~a12234 & ~a12230;
assign a12238 = ~a12236 & ~a9100;
assign a12240 = a8386 & a8372;
assign a12242 = ~a12240 & a9100;
assign a12244 = ~a12242 & ~a12238;
assign a12246 = ~a12244 & a9092;
assign a12248 = ~a12246 & ~a12218;
assign a12250 = ~a12248 & ~a9088;
assign a12252 = a8146 & a8132;
assign a12254 = ~a12252 & a9106;
assign a12256 = a12254 & ~a9104;
assign a12258 = a7906 & a7892;
assign a12260 = ~a12258 & a9104;
assign a12262 = ~a12260 & ~a12256;
assign a12264 = ~a12262 & ~a9102;
assign a12266 = a7666 & a7652;
assign a12268 = ~a12266 & a9102;
assign a12270 = ~a12268 & ~a12264;
assign a12272 = ~a12270 & ~a9100;
assign a12274 = a7426 & a7412;
assign a12276 = ~a12274 & a9100;
assign a12278 = ~a12276 & ~a12272;
assign a12280 = ~a12278 & a9088;
assign a12282 = ~a12280 & ~a12250;
assign a12284 = a11020 & a11016;
assign a12286 = ~a12284 & a9346;
assign a12288 = a12286 & ~a9344;
assign a12290 = a10780 & a10776;
assign a12292 = ~a12290 & a9344;
assign a12294 = ~a12292 & ~a12288;
assign a12296 = ~a12294 & ~a9342;
assign a12298 = a10540 & a10536;
assign a12300 = ~a12298 & a9342;
assign a12302 = ~a12300 & ~a12296;
assign a12304 = ~a12302 & ~a9340;
assign a12306 = a10300 & a10296;
assign a12308 = ~a12306 & a9340;
assign a12310 = ~a12308 & ~a12304;
assign a12312 = ~a12310 & a9338;
assign a12314 = a12312 & ~a9336;
assign a12316 = a10060 & a10056;
assign a12318 = ~a12316 & a9346;
assign a12320 = a12318 & ~a9344;
assign a12322 = a9820 & a9816;
assign a12324 = ~a12322 & a9344;
assign a12326 = ~a12324 & ~a12320;
assign a12328 = ~a12326 & ~a9342;
assign a12330 = a9580 & a9576;
assign a12332 = ~a12330 & a9342;
assign a12334 = ~a12332 & ~a12328;
assign a12336 = ~a12334 & ~a9340;
assign a12338 = a9340 & ~a9336;
assign a12340 = ~a12338 & ~a12336;
assign a12342 = ~a12340 & a9336;
assign a12344 = ~a12342 & ~a12314;
assign a12346 = ~a12344 & ~a9332;
assign a12348 = a9100 & a9096;
assign a12350 = ~a12348 & a9346;
assign a12352 = a12350 & ~a9344;
assign a12354 = a8860 & a8856;
assign a12356 = ~a12354 & a9344;
assign a12358 = ~a12356 & ~a12352;
assign a12360 = ~a12358 & ~a9342;
assign a12362 = a8620 & a8616;
assign a12364 = ~a12362 & a9342;
assign a12366 = ~a12364 & ~a12360;
assign a12368 = ~a12366 & ~a9340;
assign a12370 = a8380 & a8376;
assign a12372 = ~a12370 & a9340;
assign a12374 = ~a12372 & ~a12368;
assign a12376 = ~a12374 & a9332;
assign a12378 = ~a12376 & ~a12346;
assign a12380 = ~a12378 & ~a9328;
assign a12382 = a8140 & a8136;
assign a12384 = ~a12382 & a9346;
assign a12386 = a12384 & ~a9344;
assign a12388 = a7900 & a7896;
assign a12390 = ~a12388 & a9344;
assign a12392 = ~a12390 & ~a12386;
assign a12394 = ~a12392 & ~a9342;
assign a12396 = a7660 & a7656;
assign a12398 = ~a12396 & a9342;
assign a12400 = ~a12398 & ~a12394;
assign a12402 = ~a12400 & ~a9340;
assign a12404 = a7420 & a7416;
assign a12406 = ~a12404 & a9340;
assign a12408 = ~a12406 & ~a12402;
assign a12410 = ~a12408 & a9328;
assign a12412 = ~a12410 & ~a12380;
assign a12414 = a11022 & a11016;
assign a12416 = ~a12414 & a9586;
assign a12418 = a12416 & ~a9584;
assign a12420 = a10782 & a10776;
assign a12422 = ~a12420 & a9584;
assign a12424 = ~a12422 & ~a12418;
assign a12426 = ~a12424 & ~a9582;
assign a12428 = a10542 & a10536;
assign a12430 = ~a12428 & a9582;
assign a12432 = ~a12430 & ~a12426;
assign a12434 = ~a12432 & ~a9580;
assign a12436 = a10302 & a10296;
assign a12438 = ~a12436 & a9580;
assign a12440 = ~a12438 & ~a12434;
assign a12442 = ~a12440 & a9578;
assign a12444 = a12442 & ~a9576;
assign a12446 = a10062 & a10056;
assign a12448 = ~a12446 & a9586;
assign a12450 = a12448 & ~a9584;
assign a12452 = a9822 & a9816;
assign a12454 = ~a12452 & a9584;
assign a12456 = ~a12454 & ~a12450;
assign a12458 = ~a12456 & ~a9582;
assign a12460 = a9582 & ~a9576;
assign a12462 = ~a12460 & ~a12458;
assign a12464 = ~a12462 & ~a9580;
assign a12466 = a9342 & a9336;
assign a12468 = ~a12466 & a9580;
assign a12470 = ~a12468 & ~a12464;
assign a12472 = ~a12470 & a9576;
assign a12474 = ~a12472 & ~a12444;
assign a12476 = ~a12474 & ~a9572;
assign a12478 = a9102 & a9096;
assign a12480 = ~a12478 & a9586;
assign a12482 = a12480 & ~a9584;
assign a12484 = a8862 & a8856;
assign a12486 = ~a12484 & a9584;
assign a12488 = ~a12486 & ~a12482;
assign a12490 = ~a12488 & ~a9582;
assign a12492 = a8622 & a8616;
assign a12494 = ~a12492 & a9582;
assign a12496 = ~a12494 & ~a12490;
assign a12498 = ~a12496 & ~a9580;
assign a12500 = a8382 & a8376;
assign a12502 = ~a12500 & a9580;
assign a12504 = ~a12502 & ~a12498;
assign a12506 = ~a12504 & a9572;
assign a12508 = ~a12506 & ~a12476;
assign a12510 = ~a12508 & ~a9568;
assign a12512 = a8142 & a8136;
assign a12514 = ~a12512 & a9586;
assign a12516 = a12514 & ~a9584;
assign a12518 = a7902 & a7896;
assign a12520 = ~a12518 & a9584;
assign a12522 = ~a12520 & ~a12516;
assign a12524 = ~a12522 & ~a9582;
assign a12526 = a7662 & a7656;
assign a12528 = ~a12526 & a9582;
assign a12530 = ~a12528 & ~a12524;
assign a12532 = ~a12530 & ~a9580;
assign a12534 = a7422 & a7416;
assign a12536 = ~a12534 & a9580;
assign a12538 = ~a12536 & ~a12532;
assign a12540 = ~a12538 & a9568;
assign a12542 = ~a12540 & ~a12510;
assign a12544 = a11024 & a11016;
assign a12546 = ~a12544 & a9826;
assign a12548 = a12546 & ~a9824;
assign a12550 = a10784 & a10776;
assign a12552 = ~a12550 & a9824;
assign a12554 = ~a12552 & ~a12548;
assign a12556 = ~a12554 & ~a9822;
assign a12558 = a10544 & a10536;
assign a12560 = ~a12558 & a9822;
assign a12562 = ~a12560 & ~a12556;
assign a12564 = ~a12562 & ~a9820;
assign a12566 = a10304 & a10296;
assign a12568 = ~a12566 & a9820;
assign a12570 = ~a12568 & ~a12564;
assign a12572 = ~a12570 & a9818;
assign a12574 = a12572 & ~a9816;
assign a12576 = a10064 & a10056;
assign a12578 = ~a12576 & a9826;
assign a12580 = a12578 & ~a9824;
assign a12582 = a9824 & ~a9816;
assign a12584 = ~a12582 & ~a12580;
assign a12586 = ~a12584 & ~a9822;
assign a12588 = a9584 & a9576;
assign a12590 = ~a12588 & a9822;
assign a12592 = ~a12590 & ~a12586;
assign a12594 = ~a12592 & ~a9820;
assign a12596 = a9344 & a9336;
assign a12598 = ~a12596 & a9820;
assign a12600 = ~a12598 & ~a12594;
assign a12602 = ~a12600 & a9816;
assign a12604 = ~a12602 & ~a12574;
assign a12606 = ~a12604 & ~a9812;
assign a12608 = a9104 & a9096;
assign a12610 = ~a12608 & a9826;
assign a12612 = a12610 & ~a9824;
assign a12614 = a8864 & a8856;
assign a12616 = ~a12614 & a9824;
assign a12618 = ~a12616 & ~a12612;
assign a12620 = ~a12618 & ~a9822;
assign a12622 = a8624 & a8616;
assign a12624 = ~a12622 & a9822;
assign a12626 = ~a12624 & ~a12620;
assign a12628 = ~a12626 & ~a9820;
assign a12630 = a8384 & a8376;
assign a12632 = ~a12630 & a9820;
assign a12634 = ~a12632 & ~a12628;
assign a12636 = ~a12634 & a9812;
assign a12638 = ~a12636 & ~a12606;
assign a12640 = ~a12638 & ~a9808;
assign a12642 = a8144 & a8136;
assign a12644 = ~a12642 & a9826;
assign a12646 = a12644 & ~a9824;
assign a12648 = a7904 & a7896;
assign a12650 = ~a12648 & a9824;
assign a12652 = ~a12650 & ~a12646;
assign a12654 = ~a12652 & ~a9822;
assign a12656 = a7664 & a7656;
assign a12658 = ~a12656 & a9822;
assign a12660 = ~a12658 & ~a12654;
assign a12662 = ~a12660 & ~a9820;
assign a12664 = a7424 & a7416;
assign a12666 = ~a12664 & a9820;
assign a12668 = ~a12666 & ~a12662;
assign a12670 = ~a12668 & a9808;
assign a12672 = ~a12670 & ~a12640;
assign a12674 = a11026 & a11016;
assign a12676 = ~a12674 & a10066;
assign a12678 = a12676 & ~a10064;
assign a12680 = a10786 & a10776;
assign a12682 = ~a12680 & a10064;
assign a12684 = ~a12682 & ~a12678;
assign a12686 = ~a12684 & ~a10062;
assign a12688 = a10546 & a10536;
assign a12690 = ~a12688 & a10062;
assign a12692 = ~a12690 & ~a12686;
assign a12694 = ~a12692 & ~a10060;
assign a12696 = a10306 & a10296;
assign a12698 = ~a12696 & a10060;
assign a12700 = ~a12698 & ~a12694;
assign a12702 = ~a12700 & a10058;
assign a12704 = a12702 & ~a10056;
assign a12706 = a10066 & ~a10056;
assign a12708 = a12706 & ~a10064;
assign a12710 = a9826 & a9816;
assign a12712 = ~a12710 & a10064;
assign a12714 = ~a12712 & ~a12708;
assign a12716 = ~a12714 & ~a10062;
assign a12718 = a9586 & a9576;
assign a12720 = ~a12718 & a10062;
assign a12722 = ~a12720 & ~a12716;
assign a12724 = ~a12722 & ~a10060;
assign a12726 = a9346 & a9336;
assign a12728 = ~a12726 & a10060;
assign a12730 = ~a12728 & ~a12724;
assign a12732 = ~a12730 & a10056;
assign a12734 = ~a12732 & ~a12704;
assign a12736 = ~a12734 & ~a10052;
assign a12738 = a9106 & a9096;
assign a12740 = ~a12738 & a10066;
assign a12742 = a12740 & ~a10064;
assign a12744 = a8866 & a8856;
assign a12746 = ~a12744 & a10064;
assign a12748 = ~a12746 & ~a12742;
assign a12750 = ~a12748 & ~a10062;
assign a12752 = a8626 & a8616;
assign a12754 = ~a12752 & a10062;
assign a12756 = ~a12754 & ~a12750;
assign a12758 = ~a12756 & ~a10060;
assign a12760 = a8386 & a8376;
assign a12762 = ~a12760 & a10060;
assign a12764 = ~a12762 & ~a12758;
assign a12766 = ~a12764 & a10052;
assign a12768 = ~a12766 & ~a12736;
assign a12770 = ~a12768 & ~a10048;
assign a12772 = a8146 & a8136;
assign a12774 = ~a12772 & a10066;
assign a12776 = a12774 & ~a10064;
assign a12778 = a7906 & a7896;
assign a12780 = ~a12778 & a10064;
assign a12782 = ~a12780 & ~a12776;
assign a12784 = ~a12782 & ~a10062;
assign a12786 = a7666 & a7656;
assign a12788 = ~a12786 & a10062;
assign a12790 = ~a12788 & ~a12784;
assign a12792 = ~a12790 & ~a10060;
assign a12794 = a7426 & a7416;
assign a12796 = ~a12794 & a10060;
assign a12798 = ~a12796 & ~a12792;
assign a12800 = ~a12798 & a10048;
assign a12802 = ~a12800 & ~a12770;
assign a12804 = a11020 & a11018;
assign a12806 = ~a12804 & a10306;
assign a12808 = a12806 & ~a10304;
assign a12810 = a10780 & a10778;
assign a12812 = ~a12810 & a10304;
assign a12814 = ~a12812 & ~a12808;
assign a12816 = ~a12814 & ~a10302;
assign a12818 = a10540 & a10538;
assign a12820 = ~a12818 & a10302;
assign a12822 = ~a12820 & ~a12816;
assign a12824 = ~a12822 & ~a10300;
assign a12826 = a10300 & ~a10298;
assign a12828 = ~a12826 & ~a12824;
assign a12830 = ~a12828 & a10298;
assign a12832 = a12830 & ~a10296;
assign a12834 = a10060 & a10058;
assign a12836 = ~a12834 & a10306;
assign a12838 = a12836 & ~a10304;
assign a12840 = a9820 & a9818;
assign a12842 = ~a12840 & a10304;
assign a12844 = ~a12842 & ~a12838;
assign a12846 = ~a12844 & ~a10302;
assign a12848 = a9580 & a9578;
assign a12850 = ~a12848 & a10302;
assign a12852 = ~a12850 & ~a12846;
assign a12854 = ~a12852 & ~a10300;
assign a12856 = a9340 & a9338;
assign a12858 = ~a12856 & a10300;
assign a12860 = ~a12858 & ~a12854;
assign a12862 = ~a12860 & a10296;
assign a12864 = ~a12862 & ~a12832;
assign a12866 = ~a12864 & ~a10292;
assign a12868 = a9100 & a9098;
assign a12870 = ~a12868 & a10306;
assign a12872 = a12870 & ~a10304;
assign a12874 = a8860 & a8858;
assign a12876 = ~a12874 & a10304;
assign a12878 = ~a12876 & ~a12872;
assign a12880 = ~a12878 & ~a10302;
assign a12882 = a8620 & a8618;
assign a12884 = ~a12882 & a10302;
assign a12886 = ~a12884 & ~a12880;
assign a12888 = ~a12886 & ~a10300;
assign a12890 = a8380 & a8378;
assign a12892 = ~a12890 & a10300;
assign a12894 = ~a12892 & ~a12888;
assign a12896 = ~a12894 & a10292;
assign a12898 = ~a12896 & ~a12866;
assign a12900 = ~a12898 & ~a10288;
assign a12902 = a8140 & a8138;
assign a12904 = ~a12902 & a10306;
assign a12906 = a12904 & ~a10304;
assign a12908 = a7900 & a7898;
assign a12910 = ~a12908 & a10304;
assign a12912 = ~a12910 & ~a12906;
assign a12914 = ~a12912 & ~a10302;
assign a12916 = a7660 & a7658;
assign a12918 = ~a12916 & a10302;
assign a12920 = ~a12918 & ~a12914;
assign a12922 = ~a12920 & ~a10300;
assign a12924 = a7420 & a7418;
assign a12926 = ~a12924 & a10300;
assign a12928 = ~a12926 & ~a12922;
assign a12930 = ~a12928 & a10288;
assign a12932 = ~a12930 & ~a12900;
assign a12934 = a11022 & a11018;
assign a12936 = ~a12934 & a10546;
assign a12938 = a12936 & ~a10544;
assign a12940 = a10782 & a10778;
assign a12942 = ~a12940 & a10544;
assign a12944 = ~a12942 & ~a12938;
assign a12946 = ~a12944 & ~a10542;
assign a12948 = a10542 & ~a10538;
assign a12950 = ~a12948 & ~a12946;
assign a12952 = ~a12950 & ~a10540;
assign a12954 = a10302 & a10298;
assign a12956 = ~a12954 & a10540;
assign a12958 = ~a12956 & ~a12952;
assign a12960 = ~a12958 & a10538;
assign a12962 = a12960 & ~a10536;
assign a12964 = a10062 & a10058;
assign a12966 = ~a12964 & a10546;
assign a12968 = a12966 & ~a10544;
assign a12970 = a9822 & a9818;
assign a12972 = ~a12970 & a10544;
assign a12974 = ~a12972 & ~a12968;
assign a12976 = ~a12974 & ~a10542;
assign a12978 = a9582 & a9578;
assign a12980 = ~a12978 & a10542;
assign a12982 = ~a12980 & ~a12976;
assign a12984 = ~a12982 & ~a10540;
assign a12986 = a9342 & a9338;
assign a12988 = ~a12986 & a10540;
assign a12990 = ~a12988 & ~a12984;
assign a12992 = ~a12990 & a10536;
assign a12994 = ~a12992 & ~a12962;
assign a12996 = ~a12994 & ~a10532;
assign a12998 = a9102 & a9098;
assign a13000 = ~a12998 & a10546;
assign a13002 = a13000 & ~a10544;
assign a13004 = a8862 & a8858;
assign a13006 = ~a13004 & a10544;
assign a13008 = ~a13006 & ~a13002;
assign a13010 = ~a13008 & ~a10542;
assign a13012 = a8622 & a8618;
assign a13014 = ~a13012 & a10542;
assign a13016 = ~a13014 & ~a13010;
assign a13018 = ~a13016 & ~a10540;
assign a13020 = a8382 & a8378;
assign a13022 = ~a13020 & a10540;
assign a13024 = ~a13022 & ~a13018;
assign a13026 = ~a13024 & a10532;
assign a13028 = ~a13026 & ~a12996;
assign a13030 = ~a13028 & ~a10528;
assign a13032 = a8142 & a8138;
assign a13034 = ~a13032 & a10546;
assign a13036 = a13034 & ~a10544;
assign a13038 = a7902 & a7898;
assign a13040 = ~a13038 & a10544;
assign a13042 = ~a13040 & ~a13036;
assign a13044 = ~a13042 & ~a10542;
assign a13046 = a7662 & a7658;
assign a13048 = ~a13046 & a10542;
assign a13050 = ~a13048 & ~a13044;
assign a13052 = ~a13050 & ~a10540;
assign a13054 = a7422 & a7418;
assign a13056 = ~a13054 & a10540;
assign a13058 = ~a13056 & ~a13052;
assign a13060 = ~a13058 & a10528;
assign a13062 = ~a13060 & ~a13030;
assign a13064 = a11024 & a11018;
assign a13066 = ~a13064 & a10786;
assign a13068 = a13066 & ~a10784;
assign a13070 = a10784 & ~a10778;
assign a13072 = ~a13070 & ~a13068;
assign a13074 = ~a13072 & ~a10782;
assign a13076 = a10544 & a10538;
assign a13078 = ~a13076 & a10782;
assign a13080 = ~a13078 & ~a13074;
assign a13082 = ~a13080 & ~a10780;
assign a13084 = a10304 & a10298;
assign a13086 = ~a13084 & a10780;
assign a13088 = ~a13086 & ~a13082;
assign a13090 = ~a13088 & a10778;
assign a13092 = a13090 & ~a10776;
assign a13094 = a10064 & a10058;
assign a13096 = ~a13094 & a10786;
assign a13098 = a13096 & ~a10784;
assign a13100 = a9824 & a9818;
assign a13102 = ~a13100 & a10784;
assign a13104 = ~a13102 & ~a13098;
assign a13106 = ~a13104 & ~a10782;
assign a13108 = a9584 & a9578;
assign a13110 = ~a13108 & a10782;
assign a13112 = ~a13110 & ~a13106;
assign a13114 = ~a13112 & ~a10780;
assign a13116 = a9344 & a9338;
assign a13118 = ~a13116 & a10780;
assign a13120 = ~a13118 & ~a13114;
assign a13122 = ~a13120 & a10776;
assign a13124 = ~a13122 & ~a13092;
assign a13126 = ~a13124 & ~a10772;
assign a13128 = a9104 & a9098;
assign a13130 = ~a13128 & a10786;
assign a13132 = a13130 & ~a10784;
assign a13134 = a8864 & a8858;
assign a13136 = ~a13134 & a10784;
assign a13138 = ~a13136 & ~a13132;
assign a13140 = ~a13138 & ~a10782;
assign a13142 = a8624 & a8618;
assign a13144 = ~a13142 & a10782;
assign a13146 = ~a13144 & ~a13140;
assign a13148 = ~a13146 & ~a10780;
assign a13150 = a8384 & a8378;
assign a13152 = ~a13150 & a10780;
assign a13154 = ~a13152 & ~a13148;
assign a13156 = ~a13154 & a10772;
assign a13158 = ~a13156 & ~a13126;
assign a13160 = ~a13158 & ~a10768;
assign a13162 = a8144 & a8138;
assign a13164 = ~a13162 & a10786;
assign a13166 = a13164 & ~a10784;
assign a13168 = a7904 & a7898;
assign a13170 = ~a13168 & a10784;
assign a13172 = ~a13170 & ~a13166;
assign a13174 = ~a13172 & ~a10782;
assign a13176 = a7664 & a7658;
assign a13178 = ~a13176 & a10782;
assign a13180 = ~a13178 & ~a13174;
assign a13182 = ~a13180 & ~a10780;
assign a13184 = a7424 & a7418;
assign a13186 = ~a13184 & a10780;
assign a13188 = ~a13186 & ~a13182;
assign a13190 = ~a13188 & a10768;
assign a13192 = ~a13190 & ~a13160;
assign a13194 = a11026 & ~a11018;
assign a13196 = a13194 & ~a11024;
assign a13198 = a10786 & a10778;
assign a13200 = ~a13198 & a11024;
assign a13202 = ~a13200 & ~a13196;
assign a13204 = ~a13202 & ~a11022;
assign a13206 = a10546 & a10538;
assign a13208 = ~a13206 & a11022;
assign a13210 = ~a13208 & ~a13204;
assign a13212 = ~a13210 & ~a11020;
assign a13214 = a10306 & a10298;
assign a13216 = ~a13214 & a11020;
assign a13218 = ~a13216 & ~a13212;
assign a13220 = ~a13218 & a11018;
assign a13222 = a13220 & ~a11016;
assign a13224 = a10066 & a10058;
assign a13226 = ~a13224 & a11026;
assign a13228 = a13226 & ~a11024;
assign a13230 = a9826 & a9818;
assign a13232 = ~a13230 & a11024;
assign a13234 = ~a13232 & ~a13228;
assign a13236 = ~a13234 & ~a11022;
assign a13238 = a9586 & a9578;
assign a13240 = ~a13238 & a11022;
assign a13242 = ~a13240 & ~a13236;
assign a13244 = ~a13242 & ~a11020;
assign a13246 = a9346 & a9338;
assign a13248 = ~a13246 & a11020;
assign a13250 = ~a13248 & ~a13244;
assign a13252 = ~a13250 & a11016;
assign a13254 = ~a13252 & ~a13222;
assign a13256 = ~a13254 & ~a11012;
assign a13258 = a9106 & a9098;
assign a13260 = ~a13258 & a11026;
assign a13262 = a13260 & ~a11024;
assign a13264 = a8866 & a8858;
assign a13266 = ~a13264 & a11024;
assign a13268 = ~a13266 & ~a13262;
assign a13270 = ~a13268 & ~a11022;
assign a13272 = a8626 & a8618;
assign a13274 = ~a13272 & a11022;
assign a13276 = ~a13274 & ~a13270;
assign a13278 = ~a13276 & ~a11020;
assign a13280 = a8386 & a8378;
assign a13282 = ~a13280 & a11020;
assign a13284 = ~a13282 & ~a13278;
assign a13286 = ~a13284 & a11012;
assign a13288 = ~a13286 & ~a13256;
assign a13290 = ~a13288 & ~a11008;
assign a13292 = a8146 & a8138;
assign a13294 = ~a13292 & a11026;
assign a13296 = a13294 & ~a11024;
assign a13298 = a7906 & a7898;
assign a13300 = ~a13298 & a11024;
assign a13302 = ~a13300 & ~a13296;
assign a13304 = ~a13302 & ~a11022;
assign a13306 = a7666 & a7658;
assign a13308 = ~a13306 & a11022;
assign a13310 = ~a13308 & ~a13304;
assign a13312 = ~a13310 & ~a11020;
assign a13314 = a7426 & a7418;
assign a13316 = ~a13314 & a11020;
assign a13318 = ~a13316 & ~a13312;
assign a13320 = ~a13318 & a11008;
assign a13322 = ~a13320 & ~a13290;
assign a13324 = ~a8380 & a8368;
assign a13326 = ~a8620 & a8608;
assign a13328 = ~a13326 & ~a13324;
assign a13330 = ~a8860 & a8848;
assign a13332 = ~a13330 & a13328;
assign a13334 = ~a9100 & a9088;
assign a13336 = ~a13334 & a13332;
assign a13338 = ~a9340 & a9328;
assign a13340 = ~a8616 & ~a8376;
assign a13342 = a13340 & ~a8856;
assign a13344 = a13342 & ~a9096;
assign a13346 = ~a8618 & ~a8378;
assign a13348 = a13346 & ~a8858;
assign a13350 = a13348 & ~a9098;
assign a13352 = ~a10536 & ~a10296;
assign a13354 = a13352 & ~a10776;
assign a13356 = a13354 & ~a11016;
assign a13358 = ~a13356 & ~a13350;
assign a13360 = ~a13358 & a13344;
assign a13362 = ~a13360 & a13338;
assign a13364 = ~a9580 & a9568;
assign a13366 = a13364 & ~a13360;
assign a13368 = ~a9820 & a9808;
assign a13370 = a13368 & ~a13360;
assign a13372 = ~a10060 & a10048;
assign a13374 = a13372 & ~a13360;
assign a13376 = ~a10300 & a10288;
assign a13378 = ~a9578 & ~a9338;
assign a13380 = a13378 & ~a9818;
assign a13382 = a13380 & ~a10058;
assign a13384 = ~a13382 & ~a13344;
assign a13386 = ~a13384 & a13350;
assign a13388 = ~a13386 & a13376;
assign a13390 = ~a10540 & a10528;
assign a13392 = a13390 & ~a13386;
assign a13394 = ~a10780 & a10768;
assign a13396 = a13394 & ~a13386;
assign a13398 = ~a11020 & a11008;
assign a13400 = a13398 & ~a13386;
assign a13402 = ~a13400 & ~a13396;
assign a13404 = a13402 & ~a13392;
assign a13406 = a13404 & ~a13388;
assign a13408 = a13406 & ~a13374;
assign a13410 = a13408 & ~a13370;
assign a13412 = a13410 & ~a13366;
assign a13414 = a13412 & ~a13362;
assign a13416 = a13414 & a13336;
assign a13418 = ~a13416 & a7412;
assign a13420 = ~a8382 & a8368;
assign a13422 = ~a8622 & a8608;
assign a13424 = ~a13422 & ~a13420;
assign a13426 = ~a8862 & a8848;
assign a13428 = ~a13426 & a13424;
assign a13430 = ~a9102 & a9088;
assign a13432 = ~a13430 & a13428;
assign a13434 = ~a9342 & a9328;
assign a13436 = a13434 & ~a13360;
assign a13438 = ~a9582 & a9568;
assign a13440 = a13438 & ~a13360;
assign a13442 = ~a9822 & a9808;
assign a13444 = a13442 & ~a13360;
assign a13446 = ~a10062 & a10048;
assign a13448 = a13446 & ~a13360;
assign a13450 = ~a10302 & a10288;
assign a13452 = a13450 & ~a13386;
assign a13454 = ~a10542 & a10528;
assign a13456 = a13454 & ~a13386;
assign a13458 = ~a10782 & a10768;
assign a13460 = a13458 & ~a13386;
assign a13462 = ~a11022 & a11008;
assign a13464 = a13462 & ~a13386;
assign a13466 = ~a13464 & ~a13460;
assign a13468 = a13466 & ~a13456;
assign a13470 = a13468 & ~a13452;
assign a13472 = a13470 & ~a13448;
assign a13474 = a13472 & ~a13444;
assign a13476 = a13474 & ~a13440;
assign a13478 = a13476 & ~a13436;
assign a13480 = a13478 & a13432;
assign a13482 = ~a13480 & a7652;
assign a13484 = ~a8384 & a8368;
assign a13486 = ~a8624 & a8608;
assign a13488 = ~a13486 & ~a13484;
assign a13490 = ~a8864 & a8848;
assign a13492 = ~a13490 & a13488;
assign a13494 = ~a9104 & a9088;
assign a13496 = ~a13494 & a13492;
assign a13498 = ~a9344 & a9328;
assign a13500 = a13498 & ~a13360;
assign a13502 = ~a9584 & a9568;
assign a13504 = a13502 & ~a13360;
assign a13506 = ~a9824 & a9808;
assign a13508 = a13506 & ~a13360;
assign a13510 = ~a10064 & a10048;
assign a13512 = a13510 & ~a13360;
assign a13514 = ~a10304 & a10288;
assign a13516 = a13514 & ~a13386;
assign a13518 = ~a10544 & a10528;
assign a13520 = a13518 & ~a13386;
assign a13522 = ~a10784 & a10768;
assign a13524 = a13522 & ~a13386;
assign a13526 = ~a11024 & a11008;
assign a13528 = a13526 & ~a13386;
assign a13530 = ~a13528 & ~a13524;
assign a13532 = a13530 & ~a13520;
assign a13534 = a13532 & ~a13516;
assign a13536 = a13534 & ~a13512;
assign a13538 = a13536 & ~a13508;
assign a13540 = a13538 & ~a13504;
assign a13542 = a13540 & ~a13500;
assign a13544 = a13542 & a13496;
assign a13546 = ~a13544 & a7892;
assign a13548 = ~a8386 & a8368;
assign a13550 = ~a8626 & a8608;
assign a13552 = ~a13550 & ~a13548;
assign a13554 = ~a8866 & a8848;
assign a13556 = ~a13554 & a13552;
assign a13558 = ~a9106 & a9088;
assign a13560 = ~a13558 & a13556;
assign a13562 = ~a9346 & a9328;
assign a13564 = a13562 & ~a13360;
assign a13566 = ~a9586 & a9568;
assign a13568 = a13566 & ~a13360;
assign a13570 = ~a9826 & a9808;
assign a13572 = a13570 & ~a13360;
assign a13574 = ~a10066 & a10048;
assign a13576 = a13574 & ~a13360;
assign a13578 = ~a10306 & a10288;
assign a13580 = a13578 & ~a13386;
assign a13582 = ~a10546 & a10528;
assign a13584 = a13582 & ~a13386;
assign a13586 = ~a10786 & a10768;
assign a13588 = a13586 & ~a13386;
assign a13590 = ~a11026 & a11008;
assign a13592 = a13590 & ~a13386;
assign a13594 = ~a13592 & ~a13588;
assign a13596 = a13594 & ~a13584;
assign a13598 = a13596 & ~a13580;
assign a13600 = a13598 & ~a13576;
assign a13602 = a13600 & ~a13572;
assign a13604 = a13602 & ~a13568;
assign a13606 = a13604 & ~a13564;
assign a13608 = a13606 & a13560;
assign a13610 = ~a13608 & a8132;
assign a13612 = ~a9572 & ~a9332;
assign a13614 = a13612 & ~a9812;
assign a13616 = a13614 & ~a10052;
assign a13618 = ~a10532 & ~a10292;
assign a13620 = a13618 & ~a10772;
assign a13622 = a13620 & ~a11012;
assign a13624 = ~a13622 & ~a13382;
assign a13626 = ~a13624 & a13616;
assign a13628 = ~a13626 & ~a13336;
assign a13630 = ~a13616 & ~a13350;
assign a13632 = ~a13630 & a13382;
assign a13634 = ~a13632 & a13376;
assign a13636 = ~a13632 & a13390;
assign a13638 = ~a13632 & a13394;
assign a13640 = ~a13632 & a13398;
assign a13642 = ~a13640 & ~a13638;
assign a13644 = a13642 & ~a13636;
assign a13646 = a13644 & ~a13634;
assign a13648 = a13646 & ~a13628;
assign a13650 = a13648 & ~a13338;
assign a13652 = a13650 & ~a13364;
assign a13654 = a13652 & ~a13368;
assign a13656 = a13654 & ~a13372;
assign a13658 = ~a13656 & a7416;
assign a13660 = ~a13626 & ~a13432;
assign a13662 = ~a13632 & a13450;
assign a13664 = ~a13632 & a13454;
assign a13666 = ~a13632 & a13458;
assign a13668 = ~a13632 & a13462;
assign a13670 = ~a13668 & ~a13666;
assign a13672 = a13670 & ~a13664;
assign a13674 = a13672 & ~a13662;
assign a13676 = a13674 & ~a13660;
assign a13678 = a13676 & ~a13434;
assign a13680 = a13678 & ~a13438;
assign a13682 = a13680 & ~a13442;
assign a13684 = a13682 & ~a13446;
assign a13686 = ~a13684 & a7656;
assign a13688 = ~a13626 & ~a13496;
assign a13690 = ~a13632 & a13514;
assign a13692 = ~a13632 & a13518;
assign a13694 = ~a13632 & a13522;
assign a13696 = ~a13632 & a13526;
assign a13698 = ~a13696 & ~a13694;
assign a13700 = a13698 & ~a13692;
assign a13702 = a13700 & ~a13690;
assign a13704 = a13702 & ~a13688;
assign a13706 = a13704 & ~a13498;
assign a13708 = a13706 & ~a13502;
assign a13710 = a13708 & ~a13506;
assign a13712 = a13710 & ~a13510;
assign a13714 = ~a13712 & a7896;
assign a13716 = ~a13626 & ~a13560;
assign a13718 = ~a13632 & a13578;
assign a13720 = ~a13632 & a13582;
assign a13722 = ~a13632 & a13586;
assign a13724 = ~a13632 & a13590;
assign a13726 = ~a13724 & ~a13722;
assign a13728 = a13726 & ~a13720;
assign a13730 = a13728 & ~a13718;
assign a13732 = a13730 & ~a13716;
assign a13734 = a13732 & ~a13562;
assign a13736 = a13734 & ~a13566;
assign a13738 = a13736 & ~a13570;
assign a13740 = a13738 & ~a13574;
assign a13742 = ~a13740 & a8136;
assign a13744 = ~a13616 & ~a13356;
assign a13746 = ~a13744 & a13622;
assign a13748 = ~a13746 & ~a13336;
assign a13750 = ~a13622 & ~a13344;
assign a13752 = ~a13750 & a13356;
assign a13754 = ~a13752 & a13338;
assign a13756 = ~a13752 & a13364;
assign a13758 = ~a13752 & a13368;
assign a13760 = ~a13752 & a13372;
assign a13762 = ~a13760 & ~a13758;
assign a13764 = a13762 & ~a13756;
assign a13766 = a13764 & ~a13754;
assign a13768 = a13766 & ~a13748;
assign a13770 = a13768 & ~a13376;
assign a13772 = a13770 & ~a13390;
assign a13774 = a13772 & ~a13394;
assign a13776 = a13774 & ~a13398;
assign a13778 = ~a13776 & a7418;
assign a13780 = ~a13746 & ~a13432;
assign a13782 = ~a13752 & a13434;
assign a13784 = ~a13752 & a13438;
assign a13786 = ~a13752 & a13442;
assign a13788 = ~a13752 & a13446;
assign a13790 = ~a13788 & ~a13786;
assign a13792 = a13790 & ~a13784;
assign a13794 = a13792 & ~a13782;
assign a13796 = a13794 & ~a13780;
assign a13798 = a13796 & ~a13450;
assign a13800 = a13798 & ~a13454;
assign a13802 = a13800 & ~a13458;
assign a13804 = a13802 & ~a13462;
assign a13806 = ~a13804 & a7658;
assign a13808 = ~a13746 & ~a13496;
assign a13810 = ~a13752 & a13498;
assign a13812 = ~a13752 & a13502;
assign a13814 = ~a13752 & a13506;
assign a13816 = ~a13752 & a13510;
assign a13818 = ~a13816 & ~a13814;
assign a13820 = a13818 & ~a13812;
assign a13822 = a13820 & ~a13810;
assign a13824 = a13822 & ~a13808;
assign a13826 = a13824 & ~a13514;
assign a13828 = a13826 & ~a13518;
assign a13830 = a13828 & ~a13522;
assign a13832 = a13830 & ~a13526;
assign a13834 = ~a13832 & a7898;
assign a13836 = ~a13746 & ~a13560;
assign a13838 = ~a13752 & a13562;
assign a13840 = ~a13752 & a13566;
assign a13842 = ~a13752 & a13570;
assign a13844 = ~a13752 & a13574;
assign a13846 = ~a13844 & ~a13842;
assign a13848 = a13846 & ~a13840;
assign a13850 = a13848 & ~a13838;
assign a13852 = a13850 & ~a13836;
assign a13854 = a13852 & ~a13578;
assign a13856 = a13854 & ~a13582;
assign a13858 = a13856 & ~a13586;
assign a13860 = a13858 & ~a13590;
assign a13862 = ~a13860 & a8138;
assign a13864 = ~a7420 & a7412;
assign a13866 = ~a7660 & a7652;
assign a13868 = ~a13866 & ~a13864;
assign a13870 = ~a7900 & a7892;
assign a13872 = ~a13870 & a13868;
assign a13874 = ~a8140 & a8132;
assign a13876 = ~a13874 & a13872;
assign a13878 = ~a9340 & a9332;
assign a13880 = ~a7656 & ~a7416;
assign a13882 = a13880 & ~a7896;
assign a13884 = a13882 & ~a8136;
assign a13886 = ~a7658 & ~a7418;
assign a13888 = a13886 & ~a7898;
assign a13890 = a13888 & ~a8138;
assign a13892 = ~a13890 & ~a13356;
assign a13894 = ~a13892 & a13884;
assign a13896 = ~a13894 & a13878;
assign a13898 = ~a9580 & a9572;
assign a13900 = a13898 & ~a13894;
assign a13902 = ~a9820 & a9812;
assign a13904 = a13902 & ~a13894;
assign a13906 = ~a10060 & a10052;
assign a13908 = a13906 & ~a13894;
assign a13910 = ~a10300 & a10292;
assign a13912 = ~a13884 & ~a13382;
assign a13914 = ~a13912 & a13890;
assign a13916 = ~a13914 & a13910;
assign a13918 = ~a10540 & a10532;
assign a13920 = a13918 & ~a13914;
assign a13922 = ~a10780 & a10772;
assign a13924 = a13922 & ~a13914;
assign a13926 = ~a11020 & a11012;
assign a13928 = a13926 & ~a13914;
assign a13930 = ~a13928 & ~a13924;
assign a13932 = a13930 & ~a13920;
assign a13934 = a13932 & ~a13916;
assign a13936 = a13934 & ~a13908;
assign a13938 = a13936 & ~a13904;
assign a13940 = a13938 & ~a13900;
assign a13942 = a13940 & ~a13896;
assign a13944 = a13942 & a13876;
assign a13946 = ~a13944 & a8368;
assign a13948 = ~a7422 & a7412;
assign a13950 = ~a7662 & a7652;
assign a13952 = ~a13950 & ~a13948;
assign a13954 = ~a7902 & a7892;
assign a13956 = ~a13954 & a13952;
assign a13958 = ~a8142 & a8132;
assign a13960 = ~a13958 & a13956;
assign a13962 = ~a9342 & a9332;
assign a13964 = a13962 & ~a13894;
assign a13966 = ~a9582 & a9572;
assign a13968 = a13966 & ~a13894;
assign a13970 = ~a9822 & a9812;
assign a13972 = a13970 & ~a13894;
assign a13974 = ~a10062 & a10052;
assign a13976 = a13974 & ~a13894;
assign a13978 = ~a10302 & a10292;
assign a13980 = a13978 & ~a13914;
assign a13982 = ~a10542 & a10532;
assign a13984 = a13982 & ~a13914;
assign a13986 = ~a10782 & a10772;
assign a13988 = a13986 & ~a13914;
assign a13990 = ~a11022 & a11012;
assign a13992 = a13990 & ~a13914;
assign a13994 = ~a13992 & ~a13988;
assign a13996 = a13994 & ~a13984;
assign a13998 = a13996 & ~a13980;
assign a14000 = a13998 & ~a13976;
assign a14002 = a14000 & ~a13972;
assign a14004 = a14002 & ~a13968;
assign a14006 = a14004 & ~a13964;
assign a14008 = a14006 & a13960;
assign a14010 = ~a14008 & a8608;
assign a14012 = ~a7424 & a7412;
assign a14014 = ~a7664 & a7652;
assign a14016 = ~a14014 & ~a14012;
assign a14018 = ~a7904 & a7892;
assign a14020 = ~a14018 & a14016;
assign a14022 = ~a8144 & a8132;
assign a14024 = ~a14022 & a14020;
assign a14026 = ~a9344 & a9332;
assign a14028 = a14026 & ~a13894;
assign a14030 = ~a9584 & a9572;
assign a14032 = a14030 & ~a13894;
assign a14034 = ~a9824 & a9812;
assign a14036 = a14034 & ~a13894;
assign a14038 = ~a10064 & a10052;
assign a14040 = a14038 & ~a13894;
assign a14042 = ~a10304 & a10292;
assign a14044 = a14042 & ~a13914;
assign a14046 = ~a10544 & a10532;
assign a14048 = a14046 & ~a13914;
assign a14050 = ~a10784 & a10772;
assign a14052 = a14050 & ~a13914;
assign a14054 = ~a11024 & a11012;
assign a14056 = a14054 & ~a13914;
assign a14058 = ~a14056 & ~a14052;
assign a14060 = a14058 & ~a14048;
assign a14062 = a14060 & ~a14044;
assign a14064 = a14062 & ~a14040;
assign a14066 = a14064 & ~a14036;
assign a14068 = a14066 & ~a14032;
assign a14070 = a14068 & ~a14028;
assign a14072 = a14070 & a14024;
assign a14074 = ~a14072 & a8848;
assign a14076 = ~a7426 & a7412;
assign a14078 = ~a7666 & a7652;
assign a14080 = ~a14078 & ~a14076;
assign a14082 = ~a7906 & a7892;
assign a14084 = ~a14082 & a14080;
assign a14086 = ~a8146 & a8132;
assign a14088 = ~a14086 & a14084;
assign a14090 = ~a9346 & a9332;
assign a14092 = a14090 & ~a13894;
assign a14094 = ~a9586 & a9572;
assign a14096 = a14094 & ~a13894;
assign a14098 = ~a9826 & a9812;
assign a14100 = a14098 & ~a13894;
assign a14102 = ~a10066 & a10052;
assign a14104 = a14102 & ~a13894;
assign a14106 = ~a10306 & a10292;
assign a14108 = a14106 & ~a13914;
assign a14110 = ~a10546 & a10532;
assign a14112 = a14110 & ~a13914;
assign a14114 = ~a10786 & a10772;
assign a14116 = a14114 & ~a13914;
assign a14118 = ~a11026 & a11012;
assign a14120 = a14118 & ~a13914;
assign a14122 = ~a14120 & ~a14116;
assign a14124 = a14122 & ~a14112;
assign a14126 = a14124 & ~a14108;
assign a14128 = a14126 & ~a14104;
assign a14130 = a14128 & ~a14100;
assign a14132 = a14130 & ~a14096;
assign a14134 = a14132 & ~a14092;
assign a14136 = a14134 & a14088;
assign a14138 = ~a14136 & a9088;
assign a14140 = ~a9568 & ~a9328;
assign a14142 = a14140 & ~a9808;
assign a14144 = a14142 & ~a10048;
assign a14146 = ~a10528 & ~a10288;
assign a14148 = a14146 & ~a10768;
assign a14150 = a14148 & ~a11008;
assign a14152 = ~a14150 & ~a13382;
assign a14154 = ~a14152 & a14144;
assign a14156 = ~a14154 & ~a13876;
assign a14158 = ~a14144 & ~a13890;
assign a14160 = ~a14158 & a13382;
assign a14162 = ~a14160 & a13910;
assign a14164 = ~a14160 & a13918;
assign a14166 = ~a14160 & a13922;
assign a14168 = ~a14160 & a13926;
assign a14170 = ~a14168 & ~a14166;
assign a14172 = a14170 & ~a14164;
assign a14174 = a14172 & ~a14162;
assign a14176 = a14174 & ~a14156;
assign a14178 = a14176 & ~a13878;
assign a14180 = a14178 & ~a13898;
assign a14182 = a14180 & ~a13902;
assign a14184 = a14182 & ~a13906;
assign a14186 = ~a14184 & a8376;
assign a14188 = ~a14154 & ~a13960;
assign a14190 = ~a14160 & a13978;
assign a14192 = ~a14160 & a13982;
assign a14194 = ~a14160 & a13986;
assign a14196 = ~a14160 & a13990;
assign a14198 = ~a14196 & ~a14194;
assign a14200 = a14198 & ~a14192;
assign a14202 = a14200 & ~a14190;
assign a14204 = a14202 & ~a14188;
assign a14206 = a14204 & ~a13962;
assign a14208 = a14206 & ~a13966;
assign a14210 = a14208 & ~a13970;
assign a14212 = a14210 & ~a13974;
assign a14214 = ~a14212 & a8616;
assign a14216 = ~a14154 & ~a14024;
assign a14218 = ~a14160 & a14042;
assign a14220 = ~a14160 & a14046;
assign a14222 = ~a14160 & a14050;
assign a14224 = ~a14160 & a14054;
assign a14226 = ~a14224 & ~a14222;
assign a14228 = a14226 & ~a14220;
assign a14230 = a14228 & ~a14218;
assign a14232 = a14230 & ~a14216;
assign a14234 = a14232 & ~a14026;
assign a14236 = a14234 & ~a14030;
assign a14238 = a14236 & ~a14034;
assign a14240 = a14238 & ~a14038;
assign a14242 = ~a14240 & a8856;
assign a14244 = ~a14154 & ~a14088;
assign a14246 = ~a14160 & a14106;
assign a14248 = ~a14160 & a14110;
assign a14250 = ~a14160 & a14114;
assign a14252 = ~a14160 & a14118;
assign a14254 = ~a14252 & ~a14250;
assign a14256 = a14254 & ~a14248;
assign a14258 = a14256 & ~a14246;
assign a14260 = a14258 & ~a14244;
assign a14262 = a14260 & ~a14090;
assign a14264 = a14262 & ~a14094;
assign a14266 = a14264 & ~a14098;
assign a14268 = a14266 & ~a14102;
assign a14270 = ~a14268 & a9096;
assign a14272 = ~a14144 & ~a13356;
assign a14274 = ~a14272 & a14150;
assign a14276 = ~a14274 & ~a13876;
assign a14278 = ~a14150 & ~a13884;
assign a14280 = ~a14278 & a13356;
assign a14282 = ~a14280 & a13878;
assign a14284 = ~a14280 & a13898;
assign a14286 = ~a14280 & a13902;
assign a14288 = ~a14280 & a13906;
assign a14290 = ~a14288 & ~a14286;
assign a14292 = a14290 & ~a14284;
assign a14294 = a14292 & ~a14282;
assign a14296 = a14294 & ~a14276;
assign a14298 = a14296 & ~a13910;
assign a14300 = a14298 & ~a13918;
assign a14302 = a14300 & ~a13922;
assign a14304 = a14302 & ~a13926;
assign a14306 = ~a14304 & a8378;
assign a14308 = ~a14274 & ~a13960;
assign a14310 = ~a14280 & a13962;
assign a14312 = ~a14280 & a13966;
assign a14314 = ~a14280 & a13970;
assign a14316 = ~a14280 & a13974;
assign a14318 = ~a14316 & ~a14314;
assign a14320 = a14318 & ~a14312;
assign a14322 = a14320 & ~a14310;
assign a14324 = a14322 & ~a14308;
assign a14326 = a14324 & ~a13978;
assign a14328 = a14326 & ~a13982;
assign a14330 = a14328 & ~a13986;
assign a14332 = a14330 & ~a13990;
assign a14334 = ~a14332 & a8618;
assign a14336 = ~a14274 & ~a14024;
assign a14338 = ~a14280 & a14026;
assign a14340 = ~a14280 & a14030;
assign a14342 = ~a14280 & a14034;
assign a14344 = ~a14280 & a14038;
assign a14346 = ~a14344 & ~a14342;
assign a14348 = a14346 & ~a14340;
assign a14350 = a14348 & ~a14338;
assign a14352 = a14350 & ~a14336;
assign a14354 = a14352 & ~a14042;
assign a14356 = a14354 & ~a14046;
assign a14358 = a14356 & ~a14050;
assign a14360 = a14358 & ~a14054;
assign a14362 = ~a14360 & a8858;
assign a14364 = ~a14274 & ~a14088;
assign a14366 = ~a14280 & a14090;
assign a14368 = ~a14280 & a14094;
assign a14370 = ~a14280 & a14098;
assign a14372 = ~a14280 & a14102;
assign a14374 = ~a14372 & ~a14370;
assign a14376 = a14374 & ~a14368;
assign a14378 = a14376 & ~a14366;
assign a14380 = a14378 & ~a14364;
assign a14382 = a14380 & ~a14106;
assign a14384 = a14382 & ~a14110;
assign a14386 = a14384 & ~a14114;
assign a14388 = a14386 & ~a14118;
assign a14390 = ~a14388 & a9098;
assign a14392 = ~a7420 & a7416;
assign a14394 = ~a7660 & a7656;
assign a14396 = ~a14394 & ~a14392;
assign a14398 = ~a7900 & a7896;
assign a14400 = ~a14398 & a14396;
assign a14402 = ~a8140 & a8136;
assign a14404 = ~a14402 & a14400;
assign a14406 = ~a8380 & a8376;
assign a14408 = ~a7652 & ~a7412;
assign a14410 = a14408 & ~a7892;
assign a14412 = a14410 & ~a8132;
assign a14414 = ~a13890 & ~a13622;
assign a14416 = ~a14414 & a14412;
assign a14418 = ~a14416 & a14406;
assign a14420 = ~a8620 & a8616;
assign a14422 = a14420 & ~a14416;
assign a14424 = ~a8860 & a8856;
assign a14426 = a14424 & ~a14416;
assign a14428 = ~a9100 & a9096;
assign a14430 = a14428 & ~a14416;
assign a14432 = ~a10300 & a10296;
assign a14434 = ~a14412 & ~a13350;
assign a14436 = ~a14434 & a13890;
assign a14438 = ~a14436 & a14432;
assign a14440 = ~a10540 & a10536;
assign a14442 = a14440 & ~a14436;
assign a14444 = ~a10780 & a10776;
assign a14446 = a14444 & ~a14436;
assign a14448 = ~a11020 & a11016;
assign a14450 = a14448 & ~a14436;
assign a14452 = ~a14450 & ~a14446;
assign a14454 = a14452 & ~a14442;
assign a14456 = a14454 & ~a14438;
assign a14458 = a14456 & ~a14430;
assign a14460 = a14458 & ~a14426;
assign a14462 = a14460 & ~a14422;
assign a14464 = a14462 & ~a14418;
assign a14466 = a14464 & a14404;
assign a14468 = ~a14466 & a9328;
assign a14470 = ~a7422 & a7416;
assign a14472 = ~a7662 & a7656;
assign a14474 = ~a14472 & ~a14470;
assign a14476 = ~a7902 & a7896;
assign a14478 = ~a14476 & a14474;
assign a14480 = ~a8142 & a8136;
assign a14482 = ~a14480 & a14478;
assign a14484 = ~a8382 & a8376;
assign a14486 = a14484 & ~a14416;
assign a14488 = ~a8622 & a8616;
assign a14490 = a14488 & ~a14416;
assign a14492 = ~a8862 & a8856;
assign a14494 = a14492 & ~a14416;
assign a14496 = ~a9102 & a9096;
assign a14498 = a14496 & ~a14416;
assign a14500 = ~a10302 & a10296;
assign a14502 = a14500 & ~a14436;
assign a14504 = ~a10542 & a10536;
assign a14506 = a14504 & ~a14436;
assign a14508 = ~a10782 & a10776;
assign a14510 = a14508 & ~a14436;
assign a14512 = ~a11022 & a11016;
assign a14514 = a14512 & ~a14436;
assign a14516 = ~a14514 & ~a14510;
assign a14518 = a14516 & ~a14506;
assign a14520 = a14518 & ~a14502;
assign a14522 = a14520 & ~a14498;
assign a14524 = a14522 & ~a14494;
assign a14526 = a14524 & ~a14490;
assign a14528 = a14526 & ~a14486;
assign a14530 = a14528 & a14482;
assign a14532 = ~a14530 & a9568;
assign a14534 = ~a7424 & a7416;
assign a14536 = ~a7664 & a7656;
assign a14538 = ~a14536 & ~a14534;
assign a14540 = ~a7904 & a7896;
assign a14542 = ~a14540 & a14538;
assign a14544 = ~a8144 & a8136;
assign a14546 = ~a14544 & a14542;
assign a14548 = ~a8384 & a8376;
assign a14550 = a14548 & ~a14416;
assign a14552 = ~a8624 & a8616;
assign a14554 = a14552 & ~a14416;
assign a14556 = ~a8864 & a8856;
assign a14558 = a14556 & ~a14416;
assign a14560 = ~a9104 & a9096;
assign a14562 = a14560 & ~a14416;
assign a14564 = ~a10304 & a10296;
assign a14566 = a14564 & ~a14436;
assign a14568 = ~a10544 & a10536;
assign a14570 = a14568 & ~a14436;
assign a14572 = ~a10784 & a10776;
assign a14574 = a14572 & ~a14436;
assign a14576 = ~a11024 & a11016;
assign a14578 = a14576 & ~a14436;
assign a14580 = ~a14578 & ~a14574;
assign a14582 = a14580 & ~a14570;
assign a14584 = a14582 & ~a14566;
assign a14586 = a14584 & ~a14562;
assign a14588 = a14586 & ~a14558;
assign a14590 = a14588 & ~a14554;
assign a14592 = a14590 & ~a14550;
assign a14594 = a14592 & a14546;
assign a14596 = ~a14594 & a9808;
assign a14598 = ~a7426 & a7416;
assign a14600 = ~a7666 & a7656;
assign a14602 = ~a14600 & ~a14598;
assign a14604 = ~a7906 & a7896;
assign a14606 = ~a14604 & a14602;
assign a14608 = ~a8146 & a8136;
assign a14610 = ~a14608 & a14606;
assign a14612 = ~a8386 & a8376;
assign a14614 = a14612 & ~a14416;
assign a14616 = ~a8626 & a8616;
assign a14618 = a14616 & ~a14416;
assign a14620 = ~a8866 & a8856;
assign a14622 = a14620 & ~a14416;
assign a14624 = ~a9106 & a9096;
assign a14626 = a14624 & ~a14416;
assign a14628 = ~a10306 & a10296;
assign a14630 = a14628 & ~a14436;
assign a14632 = ~a10546 & a10536;
assign a14634 = a14632 & ~a14436;
assign a14636 = ~a10786 & a10776;
assign a14638 = a14636 & ~a14436;
assign a14640 = ~a11026 & a11016;
assign a14642 = a14640 & ~a14436;
assign a14644 = ~a14642 & ~a14638;
assign a14646 = a14644 & ~a14634;
assign a14648 = a14646 & ~a14630;
assign a14650 = a14648 & ~a14626;
assign a14652 = a14650 & ~a14622;
assign a14654 = a14652 & ~a14618;
assign a14656 = a14654 & ~a14614;
assign a14658 = a14656 & a14610;
assign a14660 = ~a14658 & a10048;
assign a14662 = ~a8608 & ~a8368;
assign a14664 = a14662 & ~a8848;
assign a14666 = a14664 & ~a9088;
assign a14668 = ~a14150 & ~a13350;
assign a14670 = ~a14668 & a14666;
assign a14672 = ~a14670 & ~a14404;
assign a14674 = ~a14666 & ~a13890;
assign a14676 = ~a14674 & a13350;
assign a14678 = ~a14676 & a14432;
assign a14680 = ~a14676 & a14440;
assign a14682 = ~a14676 & a14444;
assign a14684 = ~a14676 & a14448;
assign a14686 = ~a14684 & ~a14682;
assign a14688 = a14686 & ~a14680;
assign a14690 = a14688 & ~a14678;
assign a14692 = a14690 & ~a14672;
assign a14694 = a14692 & ~a14406;
assign a14696 = a14694 & ~a14420;
assign a14698 = a14696 & ~a14424;
assign a14700 = a14698 & ~a14428;
assign a14702 = ~a14700 & a9332;
assign a14704 = ~a14670 & ~a14482;
assign a14706 = ~a14676 & a14500;
assign a14708 = ~a14676 & a14504;
assign a14710 = ~a14676 & a14508;
assign a14712 = ~a14676 & a14512;
assign a14714 = ~a14712 & ~a14710;
assign a14716 = a14714 & ~a14708;
assign a14718 = a14716 & ~a14706;
assign a14720 = a14718 & ~a14704;
assign a14722 = a14720 & ~a14484;
assign a14724 = a14722 & ~a14488;
assign a14726 = a14724 & ~a14492;
assign a14728 = a14726 & ~a14496;
assign a14730 = ~a14728 & a9572;
assign a14732 = ~a14670 & ~a14546;
assign a14734 = ~a14676 & a14564;
assign a14736 = ~a14676 & a14568;
assign a14738 = ~a14676 & a14572;
assign a14740 = ~a14676 & a14576;
assign a14742 = ~a14740 & ~a14738;
assign a14744 = a14742 & ~a14736;
assign a14746 = a14744 & ~a14734;
assign a14748 = a14746 & ~a14732;
assign a14750 = a14748 & ~a14548;
assign a14752 = a14750 & ~a14552;
assign a14754 = a14752 & ~a14556;
assign a14756 = a14754 & ~a14560;
assign a14758 = ~a14756 & a9812;
assign a14760 = ~a14670 & ~a14610;
assign a14762 = ~a14676 & a14628;
assign a14764 = ~a14676 & a14632;
assign a14766 = ~a14676 & a14636;
assign a14768 = ~a14676 & a14640;
assign a14770 = ~a14768 & ~a14766;
assign a14772 = a14770 & ~a14764;
assign a14774 = a14772 & ~a14762;
assign a14776 = a14774 & ~a14760;
assign a14778 = a14776 & ~a14612;
assign a14780 = a14778 & ~a14616;
assign a14782 = a14780 & ~a14620;
assign a14784 = a14782 & ~a14624;
assign a14786 = ~a14784 & a10052;
assign a14788 = ~a14666 & ~a13622;
assign a14790 = ~a14788 & a14150;
assign a14792 = ~a14790 & ~a14404;
assign a14794 = ~a14412 & ~a14150;
assign a14796 = ~a14794 & a13622;
assign a14798 = ~a14796 & a14406;
assign a14800 = ~a14796 & a14420;
assign a14802 = ~a14796 & a14424;
assign a14804 = ~a14796 & a14428;
assign a14806 = ~a14804 & ~a14802;
assign a14808 = a14806 & ~a14800;
assign a14810 = a14808 & ~a14798;
assign a14812 = a14810 & ~a14792;
assign a14814 = a14812 & ~a14432;
assign a14816 = a14814 & ~a14440;
assign a14818 = a14816 & ~a14444;
assign a14820 = a14818 & ~a14448;
assign a14822 = ~a14820 & a9338;
assign a14824 = ~a14790 & ~a14482;
assign a14826 = ~a14796 & a14484;
assign a14828 = ~a14796 & a14488;
assign a14830 = ~a14796 & a14492;
assign a14832 = ~a14796 & a14496;
assign a14834 = ~a14832 & ~a14830;
assign a14836 = a14834 & ~a14828;
assign a14838 = a14836 & ~a14826;
assign a14840 = a14838 & ~a14824;
assign a14842 = a14840 & ~a14500;
assign a14844 = a14842 & ~a14504;
assign a14846 = a14844 & ~a14508;
assign a14848 = a14846 & ~a14512;
assign a14850 = ~a14848 & a9578;
assign a14852 = ~a14790 & ~a14546;
assign a14854 = ~a14796 & a14548;
assign a14856 = ~a14796 & a14552;
assign a14858 = ~a14796 & a14556;
assign a14860 = ~a14796 & a14560;
assign a14862 = ~a14860 & ~a14858;
assign a14864 = a14862 & ~a14856;
assign a14866 = a14864 & ~a14854;
assign a14868 = a14866 & ~a14852;
assign a14870 = a14868 & ~a14564;
assign a14872 = a14870 & ~a14568;
assign a14874 = a14872 & ~a14572;
assign a14876 = a14874 & ~a14576;
assign a14878 = ~a14876 & a9818;
assign a14880 = ~a14790 & ~a14610;
assign a14882 = ~a14796 & a14612;
assign a14884 = ~a14796 & a14616;
assign a14886 = ~a14796 & a14620;
assign a14888 = ~a14796 & a14624;
assign a14890 = ~a14888 & ~a14886;
assign a14892 = a14890 & ~a14884;
assign a14894 = a14892 & ~a14882;
assign a14896 = a14894 & ~a14880;
assign a14898 = a14896 & ~a14628;
assign a14900 = a14898 & ~a14632;
assign a14902 = a14900 & ~a14636;
assign a14904 = a14902 & ~a14640;
assign a14906 = ~a14904 & a10058;
assign a14908 = ~a7420 & a7418;
assign a14910 = ~a7660 & a7658;
assign a14912 = ~a14910 & ~a14908;
assign a14914 = ~a7900 & a7898;
assign a14916 = ~a14914 & a14912;
assign a14918 = ~a8140 & a8138;
assign a14920 = ~a14918 & a14916;
assign a14922 = ~a8380 & a8378;
assign a14924 = ~a13884 & ~a13616;
assign a14926 = ~a14924 & a14412;
assign a14928 = ~a14926 & a14922;
assign a14930 = ~a8620 & a8618;
assign a14932 = a14930 & ~a14926;
assign a14934 = ~a8860 & a8858;
assign a14936 = a14934 & ~a14926;
assign a14938 = ~a9100 & a9098;
assign a14940 = a14938 & ~a14926;
assign a14942 = ~a9340 & a9338;
assign a14944 = ~a14412 & ~a13344;
assign a14946 = ~a14944 & a13884;
assign a14948 = ~a14946 & a14942;
assign a14950 = ~a9580 & a9578;
assign a14952 = a14950 & ~a14946;
assign a14954 = ~a9820 & a9818;
assign a14956 = a14954 & ~a14946;
assign a14958 = ~a10060 & a10058;
assign a14960 = a14958 & ~a14946;
assign a14962 = ~a14960 & ~a14956;
assign a14964 = a14962 & ~a14952;
assign a14966 = a14964 & ~a14948;
assign a14968 = a14966 & ~a14940;
assign a14970 = a14968 & ~a14936;
assign a14972 = a14970 & ~a14932;
assign a14974 = a14972 & ~a14928;
assign a14976 = a14974 & a14920;
assign a14978 = ~a14976 & a10288;
assign a14980 = ~a7422 & a7418;
assign a14982 = ~a7662 & a7658;
assign a14984 = ~a14982 & ~a14980;
assign a14986 = ~a7902 & a7898;
assign a14988 = ~a14986 & a14984;
assign a14990 = ~a8142 & a8138;
assign a14992 = ~a14990 & a14988;
assign a14994 = ~a8382 & a8378;
assign a14996 = a14994 & ~a14926;
assign a14998 = ~a8622 & a8618;
assign a15000 = a14998 & ~a14926;
assign a15002 = ~a8862 & a8858;
assign a15004 = a15002 & ~a14926;
assign a15006 = ~a9102 & a9098;
assign a15008 = a15006 & ~a14926;
assign a15010 = ~a9342 & a9338;
assign a15012 = a15010 & ~a14946;
assign a15014 = ~a9582 & a9578;
assign a15016 = a15014 & ~a14946;
assign a15018 = ~a9822 & a9818;
assign a15020 = a15018 & ~a14946;
assign a15022 = ~a10062 & a10058;
assign a15024 = a15022 & ~a14946;
assign a15026 = ~a15024 & ~a15020;
assign a15028 = a15026 & ~a15016;
assign a15030 = a15028 & ~a15012;
assign a15032 = a15030 & ~a15008;
assign a15034 = a15032 & ~a15004;
assign a15036 = a15034 & ~a15000;
assign a15038 = a15036 & ~a14996;
assign a15040 = a15038 & a14992;
assign a15042 = ~a15040 & a10528;
assign a15044 = ~a7424 & a7418;
assign a15046 = ~a7664 & a7658;
assign a15048 = ~a15046 & ~a15044;
assign a15050 = ~a7904 & a7898;
assign a15052 = ~a15050 & a15048;
assign a15054 = ~a8144 & a8138;
assign a15056 = ~a15054 & a15052;
assign a15058 = ~a8384 & a8378;
assign a15060 = a15058 & ~a14926;
assign a15062 = ~a8624 & a8618;
assign a15064 = a15062 & ~a14926;
assign a15066 = ~a8864 & a8858;
assign a15068 = a15066 & ~a14926;
assign a15070 = ~a9104 & a9098;
assign a15072 = a15070 & ~a14926;
assign a15074 = ~a9344 & a9338;
assign a15076 = a15074 & ~a14946;
assign a15078 = ~a9584 & a9578;
assign a15080 = a15078 & ~a14946;
assign a15082 = ~a9824 & a9818;
assign a15084 = a15082 & ~a14946;
assign a15086 = ~a10064 & a10058;
assign a15088 = a15086 & ~a14946;
assign a15090 = ~a15088 & ~a15084;
assign a15092 = a15090 & ~a15080;
assign a15094 = a15092 & ~a15076;
assign a15096 = a15094 & ~a15072;
assign a15098 = a15096 & ~a15068;
assign a15100 = a15098 & ~a15064;
assign a15102 = a15100 & ~a15060;
assign a15104 = a15102 & a15056;
assign a15106 = ~a15104 & a10768;
assign a15108 = ~a7426 & a7418;
assign a15110 = ~a7666 & a7658;
assign a15112 = ~a15110 & ~a15108;
assign a15114 = ~a7906 & a7898;
assign a15116 = ~a15114 & a15112;
assign a15118 = ~a8146 & a8138;
assign a15120 = ~a15118 & a15116;
assign a15122 = ~a8386 & a8378;
assign a15124 = a15122 & ~a14926;
assign a15126 = ~a8626 & a8618;
assign a15128 = a15126 & ~a14926;
assign a15130 = ~a8866 & a8858;
assign a15132 = a15130 & ~a14926;
assign a15134 = ~a9106 & a9098;
assign a15136 = a15134 & ~a14926;
assign a15138 = ~a9346 & a9338;
assign a15140 = a15138 & ~a14946;
assign a15142 = ~a9586 & a9578;
assign a15144 = a15142 & ~a14946;
assign a15146 = ~a9826 & a9818;
assign a15148 = a15146 & ~a14946;
assign a15150 = ~a10066 & a10058;
assign a15152 = a15150 & ~a14946;
assign a15154 = ~a15152 & ~a15148;
assign a15156 = a15154 & ~a15144;
assign a15158 = a15156 & ~a15140;
assign a15160 = a15158 & ~a15136;
assign a15162 = a15160 & ~a15132;
assign a15164 = a15162 & ~a15128;
assign a15166 = a15164 & ~a15124;
assign a15168 = a15166 & a15120;
assign a15170 = ~a15168 & a11008;
assign a15172 = ~a14144 & ~a13344;
assign a15174 = ~a15172 & a14666;
assign a15176 = ~a15174 & ~a14920;
assign a15178 = ~a14666 & ~a13884;
assign a15180 = ~a15178 & a13344;
assign a15182 = ~a15180 & a14942;
assign a15184 = ~a15180 & a14950;
assign a15186 = ~a15180 & a14954;
assign a15188 = ~a15180 & a14958;
assign a15190 = ~a15188 & ~a15186;
assign a15192 = a15190 & ~a15184;
assign a15194 = a15192 & ~a15182;
assign a15196 = a15194 & ~a15176;
assign a15198 = a15196 & ~a14922;
assign a15200 = a15198 & ~a14930;
assign a15202 = a15200 & ~a14934;
assign a15204 = a15202 & ~a14938;
assign a15206 = ~a15204 & a10292;
assign a15208 = ~a15174 & ~a14992;
assign a15210 = ~a15180 & a15010;
assign a15212 = ~a15180 & a15014;
assign a15214 = ~a15180 & a15018;
assign a15216 = ~a15180 & a15022;
assign a15218 = ~a15216 & ~a15214;
assign a15220 = a15218 & ~a15212;
assign a15222 = a15220 & ~a15210;
assign a15224 = a15222 & ~a15208;
assign a15226 = a15224 & ~a14994;
assign a15228 = a15226 & ~a14998;
assign a15230 = a15228 & ~a15002;
assign a15232 = a15230 & ~a15006;
assign a15234 = ~a15232 & a10532;
assign a15236 = ~a15174 & ~a15056;
assign a15238 = ~a15180 & a15074;
assign a15240 = ~a15180 & a15078;
assign a15242 = ~a15180 & a15082;
assign a15244 = ~a15180 & a15086;
assign a15246 = ~a15244 & ~a15242;
assign a15248 = a15246 & ~a15240;
assign a15250 = a15248 & ~a15238;
assign a15252 = a15250 & ~a15236;
assign a15254 = a15252 & ~a15058;
assign a15256 = a15254 & ~a15062;
assign a15258 = a15256 & ~a15066;
assign a15260 = a15258 & ~a15070;
assign a15262 = ~a15260 & a10772;
assign a15264 = ~a15174 & ~a15120;
assign a15266 = ~a15180 & a15138;
assign a15268 = ~a15180 & a15142;
assign a15270 = ~a15180 & a15146;
assign a15272 = ~a15180 & a15150;
assign a15274 = ~a15272 & ~a15270;
assign a15276 = a15274 & ~a15268;
assign a15278 = a15276 & ~a15266;
assign a15280 = a15278 & ~a15264;
assign a15282 = a15280 & ~a15122;
assign a15284 = a15282 & ~a15126;
assign a15286 = a15284 & ~a15130;
assign a15288 = a15286 & ~a15134;
assign a15290 = ~a15288 & a11012;
assign a15292 = ~a14666 & ~a13616;
assign a15294 = ~a15292 & a14144;
assign a15296 = ~a15294 & ~a14920;
assign a15298 = ~a14412 & ~a14144;
assign a15300 = ~a15298 & a13616;
assign a15302 = ~a15300 & a14922;
assign a15304 = ~a15300 & a14930;
assign a15306 = ~a15300 & a14934;
assign a15308 = ~a15300 & a14938;
assign a15310 = ~a15308 & ~a15306;
assign a15312 = a15310 & ~a15304;
assign a15314 = a15312 & ~a15302;
assign a15316 = a15314 & ~a15296;
assign a15318 = a15316 & ~a14942;
assign a15320 = a15318 & ~a14950;
assign a15322 = a15320 & ~a14954;
assign a15324 = a15322 & ~a14958;
assign a15326 = ~a15324 & a10296;
assign a15328 = ~a15294 & ~a14992;
assign a15330 = ~a15300 & a14994;
assign a15332 = ~a15300 & a14998;
assign a15334 = ~a15300 & a15002;
assign a15336 = ~a15300 & a15006;
assign a15338 = ~a15336 & ~a15334;
assign a15340 = a15338 & ~a15332;
assign a15342 = a15340 & ~a15330;
assign a15344 = a15342 & ~a15328;
assign a15346 = a15344 & ~a15010;
assign a15348 = a15346 & ~a15014;
assign a15350 = a15348 & ~a15018;
assign a15352 = a15350 & ~a15022;
assign a15354 = ~a15352 & a10536;
assign a15356 = ~a15294 & ~a15056;
assign a15358 = ~a15300 & a15058;
assign a15360 = ~a15300 & a15062;
assign a15362 = ~a15300 & a15066;
assign a15364 = ~a15300 & a15070;
assign a15366 = ~a15364 & ~a15362;
assign a15368 = a15366 & ~a15360;
assign a15370 = a15368 & ~a15358;
assign a15372 = a15370 & ~a15356;
assign a15374 = a15372 & ~a15074;
assign a15376 = a15374 & ~a15078;
assign a15378 = a15376 & ~a15082;
assign a15380 = a15378 & ~a15086;
assign a15382 = ~a15380 & a10776;
assign a15384 = ~a15294 & ~a15120;
assign a15386 = ~a15300 & a15122;
assign a15388 = ~a15300 & a15126;
assign a15390 = ~a15300 & a15130;
assign a15392 = ~a15300 & a15134;
assign a15394 = ~a15392 & ~a15390;
assign a15396 = a15394 & ~a15388;
assign a15398 = a15396 & ~a15386;
assign a15400 = a15398 & ~a15384;
assign a15402 = a15400 & ~a15138;
assign a15404 = a15402 & ~a15142;
assign a15406 = a15404 & ~a15146;
assign a15408 = a15406 & ~a15150;
assign a15410 = ~a15408 & a11016;
assign a15412 = ~a13884 & a13624;
assign a15414 = ~a13890 & a13744;
assign a15416 = ~a15414 & ~a15412;
assign a15418 = a15416 & ~a14924;
assign a15420 = a15418 & ~a14414;
assign a15422 = a15420 & a14412;
assign a15424 = ~a14666 & a13892;
assign a15426 = a14278 & ~a13350;
assign a15428 = ~a15426 & ~a15424;
assign a15430 = a15428 & ~a15178;
assign a15432 = a15430 & ~a13358;
assign a15434 = a15432 & a13344;
assign a15436 = a14434 & ~a14144;
assign a15438 = a14674 & ~a13616;
assign a15440 = ~a15438 & ~a15436;
assign a15442 = a15440 & ~a14158;
assign a15444 = a15442 & ~a13630;
assign a15446 = a15444 & a13382;
assign a15448 = a7404 & l748;
assign a15450 = ~a7404 & ~l748;
assign a15452 = ~a15450 & ~a15448;
assign a15454 = a7644 & l762;
assign a15456 = ~a7644 & ~l762;
assign a15458 = ~a15456 & ~a15454;
assign a15460 = a7884 & l776;
assign a15462 = ~a7884 & ~l776;
assign a15464 = ~a15462 & ~a15460;
assign a15466 = a8124 & l790;
assign a15468 = ~a8124 & ~l790;
assign a15470 = ~a15468 & ~a15466;
assign a15472 = a8364 & l830;
assign a15474 = ~a8364 & ~l830;
assign a15476 = ~a15474 & ~a15472;
assign a15478 = a8604 & l844;
assign a15480 = ~a8604 & ~l844;
assign a15482 = ~a15480 & ~a15478;
assign a15484 = a8844 & l858;
assign a15486 = ~a8844 & ~l858;
assign a15488 = ~a15486 & ~a15484;
assign a15490 = a9084 & l872;
assign a15492 = ~a9084 & ~l872;
assign a15494 = ~a15492 & ~a15490;
assign a15496 = a9324 & l912;
assign a15498 = ~a9324 & ~l912;
assign a15500 = ~a15498 & ~a15496;
assign a15502 = a9564 & l926;
assign a15504 = ~a9564 & ~l926;
assign a15506 = ~a15504 & ~a15502;
assign a15508 = a9804 & l940;
assign a15510 = ~a9804 & ~l940;
assign a15512 = ~a15510 & ~a15508;
assign a15514 = a10044 & l954;
assign a15516 = ~a10044 & ~l954;
assign a15518 = ~a15516 & ~a15514;
assign a15520 = a10284 & l994;
assign a15522 = ~a10284 & ~l994;
assign a15524 = ~a15522 & ~a15520;
assign a15526 = a10524 & l1008;
assign a15528 = ~a10524 & ~l1008;
assign a15530 = ~a15528 & ~a15526;
assign a15532 = a10764 & l1022;
assign a15534 = ~a10764 & ~l1022;
assign a15536 = ~a15534 & ~a15532;
assign a15538 = a11004 & l1036;
assign a15540 = ~a11004 & ~l1036;
assign a15542 = ~a15540 & ~a15538;
assign a15544 = ~l1078 & ~l746;
assign a15546 = l1078 & l746;
assign a15548 = ~a15546 & ~a15544;
assign a15550 = ~l1076 & l744;
assign a15552 = l1076 & ~l744;
assign a15554 = ~a15552 & ~a15550;
assign a15556 = ~l1082 & ~l752;
assign a15558 = l1082 & l752;
assign a15560 = ~a15558 & ~a15556;
assign a15562 = ~l1080 & l750;
assign a15564 = l1080 & ~l750;
assign a15566 = ~a15564 & ~a15562;
assign a15568 = ~l1086 & ~l760;
assign a15570 = l1086 & l760;
assign a15572 = ~a15570 & ~a15568;
assign a15574 = ~l1084 & l758;
assign a15576 = l1084 & ~l758;
assign a15578 = ~a15576 & ~a15574;
assign a15580 = ~l1090 & ~l766;
assign a15582 = l1090 & l766;
assign a15584 = ~a15582 & ~a15580;
assign a15586 = ~l1088 & l764;
assign a15588 = l1088 & ~l764;
assign a15590 = ~a15588 & ~a15586;
assign a15592 = ~l1094 & ~l774;
assign a15594 = l1094 & l774;
assign a15596 = ~a15594 & ~a15592;
assign a15598 = ~l1092 & l772;
assign a15600 = l1092 & ~l772;
assign a15602 = ~a15600 & ~a15598;
assign a15604 = ~l1098 & ~l780;
assign a15606 = l1098 & l780;
assign a15608 = ~a15606 & ~a15604;
assign a15610 = ~l1096 & l778;
assign a15612 = l1096 & ~l778;
assign a15614 = ~a15612 & ~a15610;
assign a15616 = ~l1102 & ~l788;
assign a15618 = l1102 & l788;
assign a15620 = ~a15618 & ~a15616;
assign a15622 = ~l1100 & l786;
assign a15624 = l1100 & ~l786;
assign a15626 = ~a15624 & ~a15622;
assign a15628 = ~l1106 & ~l794;
assign a15630 = l1106 & l794;
assign a15632 = ~a15630 & ~a15628;
assign a15634 = ~l1104 & l792;
assign a15636 = l1104 & ~l792;
assign a15638 = ~a15636 & ~a15634;
assign a15640 = ~l1112 & ~l800;
assign a15642 = l1112 & l800;
assign a15644 = ~a15642 & ~a15640;
assign a15646 = ~l1110 & l798;
assign a15648 = l1110 & ~l798;
assign a15650 = ~a15648 & ~a15646;
assign a15652 = ~l1108 & l796;
assign a15654 = l1108 & ~l796;
assign a15656 = ~a15654 & ~a15652;
assign a15658 = ~l1114 & l802;
assign a15660 = l1114 & ~l802;
assign a15662 = ~a15660 & ~a15658;
assign a15664 = ~l1118 & l806;
assign a15666 = l1118 & ~l806;
assign a15668 = ~a15666 & ~a15664;
assign a15670 = ~l1116 & l804;
assign a15672 = l1116 & ~l804;
assign a15674 = ~a15672 & ~a15670;
assign a15676 = ~l1120 & l810;
assign a15678 = l1120 & ~l810;
assign a15680 = ~a15678 & ~a15676;
assign a15682 = ~l1122 & l812;
assign a15684 = l1122 & ~l812;
assign a15686 = ~a15684 & ~a15682;
assign a15688 = ~l1130 & l820;
assign a15690 = l1130 & ~l820;
assign a15692 = ~a15690 & ~a15688;
assign a15694 = ~l1128 & l818;
assign a15696 = l1128 & ~l818;
assign a15698 = ~a15696 & ~a15694;
assign a15700 = ~l1126 & l816;
assign a15702 = l1126 & ~l816;
assign a15704 = ~a15702 & ~a15700;
assign a15706 = ~l1124 & l814;
assign a15708 = l1124 & ~l814;
assign a15710 = ~a15708 & ~a15706;
assign a15712 = ~l1134 & ~l828;
assign a15714 = l1134 & l828;
assign a15716 = ~a15714 & ~a15712;
assign a15718 = ~l1132 & l826;
assign a15720 = l1132 & ~l826;
assign a15722 = ~a15720 & ~a15718;
assign a15724 = ~l1138 & ~l834;
assign a15726 = l1138 & l834;
assign a15728 = ~a15726 & ~a15724;
assign a15730 = ~l1136 & l832;
assign a15732 = l1136 & ~l832;
assign a15734 = ~a15732 & ~a15730;
assign a15736 = ~l1142 & ~l842;
assign a15738 = l1142 & l842;
assign a15740 = ~a15738 & ~a15736;
assign a15742 = ~l1140 & l840;
assign a15744 = l1140 & ~l840;
assign a15746 = ~a15744 & ~a15742;
assign a15748 = ~l1146 & ~l848;
assign a15750 = l1146 & l848;
assign a15752 = ~a15750 & ~a15748;
assign a15754 = ~l1144 & l846;
assign a15756 = l1144 & ~l846;
assign a15758 = ~a15756 & ~a15754;
assign a15760 = ~l1150 & ~l856;
assign a15762 = l1150 & l856;
assign a15764 = ~a15762 & ~a15760;
assign a15766 = ~l1148 & l854;
assign a15768 = l1148 & ~l854;
assign a15770 = ~a15768 & ~a15766;
assign a15772 = ~l1154 & ~l862;
assign a15774 = l1154 & l862;
assign a15776 = ~a15774 & ~a15772;
assign a15778 = ~l1152 & l860;
assign a15780 = l1152 & ~l860;
assign a15782 = ~a15780 & ~a15778;
assign a15784 = ~l1158 & ~l870;
assign a15786 = l1158 & l870;
assign a15788 = ~a15786 & ~a15784;
assign a15790 = ~l1156 & l868;
assign a15792 = l1156 & ~l868;
assign a15794 = ~a15792 & ~a15790;
assign a15796 = ~l1162 & ~l876;
assign a15798 = l1162 & l876;
assign a15800 = ~a15798 & ~a15796;
assign a15802 = ~l1160 & l874;
assign a15804 = l1160 & ~l874;
assign a15806 = ~a15804 & ~a15802;
assign a15808 = ~l1168 & ~l882;
assign a15810 = l1168 & l882;
assign a15812 = ~a15810 & ~a15808;
assign a15814 = ~l1166 & l880;
assign a15816 = l1166 & ~l880;
assign a15818 = ~a15816 & ~a15814;
assign a15820 = ~l1164 & l878;
assign a15822 = l1164 & ~l878;
assign a15824 = ~a15822 & ~a15820;
assign a15826 = ~l1170 & l884;
assign a15828 = l1170 & ~l884;
assign a15830 = ~a15828 & ~a15826;
assign a15832 = ~l1174 & l888;
assign a15834 = l1174 & ~l888;
assign a15836 = ~a15834 & ~a15832;
assign a15838 = ~l1172 & l886;
assign a15840 = l1172 & ~l886;
assign a15842 = ~a15840 & ~a15838;
assign a15844 = ~l1176 & l892;
assign a15846 = l1176 & ~l892;
assign a15848 = ~a15846 & ~a15844;
assign a15850 = ~l1178 & l894;
assign a15852 = l1178 & ~l894;
assign a15854 = ~a15852 & ~a15850;
assign a15856 = ~l1186 & l902;
assign a15858 = l1186 & ~l902;
assign a15860 = ~a15858 & ~a15856;
assign a15862 = ~l1184 & l900;
assign a15864 = l1184 & ~l900;
assign a15866 = ~a15864 & ~a15862;
assign a15868 = ~l1182 & l898;
assign a15870 = l1182 & ~l898;
assign a15872 = ~a15870 & ~a15868;
assign a15874 = ~l1180 & l896;
assign a15876 = l1180 & ~l896;
assign a15878 = ~a15876 & ~a15874;
assign a15880 = ~l1190 & ~l910;
assign a15882 = l1190 & l910;
assign a15884 = ~a15882 & ~a15880;
assign a15886 = ~l1188 & l908;
assign a15888 = l1188 & ~l908;
assign a15890 = ~a15888 & ~a15886;
assign a15892 = ~l1194 & ~l916;
assign a15894 = l1194 & l916;
assign a15896 = ~a15894 & ~a15892;
assign a15898 = ~l1192 & l914;
assign a15900 = l1192 & ~l914;
assign a15902 = ~a15900 & ~a15898;
assign a15904 = ~l1198 & ~l924;
assign a15906 = l1198 & l924;
assign a15908 = ~a15906 & ~a15904;
assign a15910 = ~l1196 & l922;
assign a15912 = l1196 & ~l922;
assign a15914 = ~a15912 & ~a15910;
assign a15916 = ~l1202 & ~l930;
assign a15918 = l1202 & l930;
assign a15920 = ~a15918 & ~a15916;
assign a15922 = ~l1200 & l928;
assign a15924 = l1200 & ~l928;
assign a15926 = ~a15924 & ~a15922;
assign a15928 = ~l1206 & ~l938;
assign a15930 = l1206 & l938;
assign a15932 = ~a15930 & ~a15928;
assign a15934 = ~l1204 & l936;
assign a15936 = l1204 & ~l936;
assign a15938 = ~a15936 & ~a15934;
assign a15940 = ~l1210 & ~l944;
assign a15942 = l1210 & l944;
assign a15944 = ~a15942 & ~a15940;
assign a15946 = ~l1208 & l942;
assign a15948 = l1208 & ~l942;
assign a15950 = ~a15948 & ~a15946;
assign a15952 = ~l1214 & ~l952;
assign a15954 = l1214 & l952;
assign a15956 = ~a15954 & ~a15952;
assign a15958 = ~l1212 & l950;
assign a15960 = l1212 & ~l950;
assign a15962 = ~a15960 & ~a15958;
assign a15964 = ~l1218 & ~l958;
assign a15966 = l1218 & l958;
assign a15968 = ~a15966 & ~a15964;
assign a15970 = ~l1216 & l956;
assign a15972 = l1216 & ~l956;
assign a15974 = ~a15972 & ~a15970;
assign a15976 = ~l1224 & ~l964;
assign a15978 = l1224 & l964;
assign a15980 = ~a15978 & ~a15976;
assign a15982 = ~l1222 & l962;
assign a15984 = l1222 & ~l962;
assign a15986 = ~a15984 & ~a15982;
assign a15988 = ~l1220 & l960;
assign a15990 = l1220 & ~l960;
assign a15992 = ~a15990 & ~a15988;
assign a15994 = ~l1226 & l966;
assign a15996 = l1226 & ~l966;
assign a15998 = ~a15996 & ~a15994;
assign a16000 = ~l1230 & l970;
assign a16002 = l1230 & ~l970;
assign a16004 = ~a16002 & ~a16000;
assign a16006 = ~l1228 & l968;
assign a16008 = l1228 & ~l968;
assign a16010 = ~a16008 & ~a16006;
assign a16012 = ~l1232 & l974;
assign a16014 = l1232 & ~l974;
assign a16016 = ~a16014 & ~a16012;
assign a16018 = ~l1234 & l976;
assign a16020 = l1234 & ~l976;
assign a16022 = ~a16020 & ~a16018;
assign a16024 = ~l1242 & l984;
assign a16026 = l1242 & ~l984;
assign a16028 = ~a16026 & ~a16024;
assign a16030 = ~l1240 & l982;
assign a16032 = l1240 & ~l982;
assign a16034 = ~a16032 & ~a16030;
assign a16036 = ~l1238 & l980;
assign a16038 = l1238 & ~l980;
assign a16040 = ~a16038 & ~a16036;
assign a16042 = ~l1236 & l978;
assign a16044 = l1236 & ~l978;
assign a16046 = ~a16044 & ~a16042;
assign a16048 = ~l1246 & ~l992;
assign a16050 = l1246 & l992;
assign a16052 = ~a16050 & ~a16048;
assign a16054 = ~l1244 & l990;
assign a16056 = l1244 & ~l990;
assign a16058 = ~a16056 & ~a16054;
assign a16060 = ~l1250 & ~l998;
assign a16062 = l1250 & l998;
assign a16064 = ~a16062 & ~a16060;
assign a16066 = ~l1248 & l996;
assign a16068 = l1248 & ~l996;
assign a16070 = ~a16068 & ~a16066;
assign a16072 = ~l1254 & ~l1006;
assign a16074 = l1254 & l1006;
assign a16076 = ~a16074 & ~a16072;
assign a16078 = ~l1252 & l1004;
assign a16080 = l1252 & ~l1004;
assign a16082 = ~a16080 & ~a16078;
assign a16084 = ~l1258 & ~l1012;
assign a16086 = l1258 & l1012;
assign a16088 = ~a16086 & ~a16084;
assign a16090 = ~l1256 & l1010;
assign a16092 = l1256 & ~l1010;
assign a16094 = ~a16092 & ~a16090;
assign a16096 = ~l1262 & ~l1020;
assign a16098 = l1262 & l1020;
assign a16100 = ~a16098 & ~a16096;
assign a16102 = ~l1260 & l1018;
assign a16104 = l1260 & ~l1018;
assign a16106 = ~a16104 & ~a16102;
assign a16108 = ~l1266 & ~l1026;
assign a16110 = l1266 & l1026;
assign a16112 = ~a16110 & ~a16108;
assign a16114 = ~l1264 & l1024;
assign a16116 = l1264 & ~l1024;
assign a16118 = ~a16116 & ~a16114;
assign a16120 = ~l1270 & ~l1034;
assign a16122 = l1270 & l1034;
assign a16124 = ~a16122 & ~a16120;
assign a16126 = ~l1268 & l1032;
assign a16128 = l1268 & ~l1032;
assign a16130 = ~a16128 & ~a16126;
assign a16132 = ~l1274 & ~l1040;
assign a16134 = l1274 & l1040;
assign a16136 = ~a16134 & ~a16132;
assign a16138 = ~l1272 & l1038;
assign a16140 = l1272 & ~l1038;
assign a16142 = ~a16140 & ~a16138;
assign a16144 = ~l1278 & l1044;
assign a16146 = l1278 & ~l1044;
assign a16148 = ~a16146 & ~a16144;
assign a16150 = ~l1276 & l1042;
assign a16152 = l1276 & ~l1042;
assign a16154 = ~a16152 & ~a16150;
assign a16156 = ~l1282 & l1048;
assign a16158 = l1282 & ~l1048;
assign a16160 = ~a16158 & ~a16156;
assign a16162 = ~l1286 & l1052;
assign a16164 = l1286 & ~l1052;
assign a16166 = ~a16164 & ~a16162;
assign a16168 = ~l1284 & l1050;
assign a16170 = l1284 & ~l1050;
assign a16172 = ~a16170 & ~a16168;
assign a16174 = ~l1288 & l1056;
assign a16176 = l1288 & ~l1056;
assign a16178 = ~a16176 & ~a16174;
assign a16180 = ~l1290 & l1058;
assign a16182 = l1290 & ~l1058;
assign a16184 = ~a16182 & ~a16180;
assign a16186 = ~l1298 & l1066;
assign a16188 = l1298 & ~l1066;
assign a16190 = ~a16188 & ~a16186;
assign a16192 = ~l1296 & l1064;
assign a16194 = l1296 & ~l1064;
assign a16196 = ~a16194 & ~a16192;
assign a16198 = ~l1294 & l1062;
assign a16200 = l1294 & ~l1062;
assign a16202 = ~a16200 & ~a16198;
assign a16204 = ~l1292 & l1060;
assign a16206 = l1292 & ~l1060;
assign a16208 = ~a16206 & ~a16204;
assign a16210 = ~l1300 & l1068;
assign a16212 = l1300 & ~l1068;
assign a16214 = ~a16212 & ~a16210;
assign a16216 = l1302 & ~l1070;
assign a16218 = ~l1302 & l1070;
assign a16220 = ~a16218 & ~a16216;
assign a16222 = l1304 & ~l1072;
assign a16224 = ~l1304 & l1072;
assign a16226 = ~a16224 & ~a16222;
assign a16228 = l1306 & ~l1074;
assign a16230 = ~l1306 & l1074;
assign a16232 = ~a16230 & ~a16228;
assign a16234 = a16232 & a16226;
assign a16236 = a16234 & a16220;
assign a16238 = a16236 & a16214;
assign a16240 = a16238 & a16208;
assign a16242 = a16240 & a16202;
assign a16244 = a16242 & a16196;
assign a16246 = a16244 & a16190;
assign a16248 = a16246 & a16184;
assign a16250 = a16248 & a16178;
assign a16252 = a16250 & a16172;
assign a16254 = a16252 & a16166;
assign a16256 = a16254 & a16160;
assign a16258 = a16256 & a16154;
assign a16260 = a16258 & a16148;
assign a16262 = ~l1280 & ~l1046;
assign a16264 = l1280 & l1046;
assign a16266 = ~a16264 & ~a16262;
assign a16268 = a16266 & a16260;
assign a16270 = a16268 & a16142;
assign a16272 = a16270 & a16136;
assign a16274 = a16272 & a16130;
assign a16276 = a16274 & a16124;
assign a16278 = a16276 & a16118;
assign a16280 = a16278 & a16112;
assign a16282 = a16280 & a16106;
assign a16284 = a16282 & a16100;
assign a16286 = a16284 & a16094;
assign a16288 = a16286 & a16088;
assign a16290 = a16288 & a16082;
assign a16292 = a16290 & a16076;
assign a16294 = a16292 & a16070;
assign a16296 = a16294 & a16064;
assign a16298 = a16296 & a16058;
assign a16300 = a16298 & a16052;
assign a16302 = a16300 & a16046;
assign a16304 = a16302 & a16040;
assign a16306 = a16304 & a16034;
assign a16308 = a16306 & a16028;
assign a16310 = a16308 & a16022;
assign a16312 = a16310 & a16016;
assign a16314 = a16312 & a16010;
assign a16316 = a16314 & a16004;
assign a16318 = a16316 & a15998;
assign a16320 = a16318 & a15992;
assign a16322 = a16320 & a15986;
assign a16324 = a16322 & a15980;
assign a16326 = a16324 & a15974;
assign a16328 = a16326 & a15968;
assign a16330 = a16328 & a15962;
assign a16332 = a16330 & a15956;
assign a16334 = a16332 & a15950;
assign a16336 = a16334 & a15944;
assign a16338 = a16336 & a15938;
assign a16340 = a16338 & a15932;
assign a16342 = a16340 & a15926;
assign a16344 = a16342 & a15920;
assign a16346 = a16344 & a15914;
assign a16348 = a16346 & a15908;
assign a16350 = a16348 & a15902;
assign a16352 = a16350 & a15896;
assign a16354 = a16352 & a15890;
assign a16356 = a16354 & a15884;
assign a16358 = a16356 & a15878;
assign a16360 = a16358 & a15872;
assign a16362 = a16360 & a15866;
assign a16364 = a16362 & a15860;
assign a16366 = a16364 & a15854;
assign a16368 = a16366 & a15848;
assign a16370 = a16368 & a15842;
assign a16372 = a16370 & a15836;
assign a16374 = a16372 & a15830;
assign a16376 = a16374 & a15824;
assign a16378 = a16376 & a15818;
assign a16380 = a16378 & a15812;
assign a16382 = a16380 & a15806;
assign a16384 = a16382 & a15800;
assign a16386 = a16384 & a15794;
assign a16388 = a16386 & a15788;
assign a16390 = a16388 & a15782;
assign a16392 = a16390 & a15776;
assign a16394 = a16392 & a15770;
assign a16396 = a16394 & a15764;
assign a16398 = a16396 & a15758;
assign a16400 = a16398 & a15752;
assign a16402 = a16400 & a15746;
assign a16404 = a16402 & a15740;
assign a16406 = a16404 & a15734;
assign a16408 = a16406 & a15728;
assign a16410 = a16408 & a15722;
assign a16412 = a16410 & a15716;
assign a16414 = a16412 & a15710;
assign a16416 = a16414 & a15704;
assign a16418 = a16416 & a15698;
assign a16420 = a16418 & a15692;
assign a16422 = a16420 & a15686;
assign a16424 = a16422 & a15680;
assign a16426 = a16424 & a15674;
assign a16428 = a16426 & a15668;
assign a16430 = a16428 & a15662;
assign a16432 = a16430 & a15656;
assign a16434 = a16432 & a15650;
assign a16436 = a16434 & a15644;
assign a16438 = a16436 & a15638;
assign a16440 = a16438 & a15632;
assign a16442 = a16440 & a15626;
assign a16444 = a16442 & a15620;
assign a16446 = a16444 & a15614;
assign a16448 = a16446 & a15608;
assign a16450 = a16448 & a15602;
assign a16452 = a16450 & a15596;
assign a16454 = a16452 & a15590;
assign a16456 = a16454 & a15584;
assign a16458 = a16456 & a15578;
assign a16460 = a16458 & a15572;
assign a16462 = a16460 & a15566;
assign a16464 = a16462 & a15560;
assign a16466 = a16464 & a15554;
assign a16468 = a16466 & a15548;
assign a16470 = a16468 & l1316;
assign a16472 = a16470 & l1308;
assign a16474 = a16472 & l1310;
assign a16476 = a16474 & l1312;
assign a16478 = ~a16476 & i570;
assign a16480 = ~a16478 & a15542;
assign a16482 = a16480 & a15536;
assign a16484 = a16482 & a15530;
assign a16486 = a16484 & a15524;
assign a16488 = a16486 & a15518;
assign a16490 = a16488 & a15512;
assign a16492 = a16490 & a15506;
assign a16494 = a16492 & a15500;
assign a16496 = a16494 & a15494;
assign a16498 = a16496 & a15488;
assign a16500 = a16498 & a15482;
assign a16502 = a16500 & a15476;
assign a16504 = a16502 & a15470;
assign a16506 = a16504 & a15464;
assign a16508 = a16506 & a15458;
assign a16510 = a16508 & a15452;
assign a16512 = a16510 & ~a15446;
assign a16514 = a16512 & ~a15434;
assign a16516 = a16514 & ~a15422;
assign a16518 = a16516 & ~a15410;
assign a16520 = a16518 & ~a15382;
assign a16522 = a16520 & ~a15354;
assign a16524 = a16522 & ~a15326;
assign a16526 = a16524 & ~a15290;
assign a16528 = a16526 & ~a15262;
assign a16530 = a16528 & ~a15234;
assign a16532 = a16530 & ~a15206;
assign a16534 = a16532 & ~a15170;
assign a16536 = a16534 & ~a15106;
assign a16538 = a16536 & ~a15042;
assign a16540 = a16538 & ~a14978;
assign a16542 = a16540 & ~a14906;
assign a16544 = a16542 & ~a14878;
assign a16546 = a16544 & ~a14850;
assign a16548 = a16546 & ~a14822;
assign a16550 = a16548 & ~a14786;
assign a16552 = a16550 & ~a14758;
assign a16554 = a16552 & ~a14730;
assign a16556 = a16554 & ~a14702;
assign a16558 = a16556 & ~a14660;
assign a16560 = a16558 & ~a14596;
assign a16562 = a16560 & ~a14532;
assign a16564 = a16562 & ~a14468;
assign a16566 = a16564 & ~a14390;
assign a16568 = a16566 & ~a14362;
assign a16570 = a16568 & ~a14334;
assign a16572 = a16570 & ~a14306;
assign a16574 = a16572 & ~a14270;
assign a16576 = a16574 & ~a14242;
assign a16578 = a16576 & ~a14214;
assign a16580 = a16578 & ~a14186;
assign a16582 = a16580 & ~a14138;
assign a16584 = a16582 & ~a14074;
assign a16586 = a16584 & ~a14010;
assign a16588 = a16586 & ~a13946;
assign a16590 = a16588 & ~a13862;
assign a16592 = a16590 & ~a13834;
assign a16594 = a16592 & ~a13806;
assign a16596 = a16594 & ~a13778;
assign a16598 = a16596 & ~a13742;
assign a16600 = a16598 & ~a13714;
assign a16602 = a16600 & ~a13686;
assign a16604 = a16602 & ~a13658;
assign a16606 = a16604 & ~a13610;
assign a16608 = a16606 & ~a13546;
assign a16610 = a16608 & ~a13482;
assign a16612 = a16610 & ~a13418;
assign a16614 = a16612 & a13322;
assign a16616 = a16614 & ~a11018;
assign a16618 = a16616 & a13192;
assign a16620 = a16618 & ~a10778;
assign a16622 = a16620 & a13062;
assign a16624 = a16622 & ~a10538;
assign a16626 = a16624 & a12932;
assign a16628 = a16626 & ~a10298;
assign a16630 = a16628 & a12802;
assign a16632 = a16630 & ~a10056;
assign a16634 = a16632 & a12672;
assign a16636 = a16634 & ~a9816;
assign a16638 = a16636 & a12542;
assign a16640 = a16638 & ~a9576;
assign a16642 = a16640 & a12412;
assign a16644 = a16642 & ~a9336;
assign a16646 = a16644 & a12282;
assign a16648 = a16646 & ~a9092;
assign a16650 = a16648 & a12152;
assign a16652 = a16650 & ~a8852;
assign a16654 = a16652 & a12022;
assign a16656 = a16654 & ~a8612;
assign a16658 = a16656 & a11892;
assign a16660 = a16658 & ~a8372;
assign a16662 = a16660 & a11762;
assign a16664 = a16662 & ~a8128;
assign a16666 = a16664 & a11632;
assign a16668 = a16666 & ~a7888;
assign a16670 = a16668 & a11502;
assign a16672 = a16670 & ~a7648;
assign a16674 = a16672 & a11372;
assign a16676 = a16674 & ~a7408;
assign a16678 = a16676 & ~a11242;
assign a16680 = a16678 & ~a11002;
assign a16682 = a16680 & ~a10762;
assign a16684 = a16682 & ~a10522;
assign a16686 = a16684 & ~a10282;
assign a16688 = a16686 & ~a10042;
assign a16690 = a16688 & ~a9802;
assign a16692 = a16690 & ~a9562;
assign a16694 = a16692 & ~a9322;
assign a16696 = a16694 & ~a9082;
assign a16698 = a16696 & ~a8842;
assign a16700 = a16698 & ~a8602;
assign a16702 = a16700 & ~a8362;
assign a16704 = a16702 & ~a8122;
assign a16706 = a16704 & ~a7882;
assign a16708 = a16706 & ~a7642;
assign a16710 = a16708 & ~a7402;
assign a16712 = a16710 & ~a7334;
assign a16714 = a16712 & ~a7330;
assign a16716 = a16714 & ~a7326;
assign a16718 = a16716 & ~a7324;
assign a16720 = a16718 & ~a7322;
assign a16722 = a16720 & ~a7320;
assign a16724 = a16722 & ~a7318;
assign a16726 = a16724 & ~a7314;
assign a16728 = a16726 & ~a7310;
assign a16730 = a16728 & ~a7308;
assign a16732 = a16730 & ~a7306;
assign a16734 = a16732 & ~a7304;
assign a16736 = a16734 & ~a7302;
assign a16738 = a16736 & ~a7298;
assign a16740 = a16738 & ~a7294;
assign a16742 = a16740 & ~a7292;
assign a16744 = a16742 & ~a7290;
assign a16746 = a16744 & ~a7288;
assign a16748 = a16746 & ~a7286;
assign a16750 = a16748 & ~a7282;
assign a16752 = a16750 & ~a7278;
assign a16754 = a16752 & ~a7276;
assign a16756 = a16754 & ~a7274;
assign a16758 = a16756 & ~a7272;
assign a16760 = a16758 & ~a7270;
assign a16762 = a16760 & ~a7268;
assign a16764 = a16762 & ~a7266;
assign a16766 = a16764 & ~a7264;
assign a16768 = a16766 & ~a7262;
assign a16770 = a16768 & ~a7260;
assign a16772 = a16770 & ~a7258;
assign a16774 = a16772 & ~a7256;
assign a16776 = a16774 & ~a7254;
assign a16778 = a16776 & ~a7252;
assign a16780 = a16778 & ~a7250;
assign a16782 = a16780 & ~a7248;
assign a16784 = a16782 & ~a7246;
assign a16786 = a16784 & ~a7244;
assign a16788 = a16786 & ~a7242;
assign a16790 = a16788 & ~a7240;
assign a16792 = a16790 & ~a7238;
assign a16794 = a16792 & ~a7236;
assign a16796 = a16794 & ~a7234;
assign a16798 = a16796 & ~a7232;
assign a16800 = a16798 & ~a7230;
assign a16802 = a16800 & ~a7228;
assign a16804 = a16802 & ~a7226;
assign a16806 = a16804 & ~a7224;
assign a16808 = a16806 & ~a7222;
assign a16810 = a16808 & ~a7220;
assign a16812 = a16810 & ~a7218;
assign a16814 = a16812 & ~a7216;
assign a16816 = a16814 & ~a7214;
assign a16818 = a16816 & ~a7212;
assign a16820 = a16818 & ~a7210;
assign a16822 = a16820 & ~a7208;
assign a16824 = a16822 & ~a7206;
assign a16826 = a16824 & ~a7204;
assign a16828 = a16826 & ~a7202;
assign a16830 = a16828 & ~a7200;
assign a16832 = a16830 & ~a7198;
assign a16834 = a16832 & ~a7196;
assign a16836 = a16834 & ~a7194;
assign a16838 = a16836 & ~a7192;
assign a16840 = a16838 & ~a7190;
assign a16842 = a16840 & ~a7186;
assign a16844 = a16842 & ~a7182;
assign a16846 = a16844 & ~a7178;
assign a16848 = a16846 & ~a7174;
assign a16850 = a16848 & ~a7170;
assign a16852 = a16850 & ~a7166;
assign a16854 = a16852 & ~a7162;
assign a16856 = a16854 & ~a7158;
assign a16858 = a16856 & ~a7154;
assign a16860 = a16858 & ~a7150;
assign a16862 = a16860 & ~a7146;
assign a16864 = a16862 & ~a7142;
assign a16866 = a16864 & ~a7138;
assign a16868 = a16866 & ~a7134;
assign a16870 = a16868 & ~a7130;
assign a16872 = a16870 & l1326;
assign a16874 = a16872 & a7126;
assign a16878 = a16872 & i570;
assign p0 = a16878;

assert property (~p0);

endmodule
