module m139454p (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474,i476,i478,i480,
i482,i484,i486,i488,i490,i492,i494,i496,i498,i500,i502,i504,i506,i508,i510,
i512,i514,i516,i518,i520,i522,i524,i526,i528,i530,i532,i534,i536,i538,i540,
i542,i544,i546,i548,i550,i552,i554,i556,i558,i560,i562,i564,i566,i568,i570,
i572,i574,i576,i578,i580,i582,i584,i586,i588,i590,i592,i594,i596,i598,i600,
i602,i604,i606,i608,i610,i612,i614,i616,i618,i620,i622,i624,i626,i628,i630,
i632,i634,i636,i638,i640,i642,i644,i646,i648,i650,i652,i654,i656,i658,i660,
i662,i664,i666,i668,i670,i672,i674,i676,i678,i680,i682,i684,i686,i688,i690,
i692,i694,i696,i698,i700,i702,i704,i706,i708,i710,i712,i714,i716,i718,i720,
i722,i724,i726,i728,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474,i476,i478,i480,
i482,i484,i486,i488,i490,i492,i494,i496,i498,i500,i502,i504,i506,i508,i510,
i512,i514,i516,i518,i520,i522,i524,i526,i528,i530,i532,i534,i536,i538,i540,
i542,i544,i546,i548,i550,i552,i554,i556,i558,i560,i562,i564,i566,i568,i570,
i572,i574,i576,i578,i580,i582,i584,i586,i588,i590,i592,i594,i596,i598,i600,
i602,i604,i606,i608,i610,i612,i614,i616,i618,i620,i622,i624,i626,i628,i630,
i632,i634,i636,i638,i640,i642,i644,i646,i648,i650,i652,i654,i656,i658,i660,
i662,i664,i666,i668,i670,i672,i674,i676,i678,i680,i682,i684,i686,i688,i690,
i692,i694,i696,i698,i700,i702,i704,i706,i708,i710,i712,i714,i716,i718,i720,
i722,i724,i726,i728;

output p0;

wire a1736,a1752,a1780,a1824,a1840,a1860,a1904,a1920,a1940,a1984,a2000,a2020,a2136,a2160,a2188,
a2200,a2526,a2536,a2546,a2556,a2564,a2622,a2638,a2666,a2710,a2726,a2746,a2790,a2806,a2826,
a2870,a2886,a2906,a3022,a3046,a3074,a3086,a3412,a3422,a3432,a3442,a3450,a3508,a3524,a3552,
a3596,a3612,a3632,a3676,a3692,a3712,a3756,a3772,a3792,a3908,a3932,a3960,a3972,a4298,a4308,
a4318,a4328,a4336,a4394,a4410,a4438,a4482,a4498,a4518,a4562,a4578,a4598,a4642,a4658,a4678,
a4794,a4818,a4846,a4858,a5184,a5194,a5204,a5214,a5222,a5280,a5296,a5324,a5368,a5384,a5404,
a5448,a5464,a5484,a5528,a5544,a5564,a5680,a5704,a5732,a5744,a6070,a6080,a6090,a6100,a6108,
a6114,a6122,a6132,a6140,a6142,a26802,c1,a1680,a1682,a1684,a1686,a1688,a1690,a1692,a1694,
a1696,a1698,a1700,a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,
a1726,a1728,a1730,a1732,a1734,a1738,a1740,a1742,a1744,a1746,a1748,a1750,a1754,a1756,a1758,
a1760,a1762,a1764,a1766,a1768,a1770,a1772,a1774,a1776,a1778,a1782,a1784,a1786,a1788,a1790,
a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,
a1822,a1826,a1828,a1830,a1832,a1834,a1836,a1838,a1842,a1844,a1846,a1848,a1850,a1852,a1854,
a1856,a1858,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,a1882,a1884,a1886,
a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1906,a1908,a1910,a1912,a1914,a1916,a1918,
a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,a1938,a1942,a1944,a1946,a1948,a1950,a1952,
a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,a1972,a1974,a1976,a1978,a1980,a1982,
a1986,a1988,a1990,a1992,a1994,a1996,a1998,a2002,a2004,a2006,a2008,a2010,a2012,a2014,a2016,
a2018,a2022,a2024,a2026,a2028,a2030,a2032,a2034,a2036,a2038,a2040,a2042,a2044,a2046,a2048,
a2050,a2052,a2054,a2056,a2058,a2060,a2062,a2064,a2066,a2068,a2070,a2072,a2074,a2076,a2078,
a2080,a2082,a2084,a2086,a2088,a2090,a2092,a2094,a2096,a2098,a2100,a2102,a2104,a2106,a2108,
a2110,a2112,a2114,a2116,a2118,a2120,a2122,a2124,a2126,a2128,a2130,a2132,a2134,a2138,a2140,
a2142,a2144,a2146,a2148,a2150,a2152,a2154,a2156,a2158,a2162,a2164,a2166,a2168,a2170,a2172,
a2174,a2176,a2178,a2180,a2182,a2184,a2186,a2190,a2192,a2194,a2196,a2198,a2202,a2204,a2206,
a2208,a2210,a2212,a2214,a2216,a2218,a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,
a2238,a2240,a2242,a2244,a2246,a2248,a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,
a2268,a2270,a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,
a2298,a2300,a2302,a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,
a2328,a2330,a2332,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,
a2358,a2360,a2362,a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,
a2388,a2390,a2392,a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,
a2418,a2420,a2422,a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,
a2448,a2450,a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,
a2478,a2480,a2482,a2484,a2486,a2488,a2490,a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,
a2508,a2510,a2512,a2514,a2516,a2518,a2520,a2522,a2524,a2528,a2530,a2532,a2534,a2538,a2540,
a2542,a2544,a2548,a2550,a2552,a2554,a2558,a2560,a2562,a2566,a2568,a2570,a2572,a2574,a2576,
a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,a2602,a2604,a2606,
a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2624,a2626,a2628,a2630,a2632,a2634,a2636,a2640,
a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,a2662,a2664,a2668,a2670,a2672,
a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,a2692,a2694,a2696,a2698,a2700,a2702,
a2704,a2706,a2708,a2712,a2714,a2716,a2718,a2720,a2722,a2724,a2728,a2730,a2732,a2734,a2736,
a2738,a2740,a2742,a2744,a2748,a2750,a2752,a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,
a2770,a2772,a2774,a2776,a2778,a2780,a2782,a2784,a2786,a2788,a2792,a2794,a2796,a2798,a2800,
a2802,a2804,a2808,a2810,a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2828,a2830,a2832,a2834,
a2836,a2838,a2840,a2842,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,
a2866,a2868,a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2888,a2890,a2892,a2894,a2896,a2898,
a2900,a2902,a2904,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2930,
a2932,a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,a2960,
a2962,a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,a2988,a2990,
a2992,a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,
a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3048,a3050,a3052,a3054,
a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3076,a3078,a3080,a3082,a3084,a3088,
a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,a3112,a3114,a3116,a3118,
a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,a3142,a3144,a3146,a3148,
a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,a3172,a3174,a3176,a3178,
a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3200,a3202,a3204,a3206,a3208,
a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,a3228,a3230,a3232,a3234,a3236,a3238,
a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,a3262,a3264,a3266,a3268,
a3270,a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,a3288,a3290,a3292,a3294,a3296,a3298,
a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,a3324,a3326,a3328,
a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,a3354,a3356,a3358,
a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3382,a3384,a3386,a3388,
a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,a3408,a3410,a3414,a3416,a3418,a3420,
a3424,a3426,a3428,a3430,a3434,a3436,a3438,a3440,a3444,a3446,a3448,a3452,a3454,a3456,a3458,
a3460,a3462,a3464,a3466,a3468,a3470,a3472,a3474,a3476,a3478,a3480,a3482,a3484,a3486,a3488,
a3490,a3492,a3494,a3496,a3498,a3500,a3502,a3504,a3506,a3510,a3512,a3514,a3516,a3518,a3520,
a3522,a3526,a3528,a3530,a3532,a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3554,
a3556,a3558,a3560,a3562,a3564,a3566,a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,
a3586,a3588,a3590,a3592,a3594,a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3614,a3616,a3618,
a3620,a3622,a3624,a3626,a3628,a3630,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3648,a3650,
a3652,a3654,a3656,a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3678,a3680,a3682,
a3684,a3686,a3688,a3690,a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,a3714,a3716,
a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,a3738,a3740,a3742,a3744,a3746,
a3748,a3750,a3752,a3754,a3758,a3760,a3762,a3764,a3766,a3768,a3770,a3774,a3776,a3778,a3780,
a3782,a3784,a3786,a3788,a3790,a3794,a3796,a3798,a3800,a3802,a3804,a3806,a3808,a3810,a3812,
a3814,a3816,a3818,a3820,a3822,a3824,a3826,a3828,a3830,a3832,a3834,a3836,a3838,a3840,a3842,
a3844,a3846,a3848,a3850,a3852,a3854,a3856,a3858,a3860,a3862,a3864,a3866,a3868,a3870,a3872,
a3874,a3876,a3878,a3880,a3882,a3884,a3886,a3888,a3890,a3892,a3894,a3896,a3898,a3900,a3902,
a3904,a3906,a3910,a3912,a3914,a3916,a3918,a3920,a3922,a3924,a3926,a3928,a3930,a3934,a3936,
a3938,a3940,a3942,a3944,a3946,a3948,a3950,a3952,a3954,a3956,a3958,a3962,a3964,a3966,a3968,
a3970,a3974,a3976,a3978,a3980,a3982,a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,
a4002,a4004,a4006,a4008,a4010,a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,
a4032,a4034,a4036,a4038,a4040,a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,
a4062,a4064,a4066,a4068,a4070,a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,
a4092,a4094,a4096,a4098,a4100,a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,
a4122,a4124,a4126,a4128,a4130,a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,
a4152,a4154,a4156,a4158,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,
a4182,a4184,a4186,a4188,a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,
a4212,a4214,a4216,a4218,a4220,a4222,a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,
a4242,a4244,a4246,a4248,a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,
a4272,a4274,a4276,a4278,a4280,a4282,a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4300,a4302,
a4304,a4306,a4310,a4312,a4314,a4316,a4320,a4322,a4324,a4326,a4330,a4332,a4334,a4338,a4340,
a4342,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,a4368,a4370,
a4372,a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,a4396,a4398,a4400,a4402,
a4404,a4406,a4408,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,a4432,a4434,
a4436,a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,a4458,a4460,a4462,a4464,a4466,
a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4484,a4486,a4488,a4490,a4492,a4494,a4496,a4500,
a4502,a4504,a4506,a4508,a4510,a4512,a4514,a4516,a4520,a4522,a4524,a4526,a4528,a4530,a4532,
a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,a4554,a4556,a4558,a4560,a4564,
a4566,a4568,a4570,a4572,a4574,a4576,a4580,a4582,a4584,a4586,a4588,a4590,a4592,a4594,a4596,
a4600,a4602,a4604,a4606,a4608,a4610,a4612,a4614,a4616,a4618,a4620,a4622,a4624,a4626,a4628,
a4630,a4632,a4634,a4636,a4638,a4640,a4644,a4646,a4648,a4650,a4652,a4654,a4656,a4660,a4662,
a4664,a4666,a4668,a4670,a4672,a4674,a4676,a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,
a4696,a4698,a4700,a4702,a4704,a4706,a4708,a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,
a4726,a4728,a4730,a4732,a4734,a4736,a4738,a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,
a4756,a4758,a4760,a4762,a4764,a4766,a4768,a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4784,
a4786,a4788,a4790,a4792,a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,
a4820,a4822,a4824,a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,a4844,a4848,a4850,
a4852,a4854,a4856,a4860,a4862,a4864,a4866,a4868,a4870,a4872,a4874,a4876,a4878,a4880,a4882,
a4884,a4886,a4888,a4890,a4892,a4894,a4896,a4898,a4900,a4902,a4904,a4906,a4908,a4910,a4912,
a4914,a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,a4938,a4940,a4942,
a4944,a4946,a4948,a4950,a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,a4968,a4970,a4972,
a4974,a4976,a4978,a4980,a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,a4998,a5000,a5002,
a5004,a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,a5028,a5030,a5032,
a5034,a5036,a5038,a5040,a5042,a5044,a5046,a5048,a5050,a5052,a5054,a5056,a5058,a5060,a5062,
a5064,a5066,a5068,a5070,a5072,a5074,a5076,a5078,a5080,a5082,a5084,a5086,a5088,a5090,a5092,
a5094,a5096,a5098,a5100,a5102,a5104,a5106,a5108,a5110,a5112,a5114,a5116,a5118,a5120,a5122,
a5124,a5126,a5128,a5130,a5132,a5134,a5136,a5138,a5140,a5142,a5144,a5146,a5148,a5150,a5152,
a5154,a5156,a5158,a5160,a5162,a5164,a5166,a5168,a5170,a5172,a5174,a5176,a5178,a5180,a5182,
a5186,a5188,a5190,a5192,a5196,a5198,a5200,a5202,a5206,a5208,a5210,a5212,a5216,a5218,a5220,
a5224,a5226,a5228,a5230,a5232,a5234,a5236,a5238,a5240,a5242,a5244,a5246,a5248,a5250,a5252,
a5254,a5256,a5258,a5260,a5262,a5264,a5266,a5268,a5270,a5272,a5274,a5276,a5278,a5282,a5284,
a5286,a5288,a5290,a5292,a5294,a5298,a5300,a5302,a5304,a5306,a5308,a5310,a5312,a5314,a5316,
a5318,a5320,a5322,a5326,a5328,a5330,a5332,a5334,a5336,a5338,a5340,a5342,a5344,a5346,a5348,
a5350,a5352,a5354,a5356,a5358,a5360,a5362,a5364,a5366,a5370,a5372,a5374,a5376,a5378,a5380,
a5382,a5386,a5388,a5390,a5392,a5394,a5396,a5398,a5400,a5402,a5406,a5408,a5410,a5412,a5414,
a5416,a5418,a5420,a5422,a5424,a5426,a5428,a5430,a5432,a5434,a5436,a5438,a5440,a5442,a5444,
a5446,a5450,a5452,a5454,a5456,a5458,a5460,a5462,a5466,a5468,a5470,a5472,a5474,a5476,a5478,
a5480,a5482,a5486,a5488,a5490,a5492,a5494,a5496,a5498,a5500,a5502,a5504,a5506,a5508,a5510,
a5512,a5514,a5516,a5518,a5520,a5522,a5524,a5526,a5530,a5532,a5534,a5536,a5538,a5540,a5542,
a5546,a5548,a5550,a5552,a5554,a5556,a5558,a5560,a5562,a5566,a5568,a5570,a5572,a5574,a5576,
a5578,a5580,a5582,a5584,a5586,a5588,a5590,a5592,a5594,a5596,a5598,a5600,a5602,a5604,a5606,
a5608,a5610,a5612,a5614,a5616,a5618,a5620,a5622,a5624,a5626,a5628,a5630,a5632,a5634,a5636,
a5638,a5640,a5642,a5644,a5646,a5648,a5650,a5652,a5654,a5656,a5658,a5660,a5662,a5664,a5666,
a5668,a5670,a5672,a5674,a5676,a5678,a5682,a5684,a5686,a5688,a5690,a5692,a5694,a5696,a5698,
a5700,a5702,a5706,a5708,a5710,a5712,a5714,a5716,a5718,a5720,a5722,a5724,a5726,a5728,a5730,
a5734,a5736,a5738,a5740,a5742,a5746,a5748,a5750,a5752,a5754,a5756,a5758,a5760,a5762,a5764,
a5766,a5768,a5770,a5772,a5774,a5776,a5778,a5780,a5782,a5784,a5786,a5788,a5790,a5792,a5794,
a5796,a5798,a5800,a5802,a5804,a5806,a5808,a5810,a5812,a5814,a5816,a5818,a5820,a5822,a5824,
a5826,a5828,a5830,a5832,a5834,a5836,a5838,a5840,a5842,a5844,a5846,a5848,a5850,a5852,a5854,
a5856,a5858,a5860,a5862,a5864,a5866,a5868,a5870,a5872,a5874,a5876,a5878,a5880,a5882,a5884,
a5886,a5888,a5890,a5892,a5894,a5896,a5898,a5900,a5902,a5904,a5906,a5908,a5910,a5912,a5914,
a5916,a5918,a5920,a5922,a5924,a5926,a5928,a5930,a5932,a5934,a5936,a5938,a5940,a5942,a5944,
a5946,a5948,a5950,a5952,a5954,a5956,a5958,a5960,a5962,a5964,a5966,a5968,a5970,a5972,a5974,
a5976,a5978,a5980,a5982,a5984,a5986,a5988,a5990,a5992,a5994,a5996,a5998,a6000,a6002,a6004,
a6006,a6008,a6010,a6012,a6014,a6016,a6018,a6020,a6022,a6024,a6026,a6028,a6030,a6032,a6034,
a6036,a6038,a6040,a6042,a6044,a6046,a6048,a6050,a6052,a6054,a6056,a6058,a6060,a6062,a6064,
a6066,a6068,a6072,a6074,a6076,a6078,a6082,a6084,a6086,a6088,a6092,a6094,a6096,a6098,a6102,
a6104,a6106,a6110,a6112,a6116,a6118,a6120,a6124,a6126,a6128,a6130,a6134,a6136,a6138,a6144,
a6146,a6148,a6150,a6152,a6154,a6156,a6158,a6160,a6162,a6164,a6166,a6168,a6170,a6172,a6174,
a6176,a6178,a6180,a6182,a6184,a6186,a6188,a6190,a6192,a6194,a6196,a6198,a6200,a6202,a6204,
a6206,a6208,a6210,a6212,a6214,a6216,a6218,a6220,a6222,a6224,a6226,a6228,a6230,a6232,a6234,
a6236,a6238,a6240,a6242,a6244,a6246,a6248,a6250,a6252,a6254,a6256,a6258,a6260,a6262,a6264,
a6266,a6268,a6270,a6272,a6274,a6276,a6278,a6280,a6282,a6284,a6286,a6288,a6290,a6292,a6294,
a6296,a6298,a6300,a6302,a6304,a6306,a6308,a6310,a6312,a6314,a6316,a6318,a6320,a6322,a6324,
a6326,a6328,a6330,a6332,a6334,a6336,a6338,a6340,a6342,a6344,a6346,a6348,a6350,a6352,a6354,
a6356,a6358,a6360,a6362,a6364,a6366,a6368,a6370,a6372,a6374,a6376,a6378,a6380,a6382,a6384,
a6386,a6388,a6390,a6392,a6394,a6396,a6398,a6400,a6402,a6404,a6406,a6408,a6410,a6412,a6414,
a6416,a6418,a6420,a6422,a6424,a6426,a6428,a6430,a6432,a6434,a6436,a6438,a6440,a6442,a6444,
a6446,a6448,a6450,a6452,a6454,a6456,a6458,a6460,a6462,a6464,a6466,a6468,a6470,a6472,a6474,
a6476,a6478,a6480,a6482,a6484,a6486,a6488,a6490,a6492,a6494,a6496,a6498,a6500,a6502,a6504,
a6506,a6508,a6510,a6512,a6514,a6516,a6518,a6520,a6522,a6524,a6526,a6528,a6530,a6532,a6534,
a6536,a6538,a6540,a6542,a6544,a6546,a6548,a6550,a6552,a6554,a6556,a6558,a6560,a6562,a6564,
a6566,a6568,a6570,a6572,a6574,a6576,a6578,a6580,a6582,a6584,a6586,a6588,a6590,a6592,a6594,
a6596,a6598,a6600,a6602,a6604,a6606,a6608,a6610,a6612,a6614,a6616,a6618,a6620,a6622,a6624,
a6626,a6628,a6630,a6632,a6634,a6636,a6638,a6640,a6642,a6644,a6646,a6648,a6650,a6652,a6654,
a6656,a6658,a6660,a6662,a6664,a6666,a6668,a6670,a6672,a6674,a6676,a6678,a6680,a6682,a6684,
a6686,a6688,a6690,a6692,a6694,a6696,a6698,a6700,a6702,a6704,a6706,a6708,a6710,a6712,a6714,
a6716,a6718,a6720,a6722,a6724,a6726,a6728,a6730,a6732,a6734,a6736,a6738,a6740,a6742,a6744,
a6746,a6748,a6750,a6752,a6754,a6756,a6758,a6760,a6762,a6764,a6766,a6768,a6770,a6772,a6774,
a6776,a6778,a6780,a6782,a6784,a6786,a6788,a6790,a6792,a6794,a6796,a6798,a6800,a6802,a6804,
a6806,a6808,a6810,a6812,a6814,a6816,a6818,a6820,a6822,a6824,a6826,a6828,a6830,a6832,a6834,
a6836,a6838,a6840,a6842,a6844,a6846,a6848,a6850,a6852,a6854,a6856,a6858,a6860,a6862,a6864,
a6866,a6868,a6870,a6872,a6874,a6876,a6878,a6880,a6882,a6884,a6886,a6888,a6890,a6892,a6894,
a6896,a6898,a6900,a6902,a6904,a6906,a6908,a6910,a6912,a6914,a6916,a6918,a6920,a6922,a6924,
a6926,a6928,a6930,a6932,a6934,a6936,a6938,a6940,a6942,a6944,a6946,a6948,a6950,a6952,a6954,
a6956,a6958,a6960,a6962,a6964,a6966,a6968,a6970,a6972,a6974,a6976,a6978,a6980,a6982,a6984,
a6986,a6988,a6990,a6992,a6994,a6996,a6998,a7000,a7002,a7004,a7006,a7008,a7010,a7012,a7014,
a7016,a7018,a7020,a7022,a7024,a7026,a7028,a7030,a7032,a7034,a7036,a7038,a7040,a7042,a7044,
a7046,a7048,a7050,a7052,a7054,a7056,a7058,a7060,a7062,a7064,a7066,a7068,a7070,a7072,a7074,
a7076,a7078,a7080,a7082,a7084,a7086,a7088,a7090,a7092,a7094,a7096,a7098,a7100,a7102,a7104,
a7106,a7108,a7110,a7112,a7114,a7116,a7118,a7120,a7122,a7124,a7126,a7128,a7130,a7132,a7134,
a7136,a7138,a7140,a7142,a7144,a7146,a7148,a7150,a7152,a7154,a7156,a7158,a7160,a7162,a7164,
a7166,a7168,a7170,a7172,a7174,a7176,a7178,a7180,a7182,a7184,a7186,a7188,a7190,a7192,a7194,
a7196,a7198,a7200,a7202,a7204,a7206,a7208,a7210,a7212,a7214,a7216,a7218,a7220,a7222,a7224,
a7226,a7228,a7230,a7232,a7234,a7236,a7238,a7240,a7242,a7244,a7246,a7248,a7250,a7252,a7254,
a7256,a7258,a7260,a7262,a7264,a7266,a7268,a7270,a7272,a7274,a7276,a7278,a7280,a7282,a7284,
a7286,a7288,a7290,a7292,a7294,a7296,a7298,a7300,a7302,a7304,a7306,a7308,a7310,a7312,a7314,
a7316,a7318,a7320,a7322,a7324,a7326,a7328,a7330,a7332,a7334,a7336,a7338,a7340,a7342,a7344,
a7346,a7348,a7350,a7352,a7354,a7356,a7358,a7360,a7362,a7364,a7366,a7368,a7370,a7372,a7374,
a7376,a7378,a7380,a7382,a7384,a7386,a7388,a7390,a7392,a7394,a7396,a7398,a7400,a7402,a7404,
a7406,a7408,a7410,a7412,a7414,a7416,a7418,a7420,a7422,a7424,a7426,a7428,a7430,a7432,a7434,
a7436,a7438,a7440,a7442,a7444,a7446,a7448,a7450,a7452,a7454,a7456,a7458,a7460,a7462,a7464,
a7466,a7468,a7470,a7472,a7474,a7476,a7478,a7480,a7482,a7484,a7486,a7488,a7490,a7492,a7494,
a7496,a7498,a7500,a7502,a7504,a7506,a7508,a7510,a7512,a7514,a7516,a7518,a7520,a7522,a7524,
a7526,a7528,a7530,a7532,a7534,a7536,a7538,a7540,a7542,a7544,a7546,a7548,a7550,a7552,a7554,
a7556,a7558,a7560,a7562,a7564,a7566,a7568,a7570,a7572,a7574,a7576,a7578,a7580,a7582,a7584,
a7586,a7588,a7590,a7592,a7594,a7596,a7598,a7600,a7602,a7604,a7606,a7608,a7610,a7612,a7614,
a7616,a7618,a7620,a7622,a7624,a7626,a7628,a7630,a7632,a7634,a7636,a7638,a7640,a7642,a7644,
a7646,a7648,a7650,a7652,a7654,a7656,a7658,a7660,a7662,a7664,a7666,a7668,a7670,a7672,a7674,
a7676,a7678,a7680,a7682,a7684,a7686,a7688,a7690,a7692,a7694,a7696,a7698,a7700,a7702,a7704,
a7706,a7708,a7710,a7712,a7714,a7716,a7718,a7720,a7722,a7724,a7726,a7728,a7730,a7732,a7734,
a7736,a7738,a7740,a7742,a7744,a7746,a7748,a7750,a7752,a7754,a7756,a7758,a7760,a7762,a7764,
a7766,a7768,a7770,a7772,a7774,a7776,a7778,a7780,a7782,a7784,a7786,a7788,a7790,a7792,a7794,
a7796,a7798,a7800,a7802,a7804,a7806,a7808,a7810,a7812,a7814,a7816,a7818,a7820,a7822,a7824,
a7826,a7828,a7830,a7832,a7834,a7836,a7838,a7840,a7842,a7844,a7846,a7848,a7850,a7852,a7854,
a7856,a7858,a7860,a7862,a7864,a7866,a7868,a7870,a7872,a7874,a7876,a7878,a7880,a7882,a7884,
a7886,a7888,a7890,a7892,a7894,a7896,a7898,a7900,a7902,a7904,a7906,a7908,a7910,a7912,a7914,
a7916,a7918,a7920,a7922,a7924,a7926,a7928,a7930,a7932,a7934,a7936,a7938,a7940,a7942,a7944,
a7946,a7948,a7950,a7952,a7954,a7956,a7958,a7960,a7962,a7964,a7966,a7968,a7970,a7972,a7974,
a7976,a7978,a7980,a7982,a7984,a7986,a7988,a7990,a7992,a7994,a7996,a7998,a8000,a8002,a8004,
a8006,a8008,a8010,a8012,a8014,a8016,a8018,a8020,a8022,a8024,a8026,a8028,a8030,a8032,a8034,
a8036,a8038,a8040,a8042,a8044,a8046,a8048,a8050,a8052,a8054,a8056,a8058,a8060,a8062,a8064,
a8066,a8068,a8070,a8072,a8074,a8076,a8078,a8080,a8082,a8084,a8086,a8088,a8090,a8092,a8094,
a8096,a8098,a8100,a8102,a8104,a8106,a8108,a8110,a8112,a8114,a8116,a8118,a8120,a8122,a8124,
a8126,a8128,a8130,a8132,a8134,a8136,a8138,a8140,a8142,a8144,a8146,a8148,a8150,a8152,a8154,
a8156,a8158,a8160,a8162,a8164,a8166,a8168,a8170,a8172,a8174,a8176,a8178,a8180,a8182,a8184,
a8186,a8188,a8190,a8192,a8194,a8196,a8198,a8200,a8202,a8204,a8206,a8208,a8210,a8212,a8214,
a8216,a8218,a8220,a8222,a8224,a8226,a8228,a8230,a8232,a8234,a8236,a8238,a8240,a8242,a8244,
a8246,a8248,a8250,a8252,a8254,a8256,a8258,a8260,a8262,a8264,a8266,a8268,a8270,a8272,a8274,
a8276,a8278,a8280,a8282,a8284,a8286,a8288,a8290,a8292,a8294,a8296,a8298,a8300,a8302,a8304,
a8306,a8308,a8310,a8312,a8314,a8316,a8318,a8320,a8322,a8324,a8326,a8328,a8330,a8332,a8334,
a8336,a8338,a8340,a8342,a8344,a8346,a8348,a8350,a8352,a8354,a8356,a8358,a8360,a8362,a8364,
a8366,a8368,a8370,a8372,a8374,a8376,a8378,a8380,a8382,a8384,a8386,a8388,a8390,a8392,a8394,
a8396,a8398,a8400,a8402,a8404,a8406,a8408,a8410,a8412,a8414,a8416,a8418,a8420,a8422,a8424,
a8426,a8428,a8430,a8432,a8434,a8436,a8438,a8440,a8442,a8444,a8446,a8448,a8450,a8452,a8454,
a8456,a8458,a8460,a8462,a8464,a8466,a8468,a8470,a8472,a8474,a8476,a8478,a8480,a8482,a8484,
a8486,a8488,a8490,a8492,a8494,a8496,a8498,a8500,a8502,a8504,a8506,a8508,a8510,a8512,a8514,
a8516,a8518,a8520,a8522,a8524,a8526,a8528,a8530,a8532,a8534,a8536,a8538,a8540,a8542,a8544,
a8546,a8548,a8550,a8552,a8554,a8556,a8558,a8560,a8562,a8564,a8566,a8568,a8570,a8572,a8574,
a8576,a8578,a8580,a8582,a8584,a8586,a8588,a8590,a8592,a8594,a8596,a8598,a8600,a8602,a8604,
a8606,a8608,a8610,a8612,a8614,a8616,a8618,a8620,a8622,a8624,a8626,a8628,a8630,a8632,a8634,
a8636,a8638,a8640,a8642,a8644,a8646,a8648,a8650,a8652,a8654,a8656,a8658,a8660,a8662,a8664,
a8666,a8668,a8670,a8672,a8674,a8676,a8678,a8680,a8682,a8684,a8686,a8688,a8690,a8692,a8694,
a8696,a8698,a8700,a8702,a8704,a8706,a8708,a8710,a8712,a8714,a8716,a8718,a8720,a8722,a8724,
a8726,a8728,a8730,a8732,a8734,a8736,a8738,a8740,a8742,a8744,a8746,a8748,a8750,a8752,a8754,
a8756,a8758,a8760,a8762,a8764,a8766,a8768,a8770,a8772,a8774,a8776,a8778,a8780,a8782,a8784,
a8786,a8788,a8790,a8792,a8794,a8796,a8798,a8800,a8802,a8804,a8806,a8808,a8810,a8812,a8814,
a8816,a8818,a8820,a8822,a8824,a8826,a8828,a8830,a8832,a8834,a8836,a8838,a8840,a8842,a8844,
a8846,a8848,a8850,a8852,a8854,a8856,a8858,a8860,a8862,a8864,a8866,a8868,a8870,a8872,a8874,
a8876,a8878,a8880,a8882,a8884,a8886,a8888,a8890,a8892,a8894,a8896,a8898,a8900,a8902,a8904,
a8906,a8908,a8910,a8912,a8914,a8916,a8918,a8920,a8922,a8924,a8926,a8928,a8930,a8932,a8934,
a8936,a8938,a8940,a8942,a8944,a8946,a8948,a8950,a8952,a8954,a8956,a8958,a8960,a8962,a8964,
a8966,a8968,a8970,a8972,a8974,a8976,a8978,a8980,a8982,a8984,a8986,a8988,a8990,a8992,a8994,
a8996,a8998,a9000,a9002,a9004,a9006,a9008,a9010,a9012,a9014,a9016,a9018,a9020,a9022,a9024,
a9026,a9028,a9030,a9032,a9034,a9036,a9038,a9040,a9042,a9044,a9046,a9048,a9050,a9052,a9054,
a9056,a9058,a9060,a9062,a9064,a9066,a9068,a9070,a9072,a9074,a9076,a9078,a9080,a9082,a9084,
a9086,a9088,a9090,a9092,a9094,a9096,a9098,a9100,a9102,a9104,a9106,a9108,a9110,a9112,a9114,
a9116,a9118,a9120,a9122,a9124,a9126,a9128,a9130,a9132,a9134,a9136,a9138,a9140,a9142,a9144,
a9146,a9148,a9150,a9152,a9154,a9156,a9158,a9160,a9162,a9164,a9166,a9168,a9170,a9172,a9174,
a9176,a9178,a9180,a9182,a9184,a9186,a9188,a9190,a9192,a9194,a9196,a9198,a9200,a9202,a9204,
a9206,a9208,a9210,a9212,a9214,a9216,a9218,a9220,a9222,a9224,a9226,a9228,a9230,a9232,a9234,
a9236,a9238,a9240,a9242,a9244,a9246,a9248,a9250,a9252,a9254,a9256,a9258,a9260,a9262,a9264,
a9266,a9268,a9270,a9272,a9274,a9276,a9278,a9280,a9282,a9284,a9286,a9288,a9290,a9292,a9294,
a9296,a9298,a9300,a9302,a9304,a9306,a9308,a9310,a9312,a9314,a9316,a9318,a9320,a9322,a9324,
a9326,a9328,a9330,a9332,a9334,a9336,a9338,a9340,a9342,a9344,a9346,a9348,a9350,a9352,a9354,
a9356,a9358,a9360,a9362,a9364,a9366,a9368,a9370,a9372,a9374,a9376,a9378,a9380,a9382,a9384,
a9386,a9388,a9390,a9392,a9394,a9396,a9398,a9400,a9402,a9404,a9406,a9408,a9410,a9412,a9414,
a9416,a9418,a9420,a9422,a9424,a9426,a9428,a9430,a9432,a9434,a9436,a9438,a9440,a9442,a9444,
a9446,a9448,a9450,a9452,a9454,a9456,a9458,a9460,a9462,a9464,a9466,a9468,a9470,a9472,a9474,
a9476,a9478,a9480,a9482,a9484,a9486,a9488,a9490,a9492,a9494,a9496,a9498,a9500,a9502,a9504,
a9506,a9508,a9510,a9512,a9514,a9516,a9518,a9520,a9522,a9524,a9526,a9528,a9530,a9532,a9534,
a9536,a9538,a9540,a9542,a9544,a9546,a9548,a9550,a9552,a9554,a9556,a9558,a9560,a9562,a9564,
a9566,a9568,a9570,a9572,a9574,a9576,a9578,a9580,a9582,a9584,a9586,a9588,a9590,a9592,a9594,
a9596,a9598,a9600,a9602,a9604,a9606,a9608,a9610,a9612,a9614,a9616,a9618,a9620,a9622,a9624,
a9626,a9628,a9630,a9632,a9634,a9636,a9638,a9640,a9642,a9644,a9646,a9648,a9650,a9652,a9654,
a9656,a9658,a9660,a9662,a9664,a9666,a9668,a9670,a9672,a9674,a9676,a9678,a9680,a9682,a9684,
a9686,a9688,a9690,a9692,a9694,a9696,a9698,a9700,a9702,a9704,a9706,a9708,a9710,a9712,a9714,
a9716,a9718,a9720,a9722,a9724,a9726,a9728,a9730,a9732,a9734,a9736,a9738,a9740,a9742,a9744,
a9746,a9748,a9750,a9752,a9754,a9756,a9758,a9760,a9762,a9764,a9766,a9768,a9770,a9772,a9774,
a9776,a9778,a9780,a9782,a9784,a9786,a9788,a9790,a9792,a9794,a9796,a9798,a9800,a9802,a9804,
a9806,a9808,a9810,a9812,a9814,a9816,a9818,a9820,a9822,a9824,a9826,a9828,a9830,a9832,a9834,
a9836,a9838,a9840,a9842,a9844,a9846,a9848,a9850,a9852,a9854,a9856,a9858,a9860,a9862,a9864,
a9866,a9868,a9870,a9872,a9874,a9876,a9878,a9880,a9882,a9884,a9886,a9888,a9890,a9892,a9894,
a9896,a9898,a9900,a9902,a9904,a9906,a9908,a9910,a9912,a9914,a9916,a9918,a9920,a9922,a9924,
a9926,a9928,a9930,a9932,a9934,a9936,a9938,a9940,a9942,a9944,a9946,a9948,a9950,a9952,a9954,
a9956,a9958,a9960,a9962,a9964,a9966,a9968,a9970,a9972,a9974,a9976,a9978,a9980,a9982,a9984,
a9986,a9988,a9990,a9992,a9994,a9996,a9998,a10000,a10002,a10004,a10006,a10008,a10010,a10012,a10014,
a10016,a10018,a10020,a10022,a10024,a10026,a10028,a10030,a10032,a10034,a10036,a10038,a10040,a10042,a10044,
a10046,a10048,a10050,a10052,a10054,a10056,a10058,a10060,a10062,a10064,a10066,a10068,a10070,a10072,a10074,
a10076,a10078,a10080,a10082,a10084,a10086,a10088,a10090,a10092,a10094,a10096,a10098,a10100,a10102,a10104,
a10106,a10108,a10110,a10112,a10114,a10116,a10118,a10120,a10122,a10124,a10126,a10128,a10130,a10132,a10134,
a10136,a10138,a10140,a10142,a10144,a10146,a10148,a10150,a10152,a10154,a10156,a10158,a10160,a10162,a10164,
a10166,a10168,a10170,a10172,a10174,a10176,a10178,a10180,a10182,a10184,a10186,a10188,a10190,a10192,a10194,
a10196,a10198,a10200,a10202,a10204,a10206,a10208,a10210,a10212,a10214,a10216,a10218,a10220,a10222,a10224,
a10226,a10228,a10230,a10232,a10234,a10236,a10238,a10240,a10242,a10244,a10246,a10248,a10250,a10252,a10254,
a10256,a10258,a10260,a10262,a10264,a10266,a10268,a10270,a10272,a10274,a10276,a10278,a10280,a10282,a10284,
a10286,a10288,a10290,a10292,a10294,a10296,a10298,a10300,a10302,a10304,a10306,a10308,a10310,a10312,a10314,
a10316,a10318,a10320,a10322,a10324,a10326,a10328,a10330,a10332,a10334,a10336,a10338,a10340,a10342,a10344,
a10346,a10348,a10350,a10352,a10354,a10356,a10358,a10360,a10362,a10364,a10366,a10368,a10370,a10372,a10374,
a10376,a10378,a10380,a10382,a10384,a10386,a10388,a10390,a10392,a10394,a10396,a10398,a10400,a10402,a10404,
a10406,a10408,a10410,a10412,a10414,a10416,a10418,a10420,a10422,a10424,a10426,a10428,a10430,a10432,a10434,
a10436,a10438,a10440,a10442,a10444,a10446,a10448,a10450,a10452,a10454,a10456,a10458,a10460,a10462,a10464,
a10466,a10468,a10470,a10472,a10474,a10476,a10478,a10480,a10482,a10484,a10486,a10488,a10490,a10492,a10494,
a10496,a10498,a10500,a10502,a10504,a10506,a10508,a10510,a10512,a10514,a10516,a10518,a10520,a10522,a10524,
a10526,a10528,a10530,a10532,a10534,a10536,a10538,a10540,a10542,a10544,a10546,a10548,a10550,a10552,a10554,
a10556,a10558,a10560,a10562,a10564,a10566,a10568,a10570,a10572,a10574,a10576,a10578,a10580,a10582,a10584,
a10586,a10588,a10590,a10592,a10594,a10596,a10598,a10600,a10602,a10604,a10606,a10608,a10610,a10612,a10614,
a10616,a10618,a10620,a10622,a10624,a10626,a10628,a10630,a10632,a10634,a10636,a10638,a10640,a10642,a10644,
a10646,a10648,a10650,a10652,a10654,a10656,a10658,a10660,a10662,a10664,a10666,a10668,a10670,a10672,a10674,
a10676,a10678,a10680,a10682,a10684,a10686,a10688,a10690,a10692,a10694,a10696,a10698,a10700,a10702,a10704,
a10706,a10708,a10710,a10712,a10714,a10716,a10718,a10720,a10722,a10724,a10726,a10728,a10730,a10732,a10734,
a10736,a10738,a10740,a10742,a10744,a10746,a10748,a10750,a10752,a10754,a10756,a10758,a10760,a10762,a10764,
a10766,a10768,a10770,a10772,a10774,a10776,a10778,a10780,a10782,a10784,a10786,a10788,a10790,a10792,a10794,
a10796,a10798,a10800,a10802,a10804,a10806,a10808,a10810,a10812,a10814,a10816,a10818,a10820,a10822,a10824,
a10826,a10828,a10830,a10832,a10834,a10836,a10838,a10840,a10842,a10844,a10846,a10848,a10850,a10852,a10854,
a10856,a10858,a10860,a10862,a10864,a10866,a10868,a10870,a10872,a10874,a10876,a10878,a10880,a10882,a10884,
a10886,a10888,a10890,a10892,a10894,a10896,a10898,a10900,a10902,a10904,a10906,a10908,a10910,a10912,a10914,
a10916,a10918,a10920,a10922,a10924,a10926,a10928,a10930,a10932,a10934,a10936,a10938,a10940,a10942,a10944,
a10946,a10948,a10950,a10952,a10954,a10956,a10958,a10960,a10962,a10964,a10966,a10968,a10970,a10972,a10974,
a10976,a10978,a10980,a10982,a10984,a10986,a10988,a10990,a10992,a10994,a10996,a10998,a11000,a11002,a11004,
a11006,a11008,a11010,a11012,a11014,a11016,a11018,a11020,a11022,a11024,a11026,a11028,a11030,a11032,a11034,
a11036,a11038,a11040,a11042,a11044,a11046,a11048,a11050,a11052,a11054,a11056,a11058,a11060,a11062,a11064,
a11066,a11068,a11070,a11072,a11074,a11076,a11078,a11080,a11082,a11084,a11086,a11088,a11090,a11092,a11094,
a11096,a11098,a11100,a11102,a11104,a11106,a11108,a11110,a11112,a11114,a11116,a11118,a11120,a11122,a11124,
a11126,a11128,a11130,a11132,a11134,a11136,a11138,a11140,a11142,a11144,a11146,a11148,a11150,a11152,a11154,
a11156,a11158,a11160,a11162,a11164,a11166,a11168,a11170,a11172,a11174,a11176,a11178,a11180,a11182,a11184,
a11186,a11188,a11190,a11192,a11194,a11196,a11198,a11200,a11202,a11204,a11206,a11208,a11210,a11212,a11214,
a11216,a11218,a11220,a11222,a11224,a11226,a11228,a11230,a11232,a11234,a11236,a11238,a11240,a11242,a11244,
a11246,a11248,a11250,a11252,a11254,a11256,a11258,a11260,a11262,a11264,a11266,a11268,a11270,a11272,a11274,
a11276,a11278,a11280,a11282,a11284,a11286,a11288,a11290,a11292,a11294,a11296,a11298,a11300,a11302,a11304,
a11306,a11308,a11310,a11312,a11314,a11316,a11318,a11320,a11322,a11324,a11326,a11328,a11330,a11332,a11334,
a11336,a11338,a11340,a11342,a11344,a11346,a11348,a11350,a11352,a11354,a11356,a11358,a11360,a11362,a11364,
a11366,a11368,a11370,a11372,a11374,a11376,a11378,a11380,a11382,a11384,a11386,a11388,a11390,a11392,a11394,
a11396,a11398,a11400,a11402,a11404,a11406,a11408,a11410,a11412,a11414,a11416,a11418,a11420,a11422,a11424,
a11426,a11428,a11430,a11432,a11434,a11436,a11438,a11440,a11442,a11444,a11446,a11448,a11450,a11452,a11454,
a11456,a11458,a11460,a11462,a11464,a11466,a11468,a11470,a11472,a11474,a11476,a11478,a11480,a11482,a11484,
a11486,a11488,a11490,a11492,a11494,a11496,a11498,a11500,a11502,a11504,a11506,a11508,a11510,a11512,a11514,
a11516,a11518,a11520,a11522,a11524,a11526,a11528,a11530,a11532,a11534,a11536,a11538,a11540,a11542,a11544,
a11546,a11548,a11550,a11552,a11554,a11556,a11558,a11560,a11562,a11564,a11566,a11568,a11570,a11572,a11574,
a11576,a11578,a11580,a11582,a11584,a11586,a11588,a11590,a11592,a11594,a11596,a11598,a11600,a11602,a11604,
a11606,a11608,a11610,a11612,a11614,a11616,a11618,a11620,a11622,a11624,a11626,a11628,a11630,a11632,a11634,
a11636,a11638,a11640,a11642,a11644,a11646,a11648,a11650,a11652,a11654,a11656,a11658,a11660,a11662,a11664,
a11666,a11668,a11670,a11672,a11674,a11676,a11678,a11680,a11682,a11684,a11686,a11688,a11690,a11692,a11694,
a11696,a11698,a11700,a11702,a11704,a11706,a11708,a11710,a11712,a11714,a11716,a11718,a11720,a11722,a11724,
a11726,a11728,a11730,a11732,a11734,a11736,a11738,a11740,a11742,a11744,a11746,a11748,a11750,a11752,a11754,
a11756,a11758,a11760,a11762,a11764,a11766,a11768,a11770,a11772,a11774,a11776,a11778,a11780,a11782,a11784,
a11786,a11788,a11790,a11792,a11794,a11796,a11798,a11800,a11802,a11804,a11806,a11808,a11810,a11812,a11814,
a11816,a11818,a11820,a11822,a11824,a11826,a11828,a11830,a11832,a11834,a11836,a11838,a11840,a11842,a11844,
a11846,a11848,a11850,a11852,a11854,a11856,a11858,a11860,a11862,a11864,a11866,a11868,a11870,a11872,a11874,
a11876,a11878,a11880,a11882,a11884,a11886,a11888,a11890,a11892,a11894,a11896,a11898,a11900,a11902,a11904,
a11906,a11908,a11910,a11912,a11914,a11916,a11918,a11920,a11922,a11924,a11926,a11928,a11930,a11932,a11934,
a11936,a11938,a11940,a11942,a11944,a11946,a11948,a11950,a11952,a11954,a11956,a11958,a11960,a11962,a11964,
a11966,a11968,a11970,a11972,a11974,a11976,a11978,a11980,a11982,a11984,a11986,a11988,a11990,a11992,a11994,
a11996,a11998,a12000,a12002,a12004,a12006,a12008,a12010,a12012,a12014,a12016,a12018,a12020,a12022,a12024,
a12026,a12028,a12030,a12032,a12034,a12036,a12038,a12040,a12042,a12044,a12046,a12048,a12050,a12052,a12054,
a12056,a12058,a12060,a12062,a12064,a12066,a12068,a12070,a12072,a12074,a12076,a12078,a12080,a12082,a12084,
a12086,a12088,a12090,a12092,a12094,a12096,a12098,a12100,a12102,a12104,a12106,a12108,a12110,a12112,a12114,
a12116,a12118,a12120,a12122,a12124,a12126,a12128,a12130,a12132,a12134,a12136,a12138,a12140,a12142,a12144,
a12146,a12148,a12150,a12152,a12154,a12156,a12158,a12160,a12162,a12164,a12166,a12168,a12170,a12172,a12174,
a12176,a12178,a12180,a12182,a12184,a12186,a12188,a12190,a12192,a12194,a12196,a12198,a12200,a12202,a12204,
a12206,a12208,a12210,a12212,a12214,a12216,a12218,a12220,a12222,a12224,a12226,a12228,a12230,a12232,a12234,
a12236,a12238,a12240,a12242,a12244,a12246,a12248,a12250,a12252,a12254,a12256,a12258,a12260,a12262,a12264,
a12266,a12268,a12270,a12272,a12274,a12276,a12278,a12280,a12282,a12284,a12286,a12288,a12290,a12292,a12294,
a12296,a12298,a12300,a12302,a12304,a12306,a12308,a12310,a12312,a12314,a12316,a12318,a12320,a12322,a12324,
a12326,a12328,a12330,a12332,a12334,a12336,a12338,a12340,a12342,a12344,a12346,a12348,a12350,a12352,a12354,
a12356,a12358,a12360,a12362,a12364,a12366,a12368,a12370,a12372,a12374,a12376,a12378,a12380,a12382,a12384,
a12386,a12388,a12390,a12392,a12394,a12396,a12398,a12400,a12402,a12404,a12406,a12408,a12410,a12412,a12414,
a12416,a12418,a12420,a12422,a12424,a12426,a12428,a12430,a12432,a12434,a12436,a12438,a12440,a12442,a12444,
a12446,a12448,a12450,a12452,a12454,a12456,a12458,a12460,a12462,a12464,a12466,a12468,a12470,a12472,a12474,
a12476,a12478,a12480,a12482,a12484,a12486,a12488,a12490,a12492,a12494,a12496,a12498,a12500,a12502,a12504,
a12506,a12508,a12510,a12512,a12514,a12516,a12518,a12520,a12522,a12524,a12526,a12528,a12530,a12532,a12534,
a12536,a12538,a12540,a12542,a12544,a12546,a12548,a12550,a12552,a12554,a12556,a12558,a12560,a12562,a12564,
a12566,a12568,a12570,a12572,a12574,a12576,a12578,a12580,a12582,a12584,a12586,a12588,a12590,a12592,a12594,
a12596,a12598,a12600,a12602,a12604,a12606,a12608,a12610,a12612,a12614,a12616,a12618,a12620,a12622,a12624,
a12626,a12628,a12630,a12632,a12634,a12636,a12638,a12640,a12642,a12644,a12646,a12648,a12650,a12652,a12654,
a12656,a12658,a12660,a12662,a12664,a12666,a12668,a12670,a12672,a12674,a12676,a12678,a12680,a12682,a12684,
a12686,a12688,a12690,a12692,a12694,a12696,a12698,a12700,a12702,a12704,a12706,a12708,a12710,a12712,a12714,
a12716,a12718,a12720,a12722,a12724,a12726,a12728,a12730,a12732,a12734,a12736,a12738,a12740,a12742,a12744,
a12746,a12748,a12750,a12752,a12754,a12756,a12758,a12760,a12762,a12764,a12766,a12768,a12770,a12772,a12774,
a12776,a12778,a12780,a12782,a12784,a12786,a12788,a12790,a12792,a12794,a12796,a12798,a12800,a12802,a12804,
a12806,a12808,a12810,a12812,a12814,a12816,a12818,a12820,a12822,a12824,a12826,a12828,a12830,a12832,a12834,
a12836,a12838,a12840,a12842,a12844,a12846,a12848,a12850,a12852,a12854,a12856,a12858,a12860,a12862,a12864,
a12866,a12868,a12870,a12872,a12874,a12876,a12878,a12880,a12882,a12884,a12886,a12888,a12890,a12892,a12894,
a12896,a12898,a12900,a12902,a12904,a12906,a12908,a12910,a12912,a12914,a12916,a12918,a12920,a12922,a12924,
a12926,a12928,a12930,a12932,a12934,a12936,a12938,a12940,a12942,a12944,a12946,a12948,a12950,a12952,a12954,
a12956,a12958,a12960,a12962,a12964,a12966,a12968,a12970,a12972,a12974,a12976,a12978,a12980,a12982,a12984,
a12986,a12988,a12990,a12992,a12994,a12996,a12998,a13000,a13002,a13004,a13006,a13008,a13010,a13012,a13014,
a13016,a13018,a13020,a13022,a13024,a13026,a13028,a13030,a13032,a13034,a13036,a13038,a13040,a13042,a13044,
a13046,a13048,a13050,a13052,a13054,a13056,a13058,a13060,a13062,a13064,a13066,a13068,a13070,a13072,a13074,
a13076,a13078,a13080,a13082,a13084,a13086,a13088,a13090,a13092,a13094,a13096,a13098,a13100,a13102,a13104,
a13106,a13108,a13110,a13112,a13114,a13116,a13118,a13120,a13122,a13124,a13126,a13128,a13130,a13132,a13134,
a13136,a13138,a13140,a13142,a13144,a13146,a13148,a13150,a13152,a13154,a13156,a13158,a13160,a13162,a13164,
a13166,a13168,a13170,a13172,a13174,a13176,a13178,a13180,a13182,a13184,a13186,a13188,a13190,a13192,a13194,
a13196,a13198,a13200,a13202,a13204,a13206,a13208,a13210,a13212,a13214,a13216,a13218,a13220,a13222,a13224,
a13226,a13228,a13230,a13232,a13234,a13236,a13238,a13240,a13242,a13244,a13246,a13248,a13250,a13252,a13254,
a13256,a13258,a13260,a13262,a13264,a13266,a13268,a13270,a13272,a13274,a13276,a13278,a13280,a13282,a13284,
a13286,a13288,a13290,a13292,a13294,a13296,a13298,a13300,a13302,a13304,a13306,a13308,a13310,a13312,a13314,
a13316,a13318,a13320,a13322,a13324,a13326,a13328,a13330,a13332,a13334,a13336,a13338,a13340,a13342,a13344,
a13346,a13348,a13350,a13352,a13354,a13356,a13358,a13360,a13362,a13364,a13366,a13368,a13370,a13372,a13374,
a13376,a13378,a13380,a13382,a13384,a13386,a13388,a13390,a13392,a13394,a13396,a13398,a13400,a13402,a13404,
a13406,a13408,a13410,a13412,a13414,a13416,a13418,a13420,a13422,a13424,a13426,a13428,a13430,a13432,a13434,
a13436,a13438,a13440,a13442,a13444,a13446,a13448,a13450,a13452,a13454,a13456,a13458,a13460,a13462,a13464,
a13466,a13468,a13470,a13472,a13474,a13476,a13478,a13480,a13482,a13484,a13486,a13488,a13490,a13492,a13494,
a13496,a13498,a13500,a13502,a13504,a13506,a13508,a13510,a13512,a13514,a13516,a13518,a13520,a13522,a13524,
a13526,a13528,a13530,a13532,a13534,a13536,a13538,a13540,a13542,a13544,a13546,a13548,a13550,a13552,a13554,
a13556,a13558,a13560,a13562,a13564,a13566,a13568,a13570,a13572,a13574,a13576,a13578,a13580,a13582,a13584,
a13586,a13588,a13590,a13592,a13594,a13596,a13598,a13600,a13602,a13604,a13606,a13608,a13610,a13612,a13614,
a13616,a13618,a13620,a13622,a13624,a13626,a13628,a13630,a13632,a13634,a13636,a13638,a13640,a13642,a13644,
a13646,a13648,a13650,a13652,a13654,a13656,a13658,a13660,a13662,a13664,a13666,a13668,a13670,a13672,a13674,
a13676,a13678,a13680,a13682,a13684,a13686,a13688,a13690,a13692,a13694,a13696,a13698,a13700,a13702,a13704,
a13706,a13708,a13710,a13712,a13714,a13716,a13718,a13720,a13722,a13724,a13726,a13728,a13730,a13732,a13734,
a13736,a13738,a13740,a13742,a13744,a13746,a13748,a13750,a13752,a13754,a13756,a13758,a13760,a13762,a13764,
a13766,a13768,a13770,a13772,a13774,a13776,a13778,a13780,a13782,a13784,a13786,a13788,a13790,a13792,a13794,
a13796,a13798,a13800,a13802,a13804,a13806,a13808,a13810,a13812,a13814,a13816,a13818,a13820,a13822,a13824,
a13826,a13828,a13830,a13832,a13834,a13836,a13838,a13840,a13842,a13844,a13846,a13848,a13850,a13852,a13854,
a13856,a13858,a13860,a13862,a13864,a13866,a13868,a13870,a13872,a13874,a13876,a13878,a13880,a13882,a13884,
a13886,a13888,a13890,a13892,a13894,a13896,a13898,a13900,a13902,a13904,a13906,a13908,a13910,a13912,a13914,
a13916,a13918,a13920,a13922,a13924,a13926,a13928,a13930,a13932,a13934,a13936,a13938,a13940,a13942,a13944,
a13946,a13948,a13950,a13952,a13954,a13956,a13958,a13960,a13962,a13964,a13966,a13968,a13970,a13972,a13974,
a13976,a13978,a13980,a13982,a13984,a13986,a13988,a13990,a13992,a13994,a13996,a13998,a14000,a14002,a14004,
a14006,a14008,a14010,a14012,a14014,a14016,a14018,a14020,a14022,a14024,a14026,a14028,a14030,a14032,a14034,
a14036,a14038,a14040,a14042,a14044,a14046,a14048,a14050,a14052,a14054,a14056,a14058,a14060,a14062,a14064,
a14066,a14068,a14070,a14072,a14074,a14076,a14078,a14080,a14082,a14084,a14086,a14088,a14090,a14092,a14094,
a14096,a14098,a14100,a14102,a14104,a14106,a14108,a14110,a14112,a14114,a14116,a14118,a14120,a14122,a14124,
a14126,a14128,a14130,a14132,a14134,a14136,a14138,a14140,a14142,a14144,a14146,a14148,a14150,a14152,a14154,
a14156,a14158,a14160,a14162,a14164,a14166,a14168,a14170,a14172,a14174,a14176,a14178,a14180,a14182,a14184,
a14186,a14188,a14190,a14192,a14194,a14196,a14198,a14200,a14202,a14204,a14206,a14208,a14210,a14212,a14214,
a14216,a14218,a14220,a14222,a14224,a14226,a14228,a14230,a14232,a14234,a14236,a14238,a14240,a14242,a14244,
a14246,a14248,a14250,a14252,a14254,a14256,a14258,a14260,a14262,a14264,a14266,a14268,a14270,a14272,a14274,
a14276,a14278,a14280,a14282,a14284,a14286,a14288,a14290,a14292,a14294,a14296,a14298,a14300,a14302,a14304,
a14306,a14308,a14310,a14312,a14314,a14316,a14318,a14320,a14322,a14324,a14326,a14328,a14330,a14332,a14334,
a14336,a14338,a14340,a14342,a14344,a14346,a14348,a14350,a14352,a14354,a14356,a14358,a14360,a14362,a14364,
a14366,a14368,a14370,a14372,a14374,a14376,a14378,a14380,a14382,a14384,a14386,a14388,a14390,a14392,a14394,
a14396,a14398,a14400,a14402,a14404,a14406,a14408,a14410,a14412,a14414,a14416,a14418,a14420,a14422,a14424,
a14426,a14428,a14430,a14432,a14434,a14436,a14438,a14440,a14442,a14444,a14446,a14448,a14450,a14452,a14454,
a14456,a14458,a14460,a14462,a14464,a14466,a14468,a14470,a14472,a14474,a14476,a14478,a14480,a14482,a14484,
a14486,a14488,a14490,a14492,a14494,a14496,a14498,a14500,a14502,a14504,a14506,a14508,a14510,a14512,a14514,
a14516,a14518,a14520,a14522,a14524,a14526,a14528,a14530,a14532,a14534,a14536,a14538,a14540,a14542,a14544,
a14546,a14548,a14550,a14552,a14554,a14556,a14558,a14560,a14562,a14564,a14566,a14568,a14570,a14572,a14574,
a14576,a14578,a14580,a14582,a14584,a14586,a14588,a14590,a14592,a14594,a14596,a14598,a14600,a14602,a14604,
a14606,a14608,a14610,a14612,a14614,a14616,a14618,a14620,a14622,a14624,a14626,a14628,a14630,a14632,a14634,
a14636,a14638,a14640,a14642,a14644,a14646,a14648,a14650,a14652,a14654,a14656,a14658,a14660,a14662,a14664,
a14666,a14668,a14670,a14672,a14674,a14676,a14678,a14680,a14682,a14684,a14686,a14688,a14690,a14692,a14694,
a14696,a14698,a14700,a14702,a14704,a14706,a14708,a14710,a14712,a14714,a14716,a14718,a14720,a14722,a14724,
a14726,a14728,a14730,a14732,a14734,a14736,a14738,a14740,a14742,a14744,a14746,a14748,a14750,a14752,a14754,
a14756,a14758,a14760,a14762,a14764,a14766,a14768,a14770,a14772,a14774,a14776,a14778,a14780,a14782,a14784,
a14786,a14788,a14790,a14792,a14794,a14796,a14798,a14800,a14802,a14804,a14806,a14808,a14810,a14812,a14814,
a14816,a14818,a14820,a14822,a14824,a14826,a14828,a14830,a14832,a14834,a14836,a14838,a14840,a14842,a14844,
a14846,a14848,a14850,a14852,a14854,a14856,a14858,a14860,a14862,a14864,a14866,a14868,a14870,a14872,a14874,
a14876,a14878,a14880,a14882,a14884,a14886,a14888,a14890,a14892,a14894,a14896,a14898,a14900,a14902,a14904,
a14906,a14908,a14910,a14912,a14914,a14916,a14918,a14920,a14922,a14924,a14926,a14928,a14930,a14932,a14934,
a14936,a14938,a14940,a14942,a14944,a14946,a14948,a14950,a14952,a14954,a14956,a14958,a14960,a14962,a14964,
a14966,a14968,a14970,a14972,a14974,a14976,a14978,a14980,a14982,a14984,a14986,a14988,a14990,a14992,a14994,
a14996,a14998,a15000,a15002,a15004,a15006,a15008,a15010,a15012,a15014,a15016,a15018,a15020,a15022,a15024,
a15026,a15028,a15030,a15032,a15034,a15036,a15038,a15040,a15042,a15044,a15046,a15048,a15050,a15052,a15054,
a15056,a15058,a15060,a15062,a15064,a15066,a15068,a15070,a15072,a15074,a15076,a15078,a15080,a15082,a15084,
a15086,a15088,a15090,a15092,a15094,a15096,a15098,a15100,a15102,a15104,a15106,a15108,a15110,a15112,a15114,
a15116,a15118,a15120,a15122,a15124,a15126,a15128,a15130,a15132,a15134,a15136,a15138,a15140,a15142,a15144,
a15146,a15148,a15150,a15152,a15154,a15156,a15158,a15160,a15162,a15164,a15166,a15168,a15170,a15172,a15174,
a15176,a15178,a15180,a15182,a15184,a15186,a15188,a15190,a15192,a15194,a15196,a15198,a15200,a15202,a15204,
a15206,a15208,a15210,a15212,a15214,a15216,a15218,a15220,a15222,a15224,a15226,a15228,a15230,a15232,a15234,
a15236,a15238,a15240,a15242,a15244,a15246,a15248,a15250,a15252,a15254,a15256,a15258,a15260,a15262,a15264,
a15266,a15268,a15270,a15272,a15274,a15276,a15278,a15280,a15282,a15284,a15286,a15288,a15290,a15292,a15294,
a15296,a15298,a15300,a15302,a15304,a15306,a15308,a15310,a15312,a15314,a15316,a15318,a15320,a15322,a15324,
a15326,a15328,a15330,a15332,a15334,a15336,a15338,a15340,a15342,a15344,a15346,a15348,a15350,a15352,a15354,
a15356,a15358,a15360,a15362,a15364,a15366,a15368,a15370,a15372,a15374,a15376,a15378,a15380,a15382,a15384,
a15386,a15388,a15390,a15392,a15394,a15396,a15398,a15400,a15402,a15404,a15406,a15408,a15410,a15412,a15414,
a15416,a15418,a15420,a15422,a15424,a15426,a15428,a15430,a15432,a15434,a15436,a15438,a15440,a15442,a15444,
a15446,a15448,a15450,a15452,a15454,a15456,a15458,a15460,a15462,a15464,a15466,a15468,a15470,a15472,a15474,
a15476,a15478,a15480,a15482,a15484,a15486,a15488,a15490,a15492,a15494,a15496,a15498,a15500,a15502,a15504,
a15506,a15508,a15510,a15512,a15514,a15516,a15518,a15520,a15522,a15524,a15526,a15528,a15530,a15532,a15534,
a15536,a15538,a15540,a15542,a15544,a15546,a15548,a15550,a15552,a15554,a15556,a15558,a15560,a15562,a15564,
a15566,a15568,a15570,a15572,a15574,a15576,a15578,a15580,a15582,a15584,a15586,a15588,a15590,a15592,a15594,
a15596,a15598,a15600,a15602,a15604,a15606,a15608,a15610,a15612,a15614,a15616,a15618,a15620,a15622,a15624,
a15626,a15628,a15630,a15632,a15634,a15636,a15638,a15640,a15642,a15644,a15646,a15648,a15650,a15652,a15654,
a15656,a15658,a15660,a15662,a15664,a15666,a15668,a15670,a15672,a15674,a15676,a15678,a15680,a15682,a15684,
a15686,a15688,a15690,a15692,a15694,a15696,a15698,a15700,a15702,a15704,a15706,a15708,a15710,a15712,a15714,
a15716,a15718,a15720,a15722,a15724,a15726,a15728,a15730,a15732,a15734,a15736,a15738,a15740,a15742,a15744,
a15746,a15748,a15750,a15752,a15754,a15756,a15758,a15760,a15762,a15764,a15766,a15768,a15770,a15772,a15774,
a15776,a15778,a15780,a15782,a15784,a15786,a15788,a15790,a15792,a15794,a15796,a15798,a15800,a15802,a15804,
a15806,a15808,a15810,a15812,a15814,a15816,a15818,a15820,a15822,a15824,a15826,a15828,a15830,a15832,a15834,
a15836,a15838,a15840,a15842,a15844,a15846,a15848,a15850,a15852,a15854,a15856,a15858,a15860,a15862,a15864,
a15866,a15868,a15870,a15872,a15874,a15876,a15878,a15880,a15882,a15884,a15886,a15888,a15890,a15892,a15894,
a15896,a15898,a15900,a15902,a15904,a15906,a15908,a15910,a15912,a15914,a15916,a15918,a15920,a15922,a15924,
a15926,a15928,a15930,a15932,a15934,a15936,a15938,a15940,a15942,a15944,a15946,a15948,a15950,a15952,a15954,
a15956,a15958,a15960,a15962,a15964,a15966,a15968,a15970,a15972,a15974,a15976,a15978,a15980,a15982,a15984,
a15986,a15988,a15990,a15992,a15994,a15996,a15998,a16000,a16002,a16004,a16006,a16008,a16010,a16012,a16014,
a16016,a16018,a16020,a16022,a16024,a16026,a16028,a16030,a16032,a16034,a16036,a16038,a16040,a16042,a16044,
a16046,a16048,a16050,a16052,a16054,a16056,a16058,a16060,a16062,a16064,a16066,a16068,a16070,a16072,a16074,
a16076,a16078,a16080,a16082,a16084,a16086,a16088,a16090,a16092,a16094,a16096,a16098,a16100,a16102,a16104,
a16106,a16108,a16110,a16112,a16114,a16116,a16118,a16120,a16122,a16124,a16126,a16128,a16130,a16132,a16134,
a16136,a16138,a16140,a16142,a16144,a16146,a16148,a16150,a16152,a16154,a16156,a16158,a16160,a16162,a16164,
a16166,a16168,a16170,a16172,a16174,a16176,a16178,a16180,a16182,a16184,a16186,a16188,a16190,a16192,a16194,
a16196,a16198,a16200,a16202,a16204,a16206,a16208,a16210,a16212,a16214,a16216,a16218,a16220,a16222,a16224,
a16226,a16228,a16230,a16232,a16234,a16236,a16238,a16240,a16242,a16244,a16246,a16248,a16250,a16252,a16254,
a16256,a16258,a16260,a16262,a16264,a16266,a16268,a16270,a16272,a16274,a16276,a16278,a16280,a16282,a16284,
a16286,a16288,a16290,a16292,a16294,a16296,a16298,a16300,a16302,a16304,a16306,a16308,a16310,a16312,a16314,
a16316,a16318,a16320,a16322,a16324,a16326,a16328,a16330,a16332,a16334,a16336,a16338,a16340,a16342,a16344,
a16346,a16348,a16350,a16352,a16354,a16356,a16358,a16360,a16362,a16364,a16366,a16368,a16370,a16372,a16374,
a16376,a16378,a16380,a16382,a16384,a16386,a16388,a16390,a16392,a16394,a16396,a16398,a16400,a16402,a16404,
a16406,a16408,a16410,a16412,a16414,a16416,a16418,a16420,a16422,a16424,a16426,a16428,a16430,a16432,a16434,
a16436,a16438,a16440,a16442,a16444,a16446,a16448,a16450,a16452,a16454,a16456,a16458,a16460,a16462,a16464,
a16466,a16468,a16470,a16472,a16474,a16476,a16478,a16480,a16482,a16484,a16486,a16488,a16490,a16492,a16494,
a16496,a16498,a16500,a16502,a16504,a16506,a16508,a16510,a16512,a16514,a16516,a16518,a16520,a16522,a16524,
a16526,a16528,a16530,a16532,a16534,a16536,a16538,a16540,a16542,a16544,a16546,a16548,a16550,a16552,a16554,
a16556,a16558,a16560,a16562,a16564,a16566,a16568,a16570,a16572,a16574,a16576,a16578,a16580,a16582,a16584,
a16586,a16588,a16590,a16592,a16594,a16596,a16598,a16600,a16602,a16604,a16606,a16608,a16610,a16612,a16614,
a16616,a16618,a16620,a16622,a16624,a16626,a16628,a16630,a16632,a16634,a16636,a16638,a16640,a16642,a16644,
a16646,a16648,a16650,a16652,a16654,a16656,a16658,a16660,a16662,a16664,a16666,a16668,a16670,a16672,a16674,
a16676,a16678,a16680,a16682,a16684,a16686,a16688,a16690,a16692,a16694,a16696,a16698,a16700,a16702,a16704,
a16706,a16708,a16710,a16712,a16714,a16716,a16718,a16720,a16722,a16724,a16726,a16728,a16730,a16732,a16734,
a16736,a16738,a16740,a16742,a16744,a16746,a16748,a16750,a16752,a16754,a16756,a16758,a16760,a16762,a16764,
a16766,a16768,a16770,a16772,a16774,a16776,a16778,a16780,a16782,a16784,a16786,a16788,a16790,a16792,a16794,
a16796,a16798,a16800,a16802,a16804,a16806,a16808,a16810,a16812,a16814,a16816,a16818,a16820,a16822,a16824,
a16826,a16828,a16830,a16832,a16834,a16836,a16838,a16840,a16842,a16844,a16846,a16848,a16850,a16852,a16854,
a16856,a16858,a16860,a16862,a16864,a16866,a16868,a16870,a16872,a16874,a16876,a16878,a16880,a16882,a16884,
a16886,a16888,a16890,a16892,a16894,a16896,a16898,a16900,a16902,a16904,a16906,a16908,a16910,a16912,a16914,
a16916,a16918,a16920,a16922,a16924,a16926,a16928,a16930,a16932,a16934,a16936,a16938,a16940,a16942,a16944,
a16946,a16948,a16950,a16952,a16954,a16956,a16958,a16960,a16962,a16964,a16966,a16968,a16970,a16972,a16974,
a16976,a16978,a16980,a16982,a16984,a16986,a16988,a16990,a16992,a16994,a16996,a16998,a17000,a17002,a17004,
a17006,a17008,a17010,a17012,a17014,a17016,a17018,a17020,a17022,a17024,a17026,a17028,a17030,a17032,a17034,
a17036,a17038,a17040,a17042,a17044,a17046,a17048,a17050,a17052,a17054,a17056,a17058,a17060,a17062,a17064,
a17066,a17068,a17070,a17072,a17074,a17076,a17078,a17080,a17082,a17084,a17086,a17088,a17090,a17092,a17094,
a17096,a17098,a17100,a17102,a17104,a17106,a17108,a17110,a17112,a17114,a17116,a17118,a17120,a17122,a17124,
a17126,a17128,a17130,a17132,a17134,a17136,a17138,a17140,a17142,a17144,a17146,a17148,a17150,a17152,a17154,
a17156,a17158,a17160,a17162,a17164,a17166,a17168,a17170,a17172,a17174,a17176,a17178,a17180,a17182,a17184,
a17186,a17188,a17190,a17192,a17194,a17196,a17198,a17200,a17202,a17204,a17206,a17208,a17210,a17212,a17214,
a17216,a17218,a17220,a17222,a17224,a17226,a17228,a17230,a17232,a17234,a17236,a17238,a17240,a17242,a17244,
a17246,a17248,a17250,a17252,a17254,a17256,a17258,a17260,a17262,a17264,a17266,a17268,a17270,a17272,a17274,
a17276,a17278,a17280,a17282,a17284,a17286,a17288,a17290,a17292,a17294,a17296,a17298,a17300,a17302,a17304,
a17306,a17308,a17310,a17312,a17314,a17316,a17318,a17320,a17322,a17324,a17326,a17328,a17330,a17332,a17334,
a17336,a17338,a17340,a17342,a17344,a17346,a17348,a17350,a17352,a17354,a17356,a17358,a17360,a17362,a17364,
a17366,a17368,a17370,a17372,a17374,a17376,a17378,a17380,a17382,a17384,a17386,a17388,a17390,a17392,a17394,
a17396,a17398,a17400,a17402,a17404,a17406,a17408,a17410,a17412,a17414,a17416,a17418,a17420,a17422,a17424,
a17426,a17428,a17430,a17432,a17434,a17436,a17438,a17440,a17442,a17444,a17446,a17448,a17450,a17452,a17454,
a17456,a17458,a17460,a17462,a17464,a17466,a17468,a17470,a17472,a17474,a17476,a17478,a17480,a17482,a17484,
a17486,a17488,a17490,a17492,a17494,a17496,a17498,a17500,a17502,a17504,a17506,a17508,a17510,a17512,a17514,
a17516,a17518,a17520,a17522,a17524,a17526,a17528,a17530,a17532,a17534,a17536,a17538,a17540,a17542,a17544,
a17546,a17548,a17550,a17552,a17554,a17556,a17558,a17560,a17562,a17564,a17566,a17568,a17570,a17572,a17574,
a17576,a17578,a17580,a17582,a17584,a17586,a17588,a17590,a17592,a17594,a17596,a17598,a17600,a17602,a17604,
a17606,a17608,a17610,a17612,a17614,a17616,a17618,a17620,a17622,a17624,a17626,a17628,a17630,a17632,a17634,
a17636,a17638,a17640,a17642,a17644,a17646,a17648,a17650,a17652,a17654,a17656,a17658,a17660,a17662,a17664,
a17666,a17668,a17670,a17672,a17674,a17676,a17678,a17680,a17682,a17684,a17686,a17688,a17690,a17692,a17694,
a17696,a17698,a17700,a17702,a17704,a17706,a17708,a17710,a17712,a17714,a17716,a17718,a17720,a17722,a17724,
a17726,a17728,a17730,a17732,a17734,a17736,a17738,a17740,a17742,a17744,a17746,a17748,a17750,a17752,a17754,
a17756,a17758,a17760,a17762,a17764,a17766,a17768,a17770,a17772,a17774,a17776,a17778,a17780,a17782,a17784,
a17786,a17788,a17790,a17792,a17794,a17796,a17798,a17800,a17802,a17804,a17806,a17808,a17810,a17812,a17814,
a17816,a17818,a17820,a17822,a17824,a17826,a17828,a17830,a17832,a17834,a17836,a17838,a17840,a17842,a17844,
a17846,a17848,a17850,a17852,a17854,a17856,a17858,a17860,a17862,a17864,a17866,a17868,a17870,a17872,a17874,
a17876,a17878,a17880,a17882,a17884,a17886,a17888,a17890,a17892,a17894,a17896,a17898,a17900,a17902,a17904,
a17906,a17908,a17910,a17912,a17914,a17916,a17918,a17920,a17922,a17924,a17926,a17928,a17930,a17932,a17934,
a17936,a17938,a17940,a17942,a17944,a17946,a17948,a17950,a17952,a17954,a17956,a17958,a17960,a17962,a17964,
a17966,a17968,a17970,a17972,a17974,a17976,a17978,a17980,a17982,a17984,a17986,a17988,a17990,a17992,a17994,
a17996,a17998,a18000,a18002,a18004,a18006,a18008,a18010,a18012,a18014,a18016,a18018,a18020,a18022,a18024,
a18026,a18028,a18030,a18032,a18034,a18036,a18038,a18040,a18042,a18044,a18046,a18048,a18050,a18052,a18054,
a18056,a18058,a18060,a18062,a18064,a18066,a18068,a18070,a18072,a18074,a18076,a18078,a18080,a18082,a18084,
a18086,a18088,a18090,a18092,a18094,a18096,a18098,a18100,a18102,a18104,a18106,a18108,a18110,a18112,a18114,
a18116,a18118,a18120,a18122,a18124,a18126,a18128,a18130,a18132,a18134,a18136,a18138,a18140,a18142,a18144,
a18146,a18148,a18150,a18152,a18154,a18156,a18158,a18160,a18162,a18164,a18166,a18168,a18170,a18172,a18174,
a18176,a18178,a18180,a18182,a18184,a18186,a18188,a18190,a18192,a18194,a18196,a18198,a18200,a18202,a18204,
a18206,a18208,a18210,a18212,a18214,a18216,a18218,a18220,a18222,a18224,a18226,a18228,a18230,a18232,a18234,
a18236,a18238,a18240,a18242,a18244,a18246,a18248,a18250,a18252,a18254,a18256,a18258,a18260,a18262,a18264,
a18266,a18268,a18270,a18272,a18274,a18276,a18278,a18280,a18282,a18284,a18286,a18288,a18290,a18292,a18294,
a18296,a18298,a18300,a18302,a18304,a18306,a18308,a18310,a18312,a18314,a18316,a18318,a18320,a18322,a18324,
a18326,a18328,a18330,a18332,a18334,a18336,a18338,a18340,a18342,a18344,a18346,a18348,a18350,a18352,a18354,
a18356,a18358,a18360,a18362,a18364,a18366,a18368,a18370,a18372,a18374,a18376,a18378,a18380,a18382,a18384,
a18386,a18388,a18390,a18392,a18394,a18396,a18398,a18400,a18402,a18404,a18406,a18408,a18410,a18412,a18414,
a18416,a18418,a18420,a18422,a18424,a18426,a18428,a18430,a18432,a18434,a18436,a18438,a18440,a18442,a18444,
a18446,a18448,a18450,a18452,a18454,a18456,a18458,a18460,a18462,a18464,a18466,a18468,a18470,a18472,a18474,
a18476,a18478,a18480,a18482,a18484,a18486,a18488,a18490,a18492,a18494,a18496,a18498,a18500,a18502,a18504,
a18506,a18508,a18510,a18512,a18514,a18516,a18518,a18520,a18522,a18524,a18526,a18528,a18530,a18532,a18534,
a18536,a18538,a18540,a18542,a18544,a18546,a18548,a18550,a18552,a18554,a18556,a18558,a18560,a18562,a18564,
a18566,a18568,a18570,a18572,a18574,a18576,a18578,a18580,a18582,a18584,a18586,a18588,a18590,a18592,a18594,
a18596,a18598,a18600,a18602,a18604,a18606,a18608,a18610,a18612,a18614,a18616,a18618,a18620,a18622,a18624,
a18626,a18628,a18630,a18632,a18634,a18636,a18638,a18640,a18642,a18644,a18646,a18648,a18650,a18652,a18654,
a18656,a18658,a18660,a18662,a18664,a18666,a18668,a18670,a18672,a18674,a18676,a18678,a18680,a18682,a18684,
a18686,a18688,a18690,a18692,a18694,a18696,a18698,a18700,a18702,a18704,a18706,a18708,a18710,a18712,a18714,
a18716,a18718,a18720,a18722,a18724,a18726,a18728,a18730,a18732,a18734,a18736,a18738,a18740,a18742,a18744,
a18746,a18748,a18750,a18752,a18754,a18756,a18758,a18760,a18762,a18764,a18766,a18768,a18770,a18772,a18774,
a18776,a18778,a18780,a18782,a18784,a18786,a18788,a18790,a18792,a18794,a18796,a18798,a18800,a18802,a18804,
a18806,a18808,a18810,a18812,a18814,a18816,a18818,a18820,a18822,a18824,a18826,a18828,a18830,a18832,a18834,
a18836,a18838,a18840,a18842,a18844,a18846,a18848,a18850,a18852,a18854,a18856,a18858,a18860,a18862,a18864,
a18866,a18868,a18870,a18872,a18874,a18876,a18878,a18880,a18882,a18884,a18886,a18888,a18890,a18892,a18894,
a18896,a18898,a18900,a18902,a18904,a18906,a18908,a18910,a18912,a18914,a18916,a18918,a18920,a18922,a18924,
a18926,a18928,a18930,a18932,a18934,a18936,a18938,a18940,a18942,a18944,a18946,a18948,a18950,a18952,a18954,
a18956,a18958,a18960,a18962,a18964,a18966,a18968,a18970,a18972,a18974,a18976,a18978,a18980,a18982,a18984,
a18986,a18988,a18990,a18992,a18994,a18996,a18998,a19000,a19002,a19004,a19006,a19008,a19010,a19012,a19014,
a19016,a19018,a19020,a19022,a19024,a19026,a19028,a19030,a19032,a19034,a19036,a19038,a19040,a19042,a19044,
a19046,a19048,a19050,a19052,a19054,a19056,a19058,a19060,a19062,a19064,a19066,a19068,a19070,a19072,a19074,
a19076,a19078,a19080,a19082,a19084,a19086,a19088,a19090,a19092,a19094,a19096,a19098,a19100,a19102,a19104,
a19106,a19108,a19110,a19112,a19114,a19116,a19118,a19120,a19122,a19124,a19126,a19128,a19130,a19132,a19134,
a19136,a19138,a19140,a19142,a19144,a19146,a19148,a19150,a19152,a19154,a19156,a19158,a19160,a19162,a19164,
a19166,a19168,a19170,a19172,a19174,a19176,a19178,a19180,a19182,a19184,a19186,a19188,a19190,a19192,a19194,
a19196,a19198,a19200,a19202,a19204,a19206,a19208,a19210,a19212,a19214,a19216,a19218,a19220,a19222,a19224,
a19226,a19228,a19230,a19232,a19234,a19236,a19238,a19240,a19242,a19244,a19246,a19248,a19250,a19252,a19254,
a19256,a19258,a19260,a19262,a19264,a19266,a19268,a19270,a19272,a19274,a19276,a19278,a19280,a19282,a19284,
a19286,a19288,a19290,a19292,a19294,a19296,a19298,a19300,a19302,a19304,a19306,a19308,a19310,a19312,a19314,
a19316,a19318,a19320,a19322,a19324,a19326,a19328,a19330,a19332,a19334,a19336,a19338,a19340,a19342,a19344,
a19346,a19348,a19350,a19352,a19354,a19356,a19358,a19360,a19362,a19364,a19366,a19368,a19370,a19372,a19374,
a19376,a19378,a19380,a19382,a19384,a19386,a19388,a19390,a19392,a19394,a19396,a19398,a19400,a19402,a19404,
a19406,a19408,a19410,a19412,a19414,a19416,a19418,a19420,a19422,a19424,a19426,a19428,a19430,a19432,a19434,
a19436,a19438,a19440,a19442,a19444,a19446,a19448,a19450,a19452,a19454,a19456,a19458,a19460,a19462,a19464,
a19466,a19468,a19470,a19472,a19474,a19476,a19478,a19480,a19482,a19484,a19486,a19488,a19490,a19492,a19494,
a19496,a19498,a19500,a19502,a19504,a19506,a19508,a19510,a19512,a19514,a19516,a19518,a19520,a19522,a19524,
a19526,a19528,a19530,a19532,a19534,a19536,a19538,a19540,a19542,a19544,a19546,a19548,a19550,a19552,a19554,
a19556,a19558,a19560,a19562,a19564,a19566,a19568,a19570,a19572,a19574,a19576,a19578,a19580,a19582,a19584,
a19586,a19588,a19590,a19592,a19594,a19596,a19598,a19600,a19602,a19604,a19606,a19608,a19610,a19612,a19614,
a19616,a19618,a19620,a19622,a19624,a19626,a19628,a19630,a19632,a19634,a19636,a19638,a19640,a19642,a19644,
a19646,a19648,a19650,a19652,a19654,a19656,a19658,a19660,a19662,a19664,a19666,a19668,a19670,a19672,a19674,
a19676,a19678,a19680,a19682,a19684,a19686,a19688,a19690,a19692,a19694,a19696,a19698,a19700,a19702,a19704,
a19706,a19708,a19710,a19712,a19714,a19716,a19718,a19720,a19722,a19724,a19726,a19728,a19730,a19732,a19734,
a19736,a19738,a19740,a19742,a19744,a19746,a19748,a19750,a19752,a19754,a19756,a19758,a19760,a19762,a19764,
a19766,a19768,a19770,a19772,a19774,a19776,a19778,a19780,a19782,a19784,a19786,a19788,a19790,a19792,a19794,
a19796,a19798,a19800,a19802,a19804,a19806,a19808,a19810,a19812,a19814,a19816,a19818,a19820,a19822,a19824,
a19826,a19828,a19830,a19832,a19834,a19836,a19838,a19840,a19842,a19844,a19846,a19848,a19850,a19852,a19854,
a19856,a19858,a19860,a19862,a19864,a19866,a19868,a19870,a19872,a19874,a19876,a19878,a19880,a19882,a19884,
a19886,a19888,a19890,a19892,a19894,a19896,a19898,a19900,a19902,a19904,a19906,a19908,a19910,a19912,a19914,
a19916,a19918,a19920,a19922,a19924,a19926,a19928,a19930,a19932,a19934,a19936,a19938,a19940,a19942,a19944,
a19946,a19948,a19950,a19952,a19954,a19956,a19958,a19960,a19962,a19964,a19966,a19968,a19970,a19972,a19974,
a19976,a19978,a19980,a19982,a19984,a19986,a19988,a19990,a19992,a19994,a19996,a19998,a20000,a20002,a20004,
a20006,a20008,a20010,a20012,a20014,a20016,a20018,a20020,a20022,a20024,a20026,a20028,a20030,a20032,a20034,
a20036,a20038,a20040,a20042,a20044,a20046,a20048,a20050,a20052,a20054,a20056,a20058,a20060,a20062,a20064,
a20066,a20068,a20070,a20072,a20074,a20076,a20078,a20080,a20082,a20084,a20086,a20088,a20090,a20092,a20094,
a20096,a20098,a20100,a20102,a20104,a20106,a20108,a20110,a20112,a20114,a20116,a20118,a20120,a20122,a20124,
a20126,a20128,a20130,a20132,a20134,a20136,a20138,a20140,a20142,a20144,a20146,a20148,a20150,a20152,a20154,
a20156,a20158,a20160,a20162,a20164,a20166,a20168,a20170,a20172,a20174,a20176,a20178,a20180,a20182,a20184,
a20186,a20188,a20190,a20192,a20194,a20196,a20198,a20200,a20202,a20204,a20206,a20208,a20210,a20212,a20214,
a20216,a20218,a20220,a20222,a20224,a20226,a20228,a20230,a20232,a20234,a20236,a20238,a20240,a20242,a20244,
a20246,a20248,a20250,a20252,a20254,a20256,a20258,a20260,a20262,a20264,a20266,a20268,a20270,a20272,a20274,
a20276,a20278,a20280,a20282,a20284,a20286,a20288,a20290,a20292,a20294,a20296,a20298,a20300,a20302,a20304,
a20306,a20308,a20310,a20312,a20314,a20316,a20318,a20320,a20322,a20324,a20326,a20328,a20330,a20332,a20334,
a20336,a20338,a20340,a20342,a20344,a20346,a20348,a20350,a20352,a20354,a20356,a20358,a20360,a20362,a20364,
a20366,a20368,a20370,a20372,a20374,a20376,a20378,a20380,a20382,a20384,a20386,a20388,a20390,a20392,a20394,
a20396,a20398,a20400,a20402,a20404,a20406,a20408,a20410,a20412,a20414,a20416,a20418,a20420,a20422,a20424,
a20426,a20428,a20430,a20432,a20434,a20436,a20438,a20440,a20442,a20444,a20446,a20448,a20450,a20452,a20454,
a20456,a20458,a20460,a20462,a20464,a20466,a20468,a20470,a20472,a20474,a20476,a20478,a20480,a20482,a20484,
a20486,a20488,a20490,a20492,a20494,a20496,a20498,a20500,a20502,a20504,a20506,a20508,a20510,a20512,a20514,
a20516,a20518,a20520,a20522,a20524,a20526,a20528,a20530,a20532,a20534,a20536,a20538,a20540,a20542,a20544,
a20546,a20548,a20550,a20552,a20554,a20556,a20558,a20560,a20562,a20564,a20566,a20568,a20570,a20572,a20574,
a20576,a20578,a20580,a20582,a20584,a20586,a20588,a20590,a20592,a20594,a20596,a20598,a20600,a20602,a20604,
a20606,a20608,a20610,a20612,a20614,a20616,a20618,a20620,a20622,a20624,a20626,a20628,a20630,a20632,a20634,
a20636,a20638,a20640,a20642,a20644,a20646,a20648,a20650,a20652,a20654,a20656,a20658,a20660,a20662,a20664,
a20666,a20668,a20670,a20672,a20674,a20676,a20678,a20680,a20682,a20684,a20686,a20688,a20690,a20692,a20694,
a20696,a20698,a20700,a20702,a20704,a20706,a20708,a20710,a20712,a20714,a20716,a20718,a20720,a20722,a20724,
a20726,a20728,a20730,a20732,a20734,a20736,a20738,a20740,a20742,a20744,a20746,a20748,a20750,a20752,a20754,
a20756,a20758,a20760,a20762,a20764,a20766,a20768,a20770,a20772,a20774,a20776,a20778,a20780,a20782,a20784,
a20786,a20788,a20790,a20792,a20794,a20796,a20798,a20800,a20802,a20804,a20806,a20808,a20810,a20812,a20814,
a20816,a20818,a20820,a20822,a20824,a20826,a20828,a20830,a20832,a20834,a20836,a20838,a20840,a20842,a20844,
a20846,a20848,a20850,a20852,a20854,a20856,a20858,a20860,a20862,a20864,a20866,a20868,a20870,a20872,a20874,
a20876,a20878,a20880,a20882,a20884,a20886,a20888,a20890,a20892,a20894,a20896,a20898,a20900,a20902,a20904,
a20906,a20908,a20910,a20912,a20914,a20916,a20918,a20920,a20922,a20924,a20926,a20928,a20930,a20932,a20934,
a20936,a20938,a20940,a20942,a20944,a20946,a20948,a20950,a20952,a20954,a20956,a20958,a20960,a20962,a20964,
a20966,a20968,a20970,a20972,a20974,a20976,a20978,a20980,a20982,a20984,a20986,a20988,a20990,a20992,a20994,
a20996,a20998,a21000,a21002,a21004,a21006,a21008,a21010,a21012,a21014,a21016,a21018,a21020,a21022,a21024,
a21026,a21028,a21030,a21032,a21034,a21036,a21038,a21040,a21042,a21044,a21046,a21048,a21050,a21052,a21054,
a21056,a21058,a21060,a21062,a21064,a21066,a21068,a21070,a21072,a21074,a21076,a21078,a21080,a21082,a21084,
a21086,a21088,a21090,a21092,a21094,a21096,a21098,a21100,a21102,a21104,a21106,a21108,a21110,a21112,a21114,
a21116,a21118,a21120,a21122,a21124,a21126,a21128,a21130,a21132,a21134,a21136,a21138,a21140,a21142,a21144,
a21146,a21148,a21150,a21152,a21154,a21156,a21158,a21160,a21162,a21164,a21166,a21168,a21170,a21172,a21174,
a21176,a21178,a21180,a21182,a21184,a21186,a21188,a21190,a21192,a21194,a21196,a21198,a21200,a21202,a21204,
a21206,a21208,a21210,a21212,a21214,a21216,a21218,a21220,a21222,a21224,a21226,a21228,a21230,a21232,a21234,
a21236,a21238,a21240,a21242,a21244,a21246,a21248,a21250,a21252,a21254,a21256,a21258,a21260,a21262,a21264,
a21266,a21268,a21270,a21272,a21274,a21276,a21278,a21280,a21282,a21284,a21286,a21288,a21290,a21292,a21294,
a21296,a21298,a21300,a21302,a21304,a21306,a21308,a21310,a21312,a21314,a21316,a21318,a21320,a21322,a21324,
a21326,a21328,a21330,a21332,a21334,a21336,a21338,a21340,a21342,a21344,a21346,a21348,a21350,a21352,a21354,
a21356,a21358,a21360,a21362,a21364,a21366,a21368,a21370,a21372,a21374,a21376,a21378,a21380,a21382,a21384,
a21386,a21388,a21390,a21392,a21394,a21396,a21398,a21400,a21402,a21404,a21406,a21408,a21410,a21412,a21414,
a21416,a21418,a21420,a21422,a21424,a21426,a21428,a21430,a21432,a21434,a21436,a21438,a21440,a21442,a21444,
a21446,a21448,a21450,a21452,a21454,a21456,a21458,a21460,a21462,a21464,a21466,a21468,a21470,a21472,a21474,
a21476,a21478,a21480,a21482,a21484,a21486,a21488,a21490,a21492,a21494,a21496,a21498,a21500,a21502,a21504,
a21506,a21508,a21510,a21512,a21514,a21516,a21518,a21520,a21522,a21524,a21526,a21528,a21530,a21532,a21534,
a21536,a21538,a21540,a21542,a21544,a21546,a21548,a21550,a21552,a21554,a21556,a21558,a21560,a21562,a21564,
a21566,a21568,a21570,a21572,a21574,a21576,a21578,a21580,a21582,a21584,a21586,a21588,a21590,a21592,a21594,
a21596,a21598,a21600,a21602,a21604,a21606,a21608,a21610,a21612,a21614,a21616,a21618,a21620,a21622,a21624,
a21626,a21628,a21630,a21632,a21634,a21636,a21638,a21640,a21642,a21644,a21646,a21648,a21650,a21652,a21654,
a21656,a21658,a21660,a21662,a21664,a21666,a21668,a21670,a21672,a21674,a21676,a21678,a21680,a21682,a21684,
a21686,a21688,a21690,a21692,a21694,a21696,a21698,a21700,a21702,a21704,a21706,a21708,a21710,a21712,a21714,
a21716,a21718,a21720,a21722,a21724,a21726,a21728,a21730,a21732,a21734,a21736,a21738,a21740,a21742,a21744,
a21746,a21748,a21750,a21752,a21754,a21756,a21758,a21760,a21762,a21764,a21766,a21768,a21770,a21772,a21774,
a21776,a21778,a21780,a21782,a21784,a21786,a21788,a21790,a21792,a21794,a21796,a21798,a21800,a21802,a21804,
a21806,a21808,a21810,a21812,a21814,a21816,a21818,a21820,a21822,a21824,a21826,a21828,a21830,a21832,a21834,
a21836,a21838,a21840,a21842,a21844,a21846,a21848,a21850,a21852,a21854,a21856,a21858,a21860,a21862,a21864,
a21866,a21868,a21870,a21872,a21874,a21876,a21878,a21880,a21882,a21884,a21886,a21888,a21890,a21892,a21894,
a21896,a21898,a21900,a21902,a21904,a21906,a21908,a21910,a21912,a21914,a21916,a21918,a21920,a21922,a21924,
a21926,a21928,a21930,a21932,a21934,a21936,a21938,a21940,a21942,a21944,a21946,a21948,a21950,a21952,a21954,
a21956,a21958,a21960,a21962,a21964,a21966,a21968,a21970,a21972,a21974,a21976,a21978,a21980,a21982,a21984,
a21986,a21988,a21990,a21992,a21994,a21996,a21998,a22000,a22002,a22004,a22006,a22008,a22010,a22012,a22014,
a22016,a22018,a22020,a22022,a22024,a22026,a22028,a22030,a22032,a22034,a22036,a22038,a22040,a22042,a22044,
a22046,a22048,a22050,a22052,a22054,a22056,a22058,a22060,a22062,a22064,a22066,a22068,a22070,a22072,a22074,
a22076,a22078,a22080,a22082,a22084,a22086,a22088,a22090,a22092,a22094,a22096,a22098,a22100,a22102,a22104,
a22106,a22108,a22110,a22112,a22114,a22116,a22118,a22120,a22122,a22124,a22126,a22128,a22130,a22132,a22134,
a22136,a22138,a22140,a22142,a22144,a22146,a22148,a22150,a22152,a22154,a22156,a22158,a22160,a22162,a22164,
a22166,a22168,a22170,a22172,a22174,a22176,a22178,a22180,a22182,a22184,a22186,a22188,a22190,a22192,a22194,
a22196,a22198,a22200,a22202,a22204,a22206,a22208,a22210,a22212,a22214,a22216,a22218,a22220,a22222,a22224,
a22226,a22228,a22230,a22232,a22234,a22236,a22238,a22240,a22242,a22244,a22246,a22248,a22250,a22252,a22254,
a22256,a22258,a22260,a22262,a22264,a22266,a22268,a22270,a22272,a22274,a22276,a22278,a22280,a22282,a22284,
a22286,a22288,a22290,a22292,a22294,a22296,a22298,a22300,a22302,a22304,a22306,a22308,a22310,a22312,a22314,
a22316,a22318,a22320,a22322,a22324,a22326,a22328,a22330,a22332,a22334,a22336,a22338,a22340,a22342,a22344,
a22346,a22348,a22350,a22352,a22354,a22356,a22358,a22360,a22362,a22364,a22366,a22368,a22370,a22372,a22374,
a22376,a22378,a22380,a22382,a22384,a22386,a22388,a22390,a22392,a22394,a22396,a22398,a22400,a22402,a22404,
a22406,a22408,a22410,a22412,a22414,a22416,a22418,a22420,a22422,a22424,a22426,a22428,a22430,a22432,a22434,
a22436,a22438,a22440,a22442,a22444,a22446,a22448,a22450,a22452,a22454,a22456,a22458,a22460,a22462,a22464,
a22466,a22468,a22470,a22472,a22474,a22476,a22478,a22480,a22482,a22484,a22486,a22488,a22490,a22492,a22494,
a22496,a22498,a22500,a22502,a22504,a22506,a22508,a22510,a22512,a22514,a22516,a22518,a22520,a22522,a22524,
a22526,a22528,a22530,a22532,a22534,a22536,a22538,a22540,a22542,a22544,a22546,a22548,a22550,a22552,a22554,
a22556,a22558,a22560,a22562,a22564,a22566,a22568,a22570,a22572,a22574,a22576,a22578,a22580,a22582,a22584,
a22586,a22588,a22590,a22592,a22594,a22596,a22598,a22600,a22602,a22604,a22606,a22608,a22610,a22612,a22614,
a22616,a22618,a22620,a22622,a22624,a22626,a22628,a22630,a22632,a22634,a22636,a22638,a22640,a22642,a22644,
a22646,a22648,a22650,a22652,a22654,a22656,a22658,a22660,a22662,a22664,a22666,a22668,a22670,a22672,a22674,
a22676,a22678,a22680,a22682,a22684,a22686,a22688,a22690,a22692,a22694,a22696,a22698,a22700,a22702,a22704,
a22706,a22708,a22710,a22712,a22714,a22716,a22718,a22720,a22722,a22724,a22726,a22728,a22730,a22732,a22734,
a22736,a22738,a22740,a22742,a22744,a22746,a22748,a22750,a22752,a22754,a22756,a22758,a22760,a22762,a22764,
a22766,a22768,a22770,a22772,a22774,a22776,a22778,a22780,a22782,a22784,a22786,a22788,a22790,a22792,a22794,
a22796,a22798,a22800,a22802,a22804,a22806,a22808,a22810,a22812,a22814,a22816,a22818,a22820,a22822,a22824,
a22826,a22828,a22830,a22832,a22834,a22836,a22838,a22840,a22842,a22844,a22846,a22848,a22850,a22852,a22854,
a22856,a22858,a22860,a22862,a22864,a22866,a22868,a22870,a22872,a22874,a22876,a22878,a22880,a22882,a22884,
a22886,a22888,a22890,a22892,a22894,a22896,a22898,a22900,a22902,a22904,a22906,a22908,a22910,a22912,a22914,
a22916,a22918,a22920,a22922,a22924,a22926,a22928,a22930,a22932,a22934,a22936,a22938,a22940,a22942,a22944,
a22946,a22948,a22950,a22952,a22954,a22956,a22958,a22960,a22962,a22964,a22966,a22968,a22970,a22972,a22974,
a22976,a22978,a22980,a22982,a22984,a22986,a22988,a22990,a22992,a22994,a22996,a22998,a23000,a23002,a23004,
a23006,a23008,a23010,a23012,a23014,a23016,a23018,a23020,a23022,a23024,a23026,a23028,a23030,a23032,a23034,
a23036,a23038,a23040,a23042,a23044,a23046,a23048,a23050,a23052,a23054,a23056,a23058,a23060,a23062,a23064,
a23066,a23068,a23070,a23072,a23074,a23076,a23078,a23080,a23082,a23084,a23086,a23088,a23090,a23092,a23094,
a23096,a23098,a23100,a23102,a23104,a23106,a23108,a23110,a23112,a23114,a23116,a23118,a23120,a23122,a23124,
a23126,a23128,a23130,a23132,a23134,a23136,a23138,a23140,a23142,a23144,a23146,a23148,a23150,a23152,a23154,
a23156,a23158,a23160,a23162,a23164,a23166,a23168,a23170,a23172,a23174,a23176,a23178,a23180,a23182,a23184,
a23186,a23188,a23190,a23192,a23194,a23196,a23198,a23200,a23202,a23204,a23206,a23208,a23210,a23212,a23214,
a23216,a23218,a23220,a23222,a23224,a23226,a23228,a23230,a23232,a23234,a23236,a23238,a23240,a23242,a23244,
a23246,a23248,a23250,a23252,a23254,a23256,a23258,a23260,a23262,a23264,a23266,a23268,a23270,a23272,a23274,
a23276,a23278,a23280,a23282,a23284,a23286,a23288,a23290,a23292,a23294,a23296,a23298,a23300,a23302,a23304,
a23306,a23308,a23310,a23312,a23314,a23316,a23318,a23320,a23322,a23324,a23326,a23328,a23330,a23332,a23334,
a23336,a23338,a23340,a23342,a23344,a23346,a23348,a23350,a23352,a23354,a23356,a23358,a23360,a23362,a23364,
a23366,a23368,a23370,a23372,a23374,a23376,a23378,a23380,a23382,a23384,a23386,a23388,a23390,a23392,a23394,
a23396,a23398,a23400,a23402,a23404,a23406,a23408,a23410,a23412,a23414,a23416,a23418,a23420,a23422,a23424,
a23426,a23428,a23430,a23432,a23434,a23436,a23438,a23440,a23442,a23444,a23446,a23448,a23450,a23452,a23454,
a23456,a23458,a23460,a23462,a23464,a23466,a23468,a23470,a23472,a23474,a23476,a23478,a23480,a23482,a23484,
a23486,a23488,a23490,a23492,a23494,a23496,a23498,a23500,a23502,a23504,a23506,a23508,a23510,a23512,a23514,
a23516,a23518,a23520,a23522,a23524,a23526,a23528,a23530,a23532,a23534,a23536,a23538,a23540,a23542,a23544,
a23546,a23548,a23550,a23552,a23554,a23556,a23558,a23560,a23562,a23564,a23566,a23568,a23570,a23572,a23574,
a23576,a23578,a23580,a23582,a23584,a23586,a23588,a23590,a23592,a23594,a23596,a23598,a23600,a23602,a23604,
a23606,a23608,a23610,a23612,a23614,a23616,a23618,a23620,a23622,a23624,a23626,a23628,a23630,a23632,a23634,
a23636,a23638,a23640,a23642,a23644,a23646,a23648,a23650,a23652,a23654,a23656,a23658,a23660,a23662,a23664,
a23666,a23668,a23670,a23672,a23674,a23676,a23678,a23680,a23682,a23684,a23686,a23688,a23690,a23692,a23694,
a23696,a23698,a23700,a23702,a23704,a23706,a23708,a23710,a23712,a23714,a23716,a23718,a23720,a23722,a23724,
a23726,a23728,a23730,a23732,a23734,a23736,a23738,a23740,a23742,a23744,a23746,a23748,a23750,a23752,a23754,
a23756,a23758,a23760,a23762,a23764,a23766,a23768,a23770,a23772,a23774,a23776,a23778,a23780,a23782,a23784,
a23786,a23788,a23790,a23792,a23794,a23796,a23798,a23800,a23802,a23804,a23806,a23808,a23810,a23812,a23814,
a23816,a23818,a23820,a23822,a23824,a23826,a23828,a23830,a23832,a23834,a23836,a23838,a23840,a23842,a23844,
a23846,a23848,a23850,a23852,a23854,a23856,a23858,a23860,a23862,a23864,a23866,a23868,a23870,a23872,a23874,
a23876,a23878,a23880,a23882,a23884,a23886,a23888,a23890,a23892,a23894,a23896,a23898,a23900,a23902,a23904,
a23906,a23908,a23910,a23912,a23914,a23916,a23918,a23920,a23922,a23924,a23926,a23928,a23930,a23932,a23934,
a23936,a23938,a23940,a23942,a23944,a23946,a23948,a23950,a23952,a23954,a23956,a23958,a23960,a23962,a23964,
a23966,a23968,a23970,a23972,a23974,a23976,a23978,a23980,a23982,a23984,a23986,a23988,a23990,a23992,a23994,
a23996,a23998,a24000,a24002,a24004,a24006,a24008,a24010,a24012,a24014,a24016,a24018,a24020,a24022,a24024,
a24026,a24028,a24030,a24032,a24034,a24036,a24038,a24040,a24042,a24044,a24046,a24048,a24050,a24052,a24054,
a24056,a24058,a24060,a24062,a24064,a24066,a24068,a24070,a24072,a24074,a24076,a24078,a24080,a24082,a24084,
a24086,a24088,a24090,a24092,a24094,a24096,a24098,a24100,a24102,a24104,a24106,a24108,a24110,a24112,a24114,
a24116,a24118,a24120,a24122,a24124,a24126,a24128,a24130,a24132,a24134,a24136,a24138,a24140,a24142,a24144,
a24146,a24148,a24150,a24152,a24154,a24156,a24158,a24160,a24162,a24164,a24166,a24168,a24170,a24172,a24174,
a24176,a24178,a24180,a24182,a24184,a24186,a24188,a24190,a24192,a24194,a24196,a24198,a24200,a24202,a24204,
a24206,a24208,a24210,a24212,a24214,a24216,a24218,a24220,a24222,a24224,a24226,a24228,a24230,a24232,a24234,
a24236,a24238,a24240,a24242,a24244,a24246,a24248,a24250,a24252,a24254,a24256,a24258,a24260,a24262,a24264,
a24266,a24268,a24270,a24272,a24274,a24276,a24278,a24280,a24282,a24284,a24286,a24288,a24290,a24292,a24294,
a24296,a24298,a24300,a24302,a24304,a24306,a24308,a24310,a24312,a24314,a24316,a24318,a24320,a24322,a24324,
a24326,a24328,a24330,a24332,a24334,a24336,a24338,a24340,a24342,a24344,a24346,a24348,a24350,a24352,a24354,
a24356,a24358,a24360,a24362,a24364,a24366,a24368,a24370,a24372,a24374,a24376,a24378,a24380,a24382,a24384,
a24386,a24388,a24390,a24392,a24394,a24396,a24398,a24400,a24402,a24404,a24406,a24408,a24410,a24412,a24414,
a24416,a24418,a24420,a24422,a24424,a24426,a24428,a24430,a24432,a24434,a24436,a24438,a24440,a24442,a24444,
a24446,a24448,a24450,a24452,a24454,a24456,a24458,a24460,a24462,a24464,a24466,a24468,a24470,a24472,a24474,
a24476,a24478,a24480,a24482,a24484,a24486,a24488,a24490,a24492,a24494,a24496,a24498,a24500,a24502,a24504,
a24506,a24508,a24510,a24512,a24514,a24516,a24518,a24520,a24522,a24524,a24526,a24528,a24530,a24532,a24534,
a24536,a24538,a24540,a24542,a24544,a24546,a24548,a24550,a24552,a24554,a24556,a24558,a24560,a24562,a24564,
a24566,a24568,a24570,a24572,a24574,a24576,a24578,a24580,a24582,a24584,a24586,a24588,a24590,a24592,a24594,
a24596,a24598,a24600,a24602,a24604,a24606,a24608,a24610,a24612,a24614,a24616,a24618,a24620,a24622,a24624,
a24626,a24628,a24630,a24632,a24634,a24636,a24638,a24640,a24642,a24644,a24646,a24648,a24650,a24652,a24654,
a24656,a24658,a24660,a24662,a24664,a24666,a24668,a24670,a24672,a24674,a24676,a24678,a24680,a24682,a24684,
a24686,a24688,a24690,a24692,a24694,a24696,a24698,a24700,a24702,a24704,a24706,a24708,a24710,a24712,a24714,
a24716,a24718,a24720,a24722,a24724,a24726,a24728,a24730,a24732,a24734,a24736,a24738,a24740,a24742,a24744,
a24746,a24748,a24750,a24752,a24754,a24756,a24758,a24760,a24762,a24764,a24766,a24768,a24770,a24772,a24774,
a24776,a24778,a24780,a24782,a24784,a24786,a24788,a24790,a24792,a24794,a24796,a24798,a24800,a24802,a24804,
a24806,a24808,a24810,a24812,a24814,a24816,a24818,a24820,a24822,a24824,a24826,a24828,a24830,a24832,a24834,
a24836,a24838,a24840,a24842,a24844,a24846,a24848,a24850,a24852,a24854,a24856,a24858,a24860,a24862,a24864,
a24866,a24868,a24870,a24872,a24874,a24876,a24878,a24880,a24882,a24884,a24886,a24888,a24890,a24892,a24894,
a24896,a24898,a24900,a24902,a24904,a24906,a24908,a24910,a24912,a24914,a24916,a24918,a24920,a24922,a24924,
a24926,a24928,a24930,a24932,a24934,a24936,a24938,a24940,a24942,a24944,a24946,a24948,a24950,a24952,a24954,
a24956,a24958,a24960,a24962,a24964,a24966,a24968,a24970,a24972,a24974,a24976,a24978,a24980,a24982,a24984,
a24986,a24988,a24990,a24992,a24994,a24996,a24998,a25000,a25002,a25004,a25006,a25008,a25010,a25012,a25014,
a25016,a25018,a25020,a25022,a25024,a25026,a25028,a25030,a25032,a25034,a25036,a25038,a25040,a25042,a25044,
a25046,a25048,a25050,a25052,a25054,a25056,a25058,a25060,a25062,a25064,a25066,a25068,a25070,a25072,a25074,
a25076,a25078,a25080,a25082,a25084,a25086,a25088,a25090,a25092,a25094,a25096,a25098,a25100,a25102,a25104,
a25106,a25108,a25110,a25112,a25114,a25116,a25118,a25120,a25122,a25124,a25126,a25128,a25130,a25132,a25134,
a25136,a25138,a25140,a25142,a25144,a25146,a25148,a25150,a25152,a25154,a25156,a25158,a25160,a25162,a25164,
a25166,a25168,a25170,a25172,a25174,a25176,a25178,a25180,a25182,a25184,a25186,a25188,a25190,a25192,a25194,
a25196,a25198,a25200,a25202,a25204,a25206,a25208,a25210,a25212,a25214,a25216,a25218,a25220,a25222,a25224,
a25226,a25228,a25230,a25232,a25234,a25236,a25238,a25240,a25242,a25244,a25246,a25248,a25250,a25252,a25254,
a25256,a25258,a25260,a25262,a25264,a25266,a25268,a25270,a25272,a25274,a25276,a25278,a25280,a25282,a25284,
a25286,a25288,a25290,a25292,a25294,a25296,a25298,a25300,a25302,a25304,a25306,a25308,a25310,a25312,a25314,
a25316,a25318,a25320,a25322,a25324,a25326,a25328,a25330,a25332,a25334,a25336,a25338,a25340,a25342,a25344,
a25346,a25348,a25350,a25352,a25354,a25356,a25358,a25360,a25362,a25364,a25366,a25368,a25370,a25372,a25374,
a25376,a25378,a25380,a25382,a25384,a25386,a25388,a25390,a25392,a25394,a25396,a25398,a25400,a25402,a25404,
a25406,a25408,a25410,a25412,a25414,a25416,a25418,a25420,a25422,a25424,a25426,a25428,a25430,a25432,a25434,
a25436,a25438,a25440,a25442,a25444,a25446,a25448,a25450,a25452,a25454,a25456,a25458,a25460,a25462,a25464,
a25466,a25468,a25470,a25472,a25474,a25476,a25478,a25480,a25482,a25484,a25486,a25488,a25490,a25492,a25494,
a25496,a25498,a25500,a25502,a25504,a25506,a25508,a25510,a25512,a25514,a25516,a25518,a25520,a25522,a25524,
a25526,a25528,a25530,a25532,a25534,a25536,a25538,a25540,a25542,a25544,a25546,a25548,a25550,a25552,a25554,
a25556,a25558,a25560,a25562,a25564,a25566,a25568,a25570,a25572,a25574,a25576,a25578,a25580,a25582,a25584,
a25586,a25588,a25590,a25592,a25594,a25596,a25598,a25600,a25602,a25604,a25606,a25608,a25610,a25612,a25614,
a25616,a25618,a25620,a25622,a25624,a25626,a25628,a25630,a25632,a25634,a25636,a25638,a25640,a25642,a25644,
a25646,a25648,a25650,a25652,a25654,a25656,a25658,a25660,a25662,a25664,a25666,a25668,a25670,a25672,a25674,
a25676,a25678,a25680,a25682,a25684,a25686,a25688,a25690,a25692,a25694,a25696,a25698,a25700,a25702,a25704,
a25706,a25708,a25710,a25712,a25714,a25716,a25718,a25720,a25722,a25724,a25726,a25728,a25730,a25732,a25734,
a25736,a25738,a25740,a25742,a25744,a25746,a25748,a25750,a25752,a25754,a25756,a25758,a25760,a25762,a25764,
a25766,a25768,a25770,a25772,a25774,a25776,a25778,a25780,a25782,a25784,a25786,a25788,a25790,a25792,a25794,
a25796,a25798,a25800,a25802,a25804,a25806,a25808,a25810,a25812,a25814,a25816,a25818,a25820,a25822,a25824,
a25826,a25828,a25830,a25832,a25834,a25836,a25838,a25840,a25842,a25844,a25846,a25848,a25850,a25852,a25854,
a25856,a25858,a25860,a25862,a25864,a25866,a25868,a25870,a25872,a25874,a25876,a25878,a25880,a25882,a25884,
a25886,a25888,a25890,a25892,a25894,a25896,a25898,a25900,a25902,a25904,a25906,a25908,a25910,a25912,a25914,
a25916,a25918,a25920,a25922,a25924,a25926,a25928,a25930,a25932,a25934,a25936,a25938,a25940,a25942,a25944,
a25946,a25948,a25950,a25952,a25954,a25956,a25958,a25960,a25962,a25964,a25966,a25968,a25970,a25972,a25974,
a25976,a25978,a25980,a25982,a25984,a25986,a25988,a25990,a25992,a25994,a25996,a25998,a26000,a26002,a26004,
a26006,a26008,a26010,a26012,a26014,a26016,a26018,a26020,a26022,a26024,a26026,a26028,a26030,a26032,a26034,
a26036,a26038,a26040,a26042,a26044,a26046,a26048,a26050,a26052,a26054,a26056,a26058,a26060,a26062,a26064,
a26066,a26068,a26070,a26072,a26074,a26076,a26078,a26080,a26082,a26084,a26086,a26088,a26090,a26092,a26094,
a26096,a26098,a26100,a26102,a26104,a26106,a26108,a26110,a26112,a26114,a26116,a26118,a26120,a26122,a26124,
a26126,a26128,a26130,a26132,a26134,a26136,a26138,a26140,a26142,a26144,a26146,a26148,a26150,a26152,a26154,
a26156,a26158,a26160,a26162,a26164,a26166,a26168,a26170,a26172,a26174,a26176,a26178,a26180,a26182,a26184,
a26186,a26188,a26190,a26192,a26194,a26196,a26198,a26200,a26202,a26204,a26206,a26208,a26210,a26212,a26214,
a26216,a26218,a26220,a26222,a26224,a26226,a26228,a26230,a26232,a26234,a26236,a26238,a26240,a26242,a26244,
a26246,a26248,a26250,a26252,a26254,a26256,a26258,a26260,a26262,a26264,a26266,a26268,a26270,a26272,a26274,
a26276,a26278,a26280,a26282,a26284,a26286,a26288,a26290,a26292,a26294,a26296,a26298,a26300,a26302,a26304,
a26306,a26308,a26310,a26312,a26314,a26316,a26318,a26320,a26322,a26324,a26326,a26328,a26330,a26332,a26334,
a26336,a26338,a26340,a26342,a26344,a26346,a26348,a26350,a26352,a26354,a26356,a26358,a26360,a26362,a26364,
a26366,a26368,a26370,a26372,a26374,a26376,a26378,a26380,a26382,a26384,a26386,a26388,a26390,a26392,a26394,
a26396,a26398,a26400,a26402,a26404,a26406,a26408,a26410,a26412,a26414,a26416,a26418,a26420,a26422,a26424,
a26426,a26428,a26430,a26432,a26434,a26436,a26438,a26440,a26442,a26444,a26446,a26448,a26450,a26452,a26454,
a26456,a26458,a26460,a26462,a26464,a26466,a26468,a26470,a26472,a26474,a26476,a26478,a26480,a26482,a26484,
a26486,a26488,a26490,a26492,a26494,a26496,a26498,a26500,a26502,a26504,a26506,a26508,a26510,a26512,a26514,
a26516,a26518,a26520,a26522,a26524,a26526,a26528,a26530,a26532,a26534,a26536,a26538,a26540,a26542,a26544,
a26546,a26548,a26550,a26552,a26554,a26556,a26558,a26560,a26562,a26564,a26566,a26568,a26570,a26572,a26574,
a26576,a26578,a26580,a26582,a26584,a26586,a26588,a26590,a26592,a26594,a26596,a26598,a26600,a26602,a26604,
a26606,a26608,a26610,a26612,a26614,a26616,a26618,a26620,a26622,a26624,a26626,a26628,a26630,a26632,a26634,
a26636,a26638,a26640,a26642,a26644,a26646,a26648,a26650,a26652,a26654,a26656,a26658,a26660,a26662,a26664,
a26666,a26668,a26670,a26672,a26674,a26676,a26678,a26680,a26682,a26684,a26686,a26688,a26690,a26692,a26694,
a26696,a26698,a26700,a26702,a26704,a26706,a26708,a26710,a26712,a26714,a26716,a26718,a26720,a26722,a26724,
a26726,a26728,a26730,a26732,a26734,a26736,a26738,a26740,a26742,a26744,a26746,a26748,a26750,a26752,a26754,
a26756,a26758,a26760,a26762,a26764,a26766,a26768,a26770,a26772,a26774,a26776,a26778,a26780,a26782,a26784,
a26786,a26788,a26790,a26792,a26794,a26796,a26798,a26800,a26804,p0;

reg l730,l732,l734,l736,l738,l740,l742,l744,l746,l748,l750,l752,l754,l756,l758,
l760,l762,l764,l766,l768,l770,l772,l774,l776,l778,l780,l782,l784,l786,l788,
l790,l792,l794,l796,l798,l800,l802,l804,l806,l808,l810,l812,l814,l816,l818,
l820,l822,l824,l826,l828,l830,l832,l834,l836,l838,l840,l842,l844,l846,l848,
l850,l852,l854,l856,l858,l860,l862,l864,l866,l868,l870,l872,l874,l876,l878,
l880,l882,l884,l886,l888,l890,l892,l894,l896,l898,l900,l902,l904,l906,l908,
l910,l912,l914,l916,l918,l920,l922,l924,l926,l928,l930,l932,l934,l936,l938,
l940,l942,l944,l946,l948,l950,l952,l954,l956,l958,l960,l962,l964,l966,l968,
l970,l972,l974,l976,l978,l980,l982,l984,l986,l988,l990,l992,l994,l996,l998,
l1000,l1002,l1004,l1006,l1008,l1010,l1012,l1014,l1016,l1018,l1020,l1022,l1024,l1026,l1028,
l1030,l1032,l1034,l1036,l1038,l1040,l1042,l1044,l1046,l1048,l1050,l1052,l1054,l1056,l1058,
l1060,l1062,l1064,l1066,l1068,l1070,l1072,l1074,l1076,l1078,l1080,l1082,l1084,l1086,l1088,
l1090,l1092,l1094,l1096,l1098,l1100,l1102,l1104,l1106,l1108,l1110,l1112,l1114,l1116,l1118,
l1120,l1122,l1124,l1126,l1128,l1130,l1132,l1134,l1136,l1138,l1140,l1142,l1144,l1146,l1148,
l1150,l1152,l1154,l1156,l1158,l1160,l1162,l1164,l1166,l1168,l1170,l1172,l1174,l1176,l1178,
l1180,l1182,l1184,l1186,l1188,l1190,l1192,l1194,l1196,l1198,l1200,l1202,l1204,l1206,l1208,
l1210,l1212,l1214,l1216,l1218,l1220,l1222,l1224,l1226,l1228,l1230,l1232,l1234,l1236,l1238,
l1240,l1242,l1244,l1246,l1248,l1250,l1252,l1254,l1256,l1258,l1260,l1262,l1264,l1266,l1268,
l1270,l1272,l1274,l1276,l1278,l1280,l1282,l1284,l1286,l1288,l1290,l1292,l1294,l1296,l1298,
l1300,l1302,l1304,l1306,l1308,l1310,l1312,l1314,l1316,l1318,l1320,l1322,l1324,l1326,l1328,
l1330,l1332,l1334,l1336,l1338,l1340,l1342,l1344,l1346,l1348,l1350,l1352,l1354,l1356,l1358,
l1360,l1362,l1364,l1366,l1368,l1370,l1372,l1374,l1376,l1378,l1380,l1382,l1384,l1386,l1388,
l1390,l1392,l1394,l1396,l1398,l1400,l1402,l1404,l1406,l1408,l1410,l1412,l1414,l1416,l1418,
l1420,l1422,l1424,l1426,l1428,l1430,l1432,l1434,l1436,l1438,l1440,l1442,l1444,l1446,l1448,
l1450,l1452,l1454,l1456,l1458,l1460,l1462,l1464,l1466,l1468,l1470,l1472,l1474,l1476,l1478,
l1480,l1482,l1484,l1486,l1488,l1490,l1492,l1494,l1496,l1498,l1500,l1502,l1504,l1506,l1508,
l1510,l1512,l1514,l1516,l1518,l1520,l1522,l1524,l1526,l1528,l1530,l1532,l1534,l1536,l1538,
l1540,l1542,l1544,l1546,l1548,l1550,l1552,l1554,l1556,l1558,l1560,l1562,l1564,l1566,l1568,
l1570,l1572,l1574,l1576,l1578,l1580,l1582,l1584,l1586,l1588,l1590,l1592,l1594,l1596,l1598,
l1600,l1602,l1604,l1606,l1608,l1610,l1612,l1614,l1616,l1618,l1620,l1622,l1624,l1626,l1628,
l1630,l1632,l1634,l1636,l1638,l1640,l1642,l1644,l1646,l1648,l1650,l1652,l1654,l1656,l1658,
l1660,l1662,l1664,l1666,l1668,l1670,l1672,l1674,l1676,l1678;

initial
begin
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
   l802 = 0;
   l804 = 0;
   l806 = 0;
   l808 = 0;
   l810 = 0;
   l812 = 0;
   l814 = 0;
   l816 = 0;
   l818 = 0;
   l820 = 0;
   l822 = 0;
   l824 = 0;
   l826 = 0;
   l828 = 0;
   l830 = 0;
   l832 = 0;
   l834 = 0;
   l836 = 0;
   l838 = 0;
   l840 = 0;
   l842 = 0;
   l844 = 0;
   l846 = 0;
   l848 = 0;
   l850 = 0;
   l852 = 0;
   l854 = 0;
   l856 = 0;
   l858 = 0;
   l860 = 0;
   l862 = 0;
   l864 = 0;
   l866 = 0;
   l868 = 0;
   l870 = 0;
   l872 = 0;
   l874 = 0;
   l876 = 0;
   l878 = 0;
   l880 = 0;
   l882 = 0;
   l884 = 0;
   l886 = 0;
   l888 = 0;
   l890 = 0;
   l892 = 0;
   l894 = 0;
   l896 = 0;
   l898 = 0;
   l900 = 0;
   l902 = 0;
   l904 = 0;
   l906 = 0;
   l908 = 0;
   l910 = 0;
   l912 = 0;
   l914 = 0;
   l916 = 0;
   l918 = 0;
   l920 = 0;
   l922 = 0;
   l924 = 0;
   l926 = 0;
   l928 = 0;
   l930 = 0;
   l932 = 0;
   l934 = 0;
   l936 = 0;
   l938 = 0;
   l940 = 0;
   l942 = 0;
   l944 = 0;
   l946 = 0;
   l948 = 0;
   l950 = 0;
   l952 = 0;
   l954 = 0;
   l956 = 0;
   l958 = 0;
   l960 = 0;
   l962 = 0;
   l964 = 0;
   l966 = 0;
   l968 = 0;
   l970 = 0;
   l972 = 0;
   l974 = 0;
   l976 = 0;
   l978 = 0;
   l980 = 0;
   l982 = 0;
   l984 = 0;
   l986 = 0;
   l988 = 0;
   l990 = 0;
   l992 = 0;
   l994 = 0;
   l996 = 0;
   l998 = 0;
   l1000 = 0;
   l1002 = 0;
   l1004 = 0;
   l1006 = 0;
   l1008 = 0;
   l1010 = 0;
   l1012 = 0;
   l1014 = 0;
   l1016 = 0;
   l1018 = 0;
   l1020 = 0;
   l1022 = 0;
   l1024 = 0;
   l1026 = 0;
   l1028 = 0;
   l1030 = 0;
   l1032 = 0;
   l1034 = 0;
   l1036 = 0;
   l1038 = 0;
   l1040 = 0;
   l1042 = 0;
   l1044 = 0;
   l1046 = 0;
   l1048 = 0;
   l1050 = 0;
   l1052 = 0;
   l1054 = 0;
   l1056 = 0;
   l1058 = 0;
   l1060 = 0;
   l1062 = 0;
   l1064 = 0;
   l1066 = 0;
   l1068 = 0;
   l1070 = 0;
   l1072 = 0;
   l1074 = 0;
   l1076 = 0;
   l1078 = 0;
   l1080 = 0;
   l1082 = 0;
   l1084 = 0;
   l1086 = 0;
   l1088 = 0;
   l1090 = 0;
   l1092 = 0;
   l1094 = 0;
   l1096 = 0;
   l1098 = 0;
   l1100 = 0;
   l1102 = 0;
   l1104 = 0;
   l1106 = 0;
   l1108 = 0;
   l1110 = 0;
   l1112 = 0;
   l1114 = 0;
   l1116 = 0;
   l1118 = 0;
   l1120 = 0;
   l1122 = 0;
   l1124 = 0;
   l1126 = 0;
   l1128 = 0;
   l1130 = 0;
   l1132 = 0;
   l1134 = 0;
   l1136 = 0;
   l1138 = 0;
   l1140 = 0;
   l1142 = 0;
   l1144 = 0;
   l1146 = 0;
   l1148 = 0;
   l1150 = 0;
   l1152 = 0;
   l1154 = 0;
   l1156 = 0;
   l1158 = 0;
   l1160 = 0;
   l1162 = 0;
   l1164 = 0;
   l1166 = 0;
   l1168 = 0;
   l1170 = 0;
   l1172 = 0;
   l1174 = 0;
   l1176 = 0;
   l1178 = 0;
   l1180 = 0;
   l1182 = 0;
   l1184 = 0;
   l1186 = 0;
   l1188 = 0;
   l1190 = 0;
   l1192 = 0;
   l1194 = 0;
   l1196 = 0;
   l1198 = 0;
   l1200 = 0;
   l1202 = 0;
   l1204 = 0;
   l1206 = 0;
   l1208 = 0;
   l1210 = 0;
   l1212 = 0;
   l1214 = 0;
   l1216 = 0;
   l1218 = 0;
   l1220 = 0;
   l1222 = 0;
   l1224 = 0;
   l1226 = 0;
   l1228 = 0;
   l1230 = 0;
   l1232 = 0;
   l1234 = 0;
   l1236 = 0;
   l1238 = 0;
   l1240 = 0;
   l1242 = 0;
   l1244 = 0;
   l1246 = 0;
   l1248 = 0;
   l1250 = 0;
   l1252 = 0;
   l1254 = 0;
   l1256 = 0;
   l1258 = 0;
   l1260 = 0;
   l1262 = 0;
   l1264 = 0;
   l1266 = 0;
   l1268 = 0;
   l1270 = 0;
   l1272 = 0;
   l1274 = 0;
   l1276 = 0;
   l1278 = 0;
   l1280 = 0;
   l1282 = 0;
   l1284 = 0;
   l1286 = 0;
   l1288 = 0;
   l1290 = 0;
   l1292 = 0;
   l1294 = 0;
   l1296 = 0;
   l1298 = 0;
   l1300 = 0;
   l1302 = 0;
   l1304 = 0;
   l1306 = 0;
   l1308 = 0;
   l1310 = 0;
   l1312 = 0;
   l1314 = 0;
   l1316 = 0;
   l1318 = 0;
   l1320 = 0;
   l1322 = 0;
   l1324 = 0;
   l1326 = 0;
   l1328 = 0;
   l1330 = 0;
   l1332 = 0;
   l1334 = 0;
   l1336 = 0;
   l1338 = 0;
   l1340 = 0;
   l1342 = 0;
   l1344 = 0;
   l1346 = 0;
   l1348 = 0;
   l1350 = 0;
   l1352 = 0;
   l1354 = 0;
   l1356 = 0;
   l1358 = 0;
   l1360 = 0;
   l1362 = 0;
   l1364 = 0;
   l1366 = 0;
   l1368 = 0;
   l1370 = 0;
   l1372 = 0;
   l1374 = 0;
   l1376 = 0;
   l1378 = 0;
   l1380 = 0;
   l1382 = 0;
   l1384 = 0;
   l1386 = 0;
   l1388 = 0;
   l1390 = 0;
   l1392 = 0;
   l1394 = 0;
   l1396 = 0;
   l1398 = 0;
   l1400 = 0;
   l1402 = 0;
   l1404 = 0;
   l1406 = 0;
   l1408 = 0;
   l1410 = 0;
   l1412 = 0;
   l1414 = 0;
   l1416 = 0;
   l1418 = 0;
   l1420 = 0;
   l1422 = 0;
   l1424 = 0;
   l1426 = 0;
   l1428 = 0;
   l1430 = 0;
   l1432 = 0;
   l1434 = 0;
   l1436 = 0;
   l1438 = 0;
   l1440 = 0;
   l1442 = 0;
   l1444 = 0;
   l1446 = 0;
   l1448 = 0;
   l1450 = 0;
   l1452 = 0;
   l1454 = 0;
   l1456 = 0;
   l1458 = 0;
   l1460 = 0;
   l1462 = 0;
   l1464 = 0;
   l1466 = 0;
   l1468 = 0;
   l1470 = 0;
   l1472 = 0;
   l1474 = 0;
   l1476 = 0;
   l1478 = 0;
   l1480 = 0;
   l1482 = 0;
   l1484 = 0;
   l1486 = 0;
   l1488 = 0;
   l1490 = 0;
   l1492 = 0;
   l1494 = 0;
   l1496 = 0;
   l1498 = 0;
   l1500 = 0;
   l1502 = 0;
   l1504 = 0;
   l1506 = 0;
   l1508 = 0;
   l1510 = 0;
   l1512 = 0;
   l1514 = 0;
   l1516 = 0;
   l1518 = 0;
   l1520 = 0;
   l1522 = 0;
   l1524 = 0;
   l1526 = 0;
   l1528 = 0;
   l1530 = 0;
   l1532 = 0;
   l1534 = 0;
   l1536 = 0;
   l1538 = 0;
   l1540 = 0;
   l1542 = 0;
   l1544 = 0;
   l1546 = 0;
   l1548 = 0;
   l1550 = 0;
   l1552 = 0;
   l1554 = 0;
   l1556 = 0;
   l1558 = 0;
   l1560 = 0;
   l1562 = 0;
   l1564 = 0;
   l1566 = 0;
   l1568 = 0;
   l1570 = 0;
   l1572 = 0;
   l1574 = 0;
   l1576 = 0;
   l1578 = 0;
   l1580 = 0;
   l1582 = 0;
   l1584 = 0;
   l1586 = 0;
   l1588 = 0;
   l1590 = 0;
   l1592 = 0;
   l1594 = 0;
   l1596 = 0;
   l1598 = 0;
   l1600 = 0;
   l1602 = 0;
   l1604 = 0;
   l1606 = 0;
   l1608 = 0;
   l1610 = 0;
   l1612 = 0;
   l1614 = 0;
   l1616 = 0;
   l1618 = 0;
   l1620 = 0;
   l1622 = 0;
   l1624 = 0;
   l1626 = 0;
   l1628 = 0;
   l1630 = 0;
   l1632 = 0;
   l1634 = 0;
   l1636 = 0;
   l1638 = 0;
   l1640 = 0;
   l1642 = 0;
   l1644 = 0;
   l1646 = 0;
   l1648 = 0;
   l1650 = 0;
   l1652 = 0;
   l1654 = 0;
   l1656 = 0;
   l1658 = 0;
   l1660 = 0;
   l1662 = 0;
   l1664 = 0;
   l1666 = 0;
   l1668 = 0;
   l1670 = 0;
   l1672 = 0;
   l1674 = 0;
   l1676 = 0;
   l1678 = 0;
end

always @(posedge i2)
   l730 <= i2;

always @(posedge i4)
   l732 <= i4;

always @(posedge i6)
   l734 <= i6;

always @(posedge i8)
   l736 <= i8;

always @(posedge i10)
   l738 <= i10;

always @(posedge i12)
   l740 <= i12;

always @(posedge i14)
   l742 <= i14;

always @(posedge i16)
   l744 <= i16;

always @(posedge i18)
   l746 <= i18;

always @(posedge i20)
   l748 <= i20;

always @(posedge i22)
   l750 <= i22;

always @(posedge i24)
   l752 <= i24;

always @(posedge i26)
   l754 <= i26;

always @(posedge i28)
   l756 <= i28;

always @(posedge i30)
   l758 <= i30;

always @(posedge i32)
   l760 <= i32;

always @(posedge i34)
   l762 <= i34;

always @(posedge i36)
   l764 <= i36;

always @(posedge i38)
   l766 <= i38;

always @(posedge i40)
   l768 <= i40;

always @(posedge i42)
   l770 <= i42;

always @(posedge i44)
   l772 <= i44;

always @(posedge i46)
   l774 <= i46;

always @(posedge i48)
   l776 <= i48;

always @(posedge i50)
   l778 <= i50;

always @(posedge i52)
   l780 <= i52;

always @(posedge i54)
   l782 <= i54;

always @(posedge i56)
   l784 <= i56;

always @(posedge i58)
   l786 <= i58;

always @(posedge i60)
   l788 <= i60;

always @(posedge i62)
   l790 <= i62;

always @(posedge i64)
   l792 <= i64;

always @(posedge i66)
   l794 <= i66;

always @(posedge i68)
   l796 <= i68;

always @(posedge i70)
   l798 <= i70;

always @(posedge i72)
   l800 <= i72;

always @(posedge i74)
   l802 <= i74;

always @(posedge i76)
   l804 <= i76;

always @(posedge i78)
   l806 <= i78;

always @(posedge i80)
   l808 <= i80;

always @(posedge i82)
   l810 <= i82;

always @(posedge i84)
   l812 <= i84;

always @(posedge i86)
   l814 <= i86;

always @(posedge i88)
   l816 <= i88;

always @(posedge i90)
   l818 <= i90;

always @(posedge i92)
   l820 <= i92;

always @(posedge i94)
   l822 <= i94;

always @(posedge i96)
   l824 <= i96;

always @(posedge i98)
   l826 <= i98;

always @(posedge i100)
   l828 <= i100;

always @(posedge i102)
   l830 <= i102;

always @(posedge i104)
   l832 <= i104;

always @(posedge i106)
   l834 <= i106;

always @(posedge i108)
   l836 <= i108;

always @(posedge i110)
   l838 <= i110;

always @(posedge i112)
   l840 <= i112;

always @(posedge i114)
   l842 <= i114;

always @(posedge i116)
   l844 <= i116;

always @(posedge i118)
   l846 <= i118;

always @(posedge i120)
   l848 <= i120;

always @(posedge i122)
   l850 <= i122;

always @(posedge i124)
   l852 <= i124;

always @(posedge i126)
   l854 <= i126;

always @(posedge i128)
   l856 <= i128;

always @(posedge i130)
   l858 <= i130;

always @(posedge i132)
   l860 <= i132;

always @(posedge i134)
   l862 <= i134;

always @(posedge i136)
   l864 <= i136;

always @(posedge i138)
   l866 <= i138;

always @(posedge i140)
   l868 <= i140;

always @(posedge i142)
   l870 <= i142;

always @(posedge i144)
   l872 <= i144;

always @(posedge i146)
   l874 <= i146;

always @(posedge i148)
   l876 <= i148;

always @(posedge i150)
   l878 <= i150;

always @(posedge i152)
   l880 <= i152;

always @(posedge i154)
   l882 <= i154;

always @(posedge i156)
   l884 <= i156;

always @(posedge i158)
   l886 <= i158;

always @(posedge i160)
   l888 <= i160;

always @(posedge i162)
   l890 <= i162;

always @(posedge i164)
   l892 <= i164;

always @(posedge i166)
   l894 <= i166;

always @(posedge i168)
   l896 <= i168;

always @(posedge i170)
   l898 <= i170;

always @(posedge i172)
   l900 <= i172;

always @(posedge i174)
   l902 <= i174;

always @(posedge i176)
   l904 <= i176;

always @(posedge i178)
   l906 <= i178;

always @(posedge i180)
   l908 <= i180;

always @(posedge i182)
   l910 <= i182;

always @(posedge i184)
   l912 <= i184;

always @(posedge i186)
   l914 <= i186;

always @(posedge i188)
   l916 <= i188;

always @(posedge i190)
   l918 <= i190;

always @(posedge i192)
   l920 <= i192;

always @(posedge i194)
   l922 <= i194;

always @(posedge i196)
   l924 <= i196;

always @(posedge i198)
   l926 <= i198;

always @(posedge i200)
   l928 <= i200;

always @(posedge i202)
   l930 <= i202;

always @(posedge i204)
   l932 <= i204;

always @(posedge a1736)
   l934 <= a1736;

always @(posedge a1752)
   l936 <= a1752;

always @(posedge i206)
   l938 <= i206;

always @(posedge i208)
   l940 <= i208;

always @(posedge a1780)
   l942 <= a1780;

always @(posedge i210)
   l944 <= i210;

always @(posedge i212)
   l946 <= i212;

always @(posedge a1824)
   l948 <= a1824;

always @(posedge a1840)
   l950 <= a1840;

always @(posedge i214)
   l952 <= i214;

always @(posedge i216)
   l954 <= i216;

always @(posedge a1860)
   l956 <= a1860;

always @(posedge i218)
   l958 <= i218;

always @(posedge i220)
   l960 <= i220;

always @(posedge a1904)
   l962 <= a1904;

always @(posedge a1920)
   l964 <= a1920;

always @(posedge i222)
   l966 <= i222;

always @(posedge i224)
   l968 <= i224;

always @(posedge a1940)
   l970 <= a1940;

always @(posedge i226)
   l972 <= i226;

always @(posedge i228)
   l974 <= i228;

always @(posedge a1984)
   l976 <= a1984;

always @(posedge a2000)
   l978 <= a2000;

always @(posedge i230)
   l980 <= i230;

always @(posedge i232)
   l982 <= i232;

always @(posedge a2020)
   l984 <= a2020;

always @(posedge a2136)
   l986 <= a2136;

always @(posedge a2160)
   l988 <= a2160;

always @(posedge a2188)
   l990 <= a2188;

always @(posedge i234)
   l992 <= i234;

always @(posedge i236)
   l994 <= i236;

always @(posedge i238)
   l996 <= i238;

always @(posedge i240)
   l998 <= i240;

always @(posedge i242)
   l1000 <= i242;

always @(posedge a2200)
   l1002 <= a2200;

always @(posedge a2526)
   l1004 <= a2526;

always @(posedge a2536)
   l1006 <= a2536;

always @(posedge a2546)
   l1008 <= a2546;

always @(posedge a2556)
   l1010 <= a2556;

always @(posedge a2564)
   l1012 <= a2564;

always @(posedge i244)
   l1014 <= i244;

always @(posedge i246)
   l1016 <= i246;

always @(posedge a2622)
   l1018 <= a2622;

always @(posedge a2638)
   l1020 <= a2638;

always @(posedge i248)
   l1022 <= i248;

always @(posedge i250)
   l1024 <= i250;

always @(posedge a2666)
   l1026 <= a2666;

always @(posedge i252)
   l1028 <= i252;

always @(posedge i254)
   l1030 <= i254;

always @(posedge a2710)
   l1032 <= a2710;

always @(posedge a2726)
   l1034 <= a2726;

always @(posedge i256)
   l1036 <= i256;

always @(posedge i258)
   l1038 <= i258;

always @(posedge a2746)
   l1040 <= a2746;

always @(posedge i260)
   l1042 <= i260;

always @(posedge i262)
   l1044 <= i262;

always @(posedge a2790)
   l1046 <= a2790;

always @(posedge a2806)
   l1048 <= a2806;

always @(posedge i264)
   l1050 <= i264;

always @(posedge i266)
   l1052 <= i266;

always @(posedge a2826)
   l1054 <= a2826;

always @(posedge i268)
   l1056 <= i268;

always @(posedge i270)
   l1058 <= i270;

always @(posedge a2870)
   l1060 <= a2870;

always @(posedge a2886)
   l1062 <= a2886;

always @(posedge i272)
   l1064 <= i272;

always @(posedge i274)
   l1066 <= i274;

always @(posedge a2906)
   l1068 <= a2906;

always @(posedge a3022)
   l1070 <= a3022;

always @(posedge a3046)
   l1072 <= a3046;

always @(posedge a3074)
   l1074 <= a3074;

always @(posedge i276)
   l1076 <= i276;

always @(posedge i278)
   l1078 <= i278;

always @(posedge i280)
   l1080 <= i280;

always @(posedge i282)
   l1082 <= i282;

always @(posedge i284)
   l1084 <= i284;

always @(posedge a3086)
   l1086 <= a3086;

always @(posedge a3412)
   l1088 <= a3412;

always @(posedge a3422)
   l1090 <= a3422;

always @(posedge a3432)
   l1092 <= a3432;

always @(posedge a3442)
   l1094 <= a3442;

always @(posedge a3450)
   l1096 <= a3450;

always @(posedge i286)
   l1098 <= i286;

always @(posedge i288)
   l1100 <= i288;

always @(posedge a3508)
   l1102 <= a3508;

always @(posedge a3524)
   l1104 <= a3524;

always @(posedge i290)
   l1106 <= i290;

always @(posedge i292)
   l1108 <= i292;

always @(posedge a3552)
   l1110 <= a3552;

always @(posedge i294)
   l1112 <= i294;

always @(posedge i296)
   l1114 <= i296;

always @(posedge a3596)
   l1116 <= a3596;

always @(posedge a3612)
   l1118 <= a3612;

always @(posedge i298)
   l1120 <= i298;

always @(posedge i300)
   l1122 <= i300;

always @(posedge a3632)
   l1124 <= a3632;

always @(posedge i302)
   l1126 <= i302;

always @(posedge i304)
   l1128 <= i304;

always @(posedge a3676)
   l1130 <= a3676;

always @(posedge a3692)
   l1132 <= a3692;

always @(posedge i306)
   l1134 <= i306;

always @(posedge i308)
   l1136 <= i308;

always @(posedge a3712)
   l1138 <= a3712;

always @(posedge i310)
   l1140 <= i310;

always @(posedge i312)
   l1142 <= i312;

always @(posedge a3756)
   l1144 <= a3756;

always @(posedge a3772)
   l1146 <= a3772;

always @(posedge i314)
   l1148 <= i314;

always @(posedge i316)
   l1150 <= i316;

always @(posedge a3792)
   l1152 <= a3792;

always @(posedge a3908)
   l1154 <= a3908;

always @(posedge a3932)
   l1156 <= a3932;

always @(posedge a3960)
   l1158 <= a3960;

always @(posedge i318)
   l1160 <= i318;

always @(posedge i320)
   l1162 <= i320;

always @(posedge i322)
   l1164 <= i322;

always @(posedge i324)
   l1166 <= i324;

always @(posedge i326)
   l1168 <= i326;

always @(posedge a3972)
   l1170 <= a3972;

always @(posedge a4298)
   l1172 <= a4298;

always @(posedge a4308)
   l1174 <= a4308;

always @(posedge a4318)
   l1176 <= a4318;

always @(posedge a4328)
   l1178 <= a4328;

always @(posedge a4336)
   l1180 <= a4336;

always @(posedge i328)
   l1182 <= i328;

always @(posedge i330)
   l1184 <= i330;

always @(posedge a4394)
   l1186 <= a4394;

always @(posedge a4410)
   l1188 <= a4410;

always @(posedge i332)
   l1190 <= i332;

always @(posedge i334)
   l1192 <= i334;

always @(posedge a4438)
   l1194 <= a4438;

always @(posedge i336)
   l1196 <= i336;

always @(posedge i338)
   l1198 <= i338;

always @(posedge a4482)
   l1200 <= a4482;

always @(posedge a4498)
   l1202 <= a4498;

always @(posedge i340)
   l1204 <= i340;

always @(posedge i342)
   l1206 <= i342;

always @(posedge a4518)
   l1208 <= a4518;

always @(posedge i344)
   l1210 <= i344;

always @(posedge i346)
   l1212 <= i346;

always @(posedge a4562)
   l1214 <= a4562;

always @(posedge a4578)
   l1216 <= a4578;

always @(posedge i348)
   l1218 <= i348;

always @(posedge i350)
   l1220 <= i350;

always @(posedge a4598)
   l1222 <= a4598;

always @(posedge i352)
   l1224 <= i352;

always @(posedge i354)
   l1226 <= i354;

always @(posedge a4642)
   l1228 <= a4642;

always @(posedge a4658)
   l1230 <= a4658;

always @(posedge i356)
   l1232 <= i356;

always @(posedge i358)
   l1234 <= i358;

always @(posedge a4678)
   l1236 <= a4678;

always @(posedge a4794)
   l1238 <= a4794;

always @(posedge a4818)
   l1240 <= a4818;

always @(posedge a4846)
   l1242 <= a4846;

always @(posedge i360)
   l1244 <= i360;

always @(posedge i362)
   l1246 <= i362;

always @(posedge i364)
   l1248 <= i364;

always @(posedge i366)
   l1250 <= i366;

always @(posedge i368)
   l1252 <= i368;

always @(posedge a4858)
   l1254 <= a4858;

always @(posedge a5184)
   l1256 <= a5184;

always @(posedge a5194)
   l1258 <= a5194;

always @(posedge a5204)
   l1260 <= a5204;

always @(posedge a5214)
   l1262 <= a5214;

always @(posedge a5222)
   l1264 <= a5222;

always @(posedge i370)
   l1266 <= i370;

always @(posedge i372)
   l1268 <= i372;

always @(posedge a5280)
   l1270 <= a5280;

always @(posedge a5296)
   l1272 <= a5296;

always @(posedge i374)
   l1274 <= i374;

always @(posedge i376)
   l1276 <= i376;

always @(posedge a5324)
   l1278 <= a5324;

always @(posedge i378)
   l1280 <= i378;

always @(posedge i380)
   l1282 <= i380;

always @(posedge a5368)
   l1284 <= a5368;

always @(posedge a5384)
   l1286 <= a5384;

always @(posedge i382)
   l1288 <= i382;

always @(posedge i384)
   l1290 <= i384;

always @(posedge a5404)
   l1292 <= a5404;

always @(posedge i386)
   l1294 <= i386;

always @(posedge i388)
   l1296 <= i388;

always @(posedge a5448)
   l1298 <= a5448;

always @(posedge a5464)
   l1300 <= a5464;

always @(posedge i390)
   l1302 <= i390;

always @(posedge i392)
   l1304 <= i392;

always @(posedge a5484)
   l1306 <= a5484;

always @(posedge i394)
   l1308 <= i394;

always @(posedge i396)
   l1310 <= i396;

always @(posedge a5528)
   l1312 <= a5528;

always @(posedge a5544)
   l1314 <= a5544;

always @(posedge i398)
   l1316 <= i398;

always @(posedge i400)
   l1318 <= i400;

always @(posedge a5564)
   l1320 <= a5564;

always @(posedge a5680)
   l1322 <= a5680;

always @(posedge a5704)
   l1324 <= a5704;

always @(posedge a5732)
   l1326 <= a5732;

always @(posedge i402)
   l1328 <= i402;

always @(posedge i404)
   l1330 <= i404;

always @(posedge i406)
   l1332 <= i406;

always @(posedge i408)
   l1334 <= i408;

always @(posedge i410)
   l1336 <= i410;

always @(posedge a5744)
   l1338 <= a5744;

always @(posedge a6070)
   l1340 <= a6070;

always @(posedge a6080)
   l1342 <= a6080;

always @(posedge a6090)
   l1344 <= a6090;

always @(posedge a6100)
   l1346 <= a6100;

always @(posedge a6108)
   l1348 <= a6108;

always @(posedge i412)
   l1350 <= i412;

always @(posedge a6114)
   l1352 <= a6114;

always @(posedge i414)
   l1354 <= i414;

always @(posedge i416)
   l1356 <= i416;

always @(posedge i418)
   l1358 <= i418;

always @(posedge i420)
   l1360 <= i420;

always @(posedge i422)
   l1362 <= i422;

always @(posedge i424)
   l1364 <= i424;

always @(posedge i426)
   l1366 <= i426;

always @(posedge i428)
   l1368 <= i428;

always @(posedge i430)
   l1370 <= i430;

always @(posedge i432)
   l1372 <= i432;

always @(posedge i434)
   l1374 <= i434;

always @(posedge i436)
   l1376 <= i436;

always @(posedge i438)
   l1378 <= i438;

always @(posedge i440)
   l1380 <= i440;

always @(posedge i442)
   l1382 <= i442;

always @(posedge i444)
   l1384 <= i444;

always @(posedge i446)
   l1386 <= i446;

always @(posedge i448)
   l1388 <= i448;

always @(posedge i450)
   l1390 <= i450;

always @(posedge i452)
   l1392 <= i452;

always @(posedge i454)
   l1394 <= i454;

always @(posedge i456)
   l1396 <= i456;

always @(posedge i458)
   l1398 <= i458;

always @(posedge i460)
   l1400 <= i460;

always @(posedge i462)
   l1402 <= i462;

always @(posedge i464)
   l1404 <= i464;

always @(posedge i466)
   l1406 <= i466;

always @(posedge i468)
   l1408 <= i468;

always @(posedge i470)
   l1410 <= i470;

always @(posedge i472)
   l1412 <= i472;

always @(posedge i474)
   l1414 <= i474;

always @(posedge i476)
   l1416 <= i476;

always @(posedge i478)
   l1418 <= i478;

always @(posedge i480)
   l1420 <= i480;

always @(posedge i482)
   l1422 <= i482;

always @(posedge i484)
   l1424 <= i484;

always @(posedge i486)
   l1426 <= i486;

always @(posedge i488)
   l1428 <= i488;

always @(posedge i490)
   l1430 <= i490;

always @(posedge i492)
   l1432 <= i492;

always @(posedge i494)
   l1434 <= i494;

always @(posedge i496)
   l1436 <= i496;

always @(posedge i498)
   l1438 <= i498;

always @(posedge i500)
   l1440 <= i500;

always @(posedge i502)
   l1442 <= i502;

always @(posedge i504)
   l1444 <= i504;

always @(posedge i506)
   l1446 <= i506;

always @(posedge i508)
   l1448 <= i508;

always @(posedge i510)
   l1450 <= i510;

always @(posedge i512)
   l1452 <= i512;

always @(posedge i514)
   l1454 <= i514;

always @(posedge i516)
   l1456 <= i516;

always @(posedge i518)
   l1458 <= i518;

always @(posedge i520)
   l1460 <= i520;

always @(posedge i522)
   l1462 <= i522;

always @(posedge i524)
   l1464 <= i524;

always @(posedge i526)
   l1466 <= i526;

always @(posedge i528)
   l1468 <= i528;

always @(posedge i530)
   l1470 <= i530;

always @(posedge i532)
   l1472 <= i532;

always @(posedge i534)
   l1474 <= i534;

always @(posedge i536)
   l1476 <= i536;

always @(posedge i538)
   l1478 <= i538;

always @(posedge i540)
   l1480 <= i540;

always @(posedge i542)
   l1482 <= i542;

always @(posedge i544)
   l1484 <= i544;

always @(posedge i546)
   l1486 <= i546;

always @(posedge i548)
   l1488 <= i548;

always @(posedge i550)
   l1490 <= i550;

always @(posedge i552)
   l1492 <= i552;

always @(posedge i554)
   l1494 <= i554;

always @(posedge i556)
   l1496 <= i556;

always @(posedge i558)
   l1498 <= i558;

always @(posedge i560)
   l1500 <= i560;

always @(posedge i562)
   l1502 <= i562;

always @(posedge i564)
   l1504 <= i564;

always @(posedge i566)
   l1506 <= i566;

always @(posedge i568)
   l1508 <= i568;

always @(posedge i570)
   l1510 <= i570;

always @(posedge i572)
   l1512 <= i572;

always @(posedge i574)
   l1514 <= i574;

always @(posedge i576)
   l1516 <= i576;

always @(posedge i578)
   l1518 <= i578;

always @(posedge i580)
   l1520 <= i580;

always @(posedge i582)
   l1522 <= i582;

always @(posedge i584)
   l1524 <= i584;

always @(posedge i586)
   l1526 <= i586;

always @(posedge i588)
   l1528 <= i588;

always @(posedge i590)
   l1530 <= i590;

always @(posedge i592)
   l1532 <= i592;

always @(posedge i594)
   l1534 <= i594;

always @(posedge i596)
   l1536 <= i596;

always @(posedge i598)
   l1538 <= i598;

always @(posedge i600)
   l1540 <= i600;

always @(posedge i602)
   l1542 <= i602;

always @(posedge i604)
   l1544 <= i604;

always @(posedge i606)
   l1546 <= i606;

always @(posedge i608)
   l1548 <= i608;

always @(posedge i610)
   l1550 <= i610;

always @(posedge i612)
   l1552 <= i612;

always @(posedge i614)
   l1554 <= i614;

always @(posedge i616)
   l1556 <= i616;

always @(posedge i618)
   l1558 <= i618;

always @(posedge i620)
   l1560 <= i620;

always @(posedge i622)
   l1562 <= i622;

always @(posedge i624)
   l1564 <= i624;

always @(posedge i626)
   l1566 <= i626;

always @(posedge i628)
   l1568 <= i628;

always @(posedge i630)
   l1570 <= i630;

always @(posedge i632)
   l1572 <= i632;

always @(posedge i634)
   l1574 <= i634;

always @(posedge i636)
   l1576 <= i636;

always @(posedge i638)
   l1578 <= i638;

always @(posedge i640)
   l1580 <= i640;

always @(posedge i642)
   l1582 <= i642;

always @(posedge i644)
   l1584 <= i644;

always @(posedge i646)
   l1586 <= i646;

always @(posedge i648)
   l1588 <= i648;

always @(posedge i650)
   l1590 <= i650;

always @(posedge i652)
   l1592 <= i652;

always @(posedge i654)
   l1594 <= i654;

always @(posedge i656)
   l1596 <= i656;

always @(posedge i658)
   l1598 <= i658;

always @(posedge i660)
   l1600 <= i660;

always @(posedge i662)
   l1602 <= i662;

always @(posedge i664)
   l1604 <= i664;

always @(posedge i666)
   l1606 <= i666;

always @(posedge i668)
   l1608 <= i668;

always @(posedge i670)
   l1610 <= i670;

always @(posedge i672)
   l1612 <= i672;

always @(posedge i674)
   l1614 <= i674;

always @(posedge i676)
   l1616 <= i676;

always @(posedge i678)
   l1618 <= i678;

always @(posedge i680)
   l1620 <= i680;

always @(posedge i682)
   l1622 <= i682;

always @(posedge i684)
   l1624 <= i684;

always @(posedge i686)
   l1626 <= i686;

always @(posedge i688)
   l1628 <= i688;

always @(posedge i690)
   l1630 <= i690;

always @(posedge i692)
   l1632 <= i692;

always @(posedge i694)
   l1634 <= i694;

always @(posedge i696)
   l1636 <= i696;

always @(posedge i698)
   l1638 <= i698;

always @(posedge i700)
   l1640 <= i700;

always @(posedge i702)
   l1642 <= i702;

always @(posedge i704)
   l1644 <= i704;

always @(posedge i706)
   l1646 <= i706;

always @(posedge i708)
   l1648 <= i708;

always @(posedge i710)
   l1650 <= i710;

always @(posedge i712)
   l1652 <= i712;

always @(posedge i714)
   l1654 <= i714;

always @(posedge a6122)
   l1656 <= a6122;

always @(posedge a6132)
   l1658 <= a6132;

always @(posedge a6140)
   l1660 <= a6140;

always @(posedge i716)
   l1662 <= i716;

always @(posedge a6142)
   l1664 <= a6142;

always @(posedge i720)
   l1666 <= i720;

always @(posedge i722)
   l1668 <= i722;

always @(posedge i724)
   l1670 <= i724;

always @(posedge i726)
   l1672 <= i726;

always @(posedge i728)
   l1674 <= i728;

always @(posedge a26802)
   l1676 <= a26802;

always @(posedge c1)
   l1678 <= c1;


assign a1736 = a1734 & l1678;
assign a1752 = ~a1750 & l1678;
assign a1780 = ~a1778 & l1678;
assign a1824 = a1822 & l1678;
assign a1840 = ~a1838 & l1678;
assign a1860 = ~a1858 & l1678;
assign a1904 = a1902 & l1678;
assign a1920 = ~a1918 & l1678;
assign a1940 = ~a1938 & l1678;
assign a1984 = a1982 & l1678;
assign a2000 = ~a1998 & l1678;
assign a2020 = ~a2018 & l1678;
assign a2136 = a2134 & l1678;
assign a2160 = ~a2158 & l1678;
assign a2188 = ~a2186 & l1678;
assign a2200 = ~a2198 & l1678;
assign a2526 = a2524 & l1678;
assign a2536 = a2534 & l1678;
assign a2546 = a2544 & l1678;
assign a2556 = a2554 & l1678;
assign a2564 = a2562 & l1678;
assign a2622 = a2620 & l1678;
assign a2638 = ~a2636 & l1678;
assign a2666 = ~a2664 & l1678;
assign a2710 = a2708 & l1678;
assign a2726 = ~a2724 & l1678;
assign a2746 = ~a2744 & l1678;
assign a2790 = a2788 & l1678;
assign a2806 = ~a2804 & l1678;
assign a2826 = ~a2824 & l1678;
assign a2870 = a2868 & l1678;
assign a2886 = ~a2884 & l1678;
assign a2906 = ~a2904 & l1678;
assign a3022 = a3020 & l1678;
assign a3046 = ~a3044 & l1678;
assign a3074 = ~a3072 & l1678;
assign a3086 = ~a3084 & l1678;
assign a3412 = a3410 & l1678;
assign a3422 = a3420 & l1678;
assign a3432 = a3430 & l1678;
assign a3442 = a3440 & l1678;
assign a3450 = a3448 & l1678;
assign a3508 = a3506 & l1678;
assign a3524 = ~a3522 & l1678;
assign a3552 = ~a3550 & l1678;
assign a3596 = a3594 & l1678;
assign a3612 = ~a3610 & l1678;
assign a3632 = ~a3630 & l1678;
assign a3676 = a3674 & l1678;
assign a3692 = ~a3690 & l1678;
assign a3712 = ~a3710 & l1678;
assign a3756 = a3754 & l1678;
assign a3772 = ~a3770 & l1678;
assign a3792 = ~a3790 & l1678;
assign a3908 = a3906 & l1678;
assign a3932 = ~a3930 & l1678;
assign a3960 = ~a3958 & l1678;
assign a3972 = ~a3970 & l1678;
assign a4298 = a4296 & l1678;
assign a4308 = a4306 & l1678;
assign a4318 = a4316 & l1678;
assign a4328 = a4326 & l1678;
assign a4336 = a4334 & l1678;
assign a4394 = a4392 & l1678;
assign a4410 = ~a4408 & l1678;
assign a4438 = ~a4436 & l1678;
assign a4482 = a4480 & l1678;
assign a4498 = ~a4496 & l1678;
assign a4518 = ~a4516 & l1678;
assign a4562 = a4560 & l1678;
assign a4578 = ~a4576 & l1678;
assign a4598 = ~a4596 & l1678;
assign a4642 = a4640 & l1678;
assign a4658 = ~a4656 & l1678;
assign a4678 = ~a4676 & l1678;
assign a4794 = a4792 & l1678;
assign a4818 = ~a4816 & l1678;
assign a4846 = ~a4844 & l1678;
assign a4858 = ~a4856 & l1678;
assign a5184 = a5182 & l1678;
assign a5194 = a5192 & l1678;
assign a5204 = a5202 & l1678;
assign a5214 = a5212 & l1678;
assign a5222 = a5220 & l1678;
assign a5280 = a5278 & l1678;
assign a5296 = ~a5294 & l1678;
assign a5324 = ~a5322 & l1678;
assign a5368 = a5366 & l1678;
assign a5384 = ~a5382 & l1678;
assign a5404 = ~a5402 & l1678;
assign a5448 = a5446 & l1678;
assign a5464 = ~a5462 & l1678;
assign a5484 = ~a5482 & l1678;
assign a5528 = a5526 & l1678;
assign a5544 = ~a5542 & l1678;
assign a5564 = ~a5562 & l1678;
assign a5680 = a5678 & l1678;
assign a5704 = ~a5702 & l1678;
assign a5732 = ~a5730 & l1678;
assign a5744 = ~a5742 & l1678;
assign a6070 = a6068 & l1678;
assign a6080 = a6078 & l1678;
assign a6090 = a6088 & l1678;
assign a6100 = a6098 & l1678;
assign a6108 = a6106 & l1678;
assign a6114 = ~a6112 & l1678;
assign a6122 = ~a6120 & l1678;
assign a6132 = ~a6130 & l1678;
assign a6140 = ~a6138 & l1678;
assign a6142 = ~a6116 & l1678;
assign a26802 = a26800 & l1678;
assign c1 = 1;
assign a1680 = l942 & ~l940;
assign a1682 = l990 & l988;
assign a1684 = a1682 & ~l986;
assign a1686 = a1684 & a1680;
assign a1688 = ~l942 & l940;
assign a1690 = a1688 & a1684;
assign a1692 = l990 & ~l988;
assign a1694 = a1692 & l986;
assign a1696 = a1694 & a1688;
assign a1698 = l932 & ~l930;
assign a1700 = a1682 & l986;
assign a1702 = a1700 & a1688;
assign a1704 = a1702 & a1698;
assign a1706 = ~l932 & ~l930;
assign a1708 = l942 & l940;
assign a1710 = a1692 & ~l986;
assign a1712 = a1710 & a1708;
assign a1714 = a1712 & a1706;
assign a1716 = a1710 & a1680;
assign a1718 = a1716 & a1698;
assign a1720 = a1710 & l992;
assign a1722 = ~a1720 & l934;
assign a1724 = a1722 & ~a1718;
assign a1726 = a1724 & ~a1714;
assign a1728 = ~a1726 & ~a1704;
assign a1730 = ~a1728 & ~a1696;
assign a1732 = ~a1730 & ~a1690;
assign a1734 = ~a1732 & ~a1686;
assign a1738 = ~a1720 & l936;
assign a1740 = a1738 & ~a1718;
assign a1742 = a1740 & ~a1714;
assign a1744 = ~a1742 & ~a1704;
assign a1746 = ~a1744 & ~a1696;
assign a1748 = ~a1746 & ~a1690;
assign a1750 = a1748 & ~a1686;
assign a1754 = ~l932 & l930;
assign a1756 = ~l990 & ~l988;
assign a1758 = a1756 & ~l986;
assign a1760 = a1758 & a1688;
assign a1762 = a1760 & a1754;
assign a1764 = ~l990 & l988;
assign a1766 = a1764 & ~l986;
assign a1768 = a1766 & a1688;
assign a1770 = a1768 & a1706;
assign a1772 = a1754 & a1702;
assign a1774 = ~a1772 & ~l942;
assign a1776 = a1774 & ~a1770;
assign a1778 = a1776 & ~a1762;
assign a1782 = l956 & ~l954;
assign a1784 = a1782 & a1684;
assign a1786 = ~l956 & l954;
assign a1788 = a1786 & a1684;
assign a1790 = a1786 & a1694;
assign a1792 = l946 & ~l944;
assign a1794 = a1786 & a1700;
assign a1796 = a1794 & a1792;
assign a1798 = ~l946 & ~l944;
assign a1800 = l956 & l954;
assign a1802 = a1800 & a1710;
assign a1804 = a1802 & a1798;
assign a1806 = a1782 & a1710;
assign a1808 = a1806 & a1792;
assign a1810 = ~a1720 & l948;
assign a1812 = a1810 & ~a1808;
assign a1814 = a1812 & ~a1804;
assign a1816 = ~a1814 & ~a1796;
assign a1818 = ~a1816 & ~a1790;
assign a1820 = ~a1818 & ~a1788;
assign a1822 = ~a1820 & ~a1784;
assign a1826 = ~a1720 & l950;
assign a1828 = a1826 & ~a1808;
assign a1830 = a1828 & ~a1804;
assign a1832 = ~a1830 & ~a1796;
assign a1834 = ~a1832 & ~a1790;
assign a1836 = ~a1834 & ~a1788;
assign a1838 = a1836 & ~a1784;
assign a1842 = ~l946 & l944;
assign a1844 = a1786 & a1758;
assign a1846 = a1844 & a1842;
assign a1848 = a1786 & a1766;
assign a1850 = a1848 & a1798;
assign a1852 = a1842 & a1794;
assign a1854 = ~a1852 & ~l956;
assign a1856 = a1854 & ~a1850;
assign a1858 = a1856 & ~a1846;
assign a1862 = l970 & ~l968;
assign a1864 = a1862 & a1684;
assign a1866 = ~l970 & l968;
assign a1868 = a1866 & a1684;
assign a1870 = a1866 & a1694;
assign a1872 = l960 & ~l958;
assign a1874 = a1866 & a1700;
assign a1876 = a1874 & a1872;
assign a1878 = ~l960 & ~l958;
assign a1880 = l970 & l968;
assign a1882 = a1880 & a1710;
assign a1884 = a1882 & a1878;
assign a1886 = a1862 & a1710;
assign a1888 = a1886 & a1872;
assign a1890 = ~a1720 & l962;
assign a1892 = a1890 & ~a1888;
assign a1894 = a1892 & ~a1884;
assign a1896 = ~a1894 & ~a1876;
assign a1898 = ~a1896 & ~a1870;
assign a1900 = ~a1898 & ~a1868;
assign a1902 = ~a1900 & ~a1864;
assign a1906 = ~a1720 & l964;
assign a1908 = a1906 & ~a1888;
assign a1910 = a1908 & ~a1884;
assign a1912 = ~a1910 & ~a1876;
assign a1914 = ~a1912 & ~a1870;
assign a1916 = ~a1914 & ~a1868;
assign a1918 = a1916 & ~a1864;
assign a1922 = ~l960 & l958;
assign a1924 = a1866 & a1758;
assign a1926 = a1924 & a1922;
assign a1928 = a1866 & a1766;
assign a1930 = a1928 & a1878;
assign a1932 = a1922 & a1874;
assign a1934 = ~a1932 & ~l970;
assign a1936 = a1934 & ~a1930;
assign a1938 = a1936 & ~a1926;
assign a1942 = l984 & ~l982;
assign a1944 = a1942 & a1684;
assign a1946 = ~l984 & l982;
assign a1948 = a1946 & a1684;
assign a1950 = a1946 & a1694;
assign a1952 = l974 & ~l972;
assign a1954 = a1946 & a1700;
assign a1956 = a1954 & a1952;
assign a1958 = ~l974 & ~l972;
assign a1960 = l984 & l982;
assign a1962 = a1960 & a1710;
assign a1964 = a1962 & a1958;
assign a1966 = a1942 & a1710;
assign a1968 = a1966 & a1952;
assign a1970 = ~a1720 & l976;
assign a1972 = a1970 & ~a1968;
assign a1974 = a1972 & ~a1964;
assign a1976 = ~a1974 & ~a1956;
assign a1978 = ~a1976 & ~a1950;
assign a1980 = ~a1978 & ~a1948;
assign a1982 = ~a1980 & ~a1944;
assign a1986 = ~a1720 & l978;
assign a1988 = a1986 & ~a1968;
assign a1990 = a1988 & ~a1964;
assign a1992 = ~a1990 & ~a1956;
assign a1994 = ~a1992 & ~a1950;
assign a1996 = ~a1994 & ~a1948;
assign a1998 = a1996 & ~a1944;
assign a2002 = ~l974 & l972;
assign a2004 = a1946 & a1758;
assign a2006 = a2004 & a2002;
assign a2008 = a1946 & a1766;
assign a2010 = a2008 & a1958;
assign a2012 = a2002 & a1954;
assign a2014 = ~a2012 & ~l984;
assign a2016 = a2014 & ~a2010;
assign a2018 = a2016 & ~a2006;
assign a2022 = l1012 & l1010;
assign a2024 = ~a2022 & ~l1008;
assign a2026 = ~a2024 & l1006;
assign a2028 = ~a2026 & ~l1004;
assign a2030 = a2028 & l998;
assign a2032 = ~a1786 & ~a1688;
assign a2034 = a2032 & ~a1866;
assign a2036 = a1786 & a1688;
assign a2038 = ~a2036 & ~a1866;
assign a2040 = ~a2038 & ~a2032;
assign a2042 = ~a2040 & ~a1946;
assign a2044 = ~a2042 & ~a2034;
assign a2046 = ~a2044 & a1758;
assign a2048 = a2046 & ~a2030;
assign a2050 = ~a1698 & a1680;
assign a2052 = ~a2050 & a1684;
assign a2054 = ~a1792 & a1782;
assign a2056 = ~a2054 & a2052;
assign a2058 = ~a1872 & a1862;
assign a2060 = ~a2058 & a2056;
assign a2062 = ~a1952 & a1942;
assign a2064 = ~a2062 & a2060;
assign a2066 = ~a1706 & a1688;
assign a2068 = ~a2066 & a1766;
assign a2070 = ~a1798 & a1786;
assign a2072 = ~a2070 & a2068;
assign a2074 = ~a1878 & a1866;
assign a2076 = ~a2074 & a2072;
assign a2078 = ~a1958 & a1946;
assign a2080 = ~a2078 & a2076;
assign a2082 = ~a2002 & a1946;
assign a2084 = ~a1922 & a1866;
assign a2086 = ~a1842 & a1786;
assign a2088 = ~a1754 & a1688;
assign a2090 = ~a2088 & a1766;
assign a2092 = a2090 & ~a2086;
assign a2094 = a2092 & ~a2084;
assign a2096 = a2094 & ~a2082;
assign a2098 = ~a1952 & a1946;
assign a2100 = ~a1872 & a1866;
assign a2102 = ~a1698 & a1688;
assign a2104 = ~a1792 & a1786;
assign a2106 = ~a2104 & ~a2102;
assign a2108 = a2106 & ~a2100;
assign a2110 = a2108 & ~a2098;
assign a2112 = ~a2088 & ~a2086;
assign a2114 = a2112 & ~a2084;
assign a2116 = a2114 & ~a2082;
assign a2118 = ~a2116 & ~a2110;
assign a2120 = ~a2118 & ~a1692;
assign a2122 = a2120 & a1700;
assign a2124 = a2122 & ~a1756;
assign a2126 = ~a2124 & l986;
assign a2128 = ~a2126 & ~a2096;
assign a2130 = ~a2128 & ~a2080;
assign a2132 = a2130 & ~a2064;
assign a2134 = a2132 & ~a2048;
assign a2138 = a1694 & ~l1000;
assign a2140 = a1756 & l986;
assign a2142 = l990 & l986;
assign a2144 = a2142 & l1000;
assign a2146 = ~a2144 & a2140;
assign a2148 = ~a2146 & ~l988;
assign a2150 = a2148 & ~a2138;
assign a2152 = ~a2150 & ~a2096;
assign a2154 = a2152 & ~a2080;
assign a2156 = ~a2154 & ~a2064;
assign a2158 = a2156 & ~a2048;
assign a2162 = a1694 & l1000;
assign a2164 = ~a2100 & ~a2098;
assign a2166 = a2164 & ~a2104;
assign a2168 = a2166 & ~a2102;
assign a2170 = a2168 & a1700;
assign a2172 = ~a2170 & l990;
assign a2174 = ~a2172 & ~a2140;
assign a2176 = ~a2174 & ~a2162;
assign a2178 = ~a2176 & ~a2138;
assign a2180 = a2178 & ~a2096;
assign a2182 = a2180 & ~a2080;
assign a2184 = ~a2182 & ~a2064;
assign a2186 = ~a2184 & ~a2048;
assign a2190 = ~l1010 & ~l1008;
assign a2192 = a2190 & ~l1006;
assign a2194 = ~a2192 & l1004;
assign a2196 = a2194 & a1758;
assign a2198 = ~a2196 & ~l1002;
assign a2202 = ~l1012 & ~l1010;
assign a2204 = a2202 & ~l1008;
assign a2206 = a2204 & ~l1006;
assign a2208 = a2206 & ~l1004;
assign a2210 = l1012 & ~l1010;
assign a2212 = a2210 & ~l1008;
assign a2214 = a2212 & ~l1006;
assign a2216 = a2214 & ~l1004;
assign a2218 = ~l1012 & l1010;
assign a2220 = a2218 & ~l1008;
assign a2222 = a2220 & ~l1006;
assign a2224 = a2222 & ~l1004;
assign a2226 = a2022 & ~l1008;
assign a2228 = a2226 & ~l1006;
assign a2230 = a2228 & ~l1004;
assign a2232 = a2202 & l1008;
assign a2234 = a2232 & ~l1006;
assign a2236 = a2234 & ~l1004;
assign a2238 = a2210 & l1008;
assign a2240 = a2238 & ~l1006;
assign a2242 = a2240 & ~l1004;
assign a2244 = a2218 & l1008;
assign a2246 = a2244 & ~l1006;
assign a2248 = a2246 & ~l1004;
assign a2250 = a2022 & l1008;
assign a2252 = a2250 & ~l1006;
assign a2254 = a2252 & ~l1004;
assign a2256 = l1006 & ~l1004;
assign a2258 = ~a2218 & a2024;
assign a2260 = a2258 & ~a2212;
assign a2262 = a2260 & ~a2204;
assign a2264 = ~a2262 & a2256;
assign a2266 = a2264 & ~a2254;
assign a2268 = a2266 & ~a2248;
assign a2270 = a2268 & ~a2242;
assign a2272 = a2270 & ~a2236;
assign a2274 = a2272 & ~a2230;
assign a2276 = a2274 & ~a2224;
assign a2278 = a2276 & ~a2216;
assign a2280 = a2278 & ~a2208;
assign a2282 = l1008 & ~l1004;
assign a2284 = a2022 & ~l1006;
assign a2286 = a2204 & l1006;
assign a2288 = a2286 & ~l1004;
assign a2290 = a2212 & l1006;
assign a2292 = a2290 & ~l1004;
assign a2294 = a2220 & l1006;
assign a2296 = a2294 & ~l1004;
assign a2298 = a2226 & l1006;
assign a2300 = a2298 & ~l1004;
assign a2302 = ~a2300 & l1006;
assign a2304 = a2302 & ~a2296;
assign a2306 = a2304 & ~a2292;
assign a2308 = a2306 & ~a2288;
assign a2310 = ~a2308 & ~a2284;
assign a2312 = a2218 & ~l1006;
assign a2314 = ~a2312 & a2310;
assign a2316 = a2210 & ~l1006;
assign a2318 = ~a2316 & a2314;
assign a2320 = a2202 & ~l1006;
assign a2322 = ~a2320 & a2318;
assign a2324 = ~a2322 & a2282;
assign a2326 = a2324 & ~a2230;
assign a2328 = a2326 & ~a2224;
assign a2330 = a2328 & ~a2216;
assign a2332 = a2330 & ~a2208;
assign a2334 = a2192 & ~l1004;
assign a2336 = l1010 & ~l1008;
assign a2338 = a2336 & ~l1006;
assign a2340 = a2338 & ~l1004;
assign a2342 = ~l1010 & l1008;
assign a2344 = a2342 & ~l1006;
assign a2346 = a2344 & ~l1004;
assign a2348 = l1010 & l1008;
assign a2350 = a2348 & ~l1006;
assign a2352 = a2350 & ~l1004;
assign a2354 = a2190 & l1006;
assign a2356 = a2354 & ~l1004;
assign a2358 = a2336 & l1006;
assign a2360 = a2358 & ~l1004;
assign a2362 = a2232 & l1006;
assign a2364 = a2362 & ~l1004;
assign a2366 = a2342 & l1006;
assign a2368 = a2366 & ~l1004;
assign a2370 = a2244 & l1006;
assign a2372 = a2370 & ~l1004;
assign a2374 = a2348 & l1006;
assign a2376 = a2374 & ~l1004;
assign a2378 = a2192 & l1004;
assign a2380 = a2378 & ~a2206;
assign a2382 = ~a2380 & ~a2376;
assign a2384 = ~a2382 & ~a2372;
assign a2386 = ~a2384 & ~a2368;
assign a2388 = ~a2386 & ~a2364;
assign a2390 = ~a2388 & ~a2360;
assign a2392 = ~a2390 & ~a2296;
assign a2394 = ~a2392 & ~a2356;
assign a2396 = ~a2394 & ~a2288;
assign a2398 = ~a2396 & ~a2352;
assign a2400 = ~a2398 & ~a2248;
assign a2402 = ~a2400 & ~a2346;
assign a2404 = ~a2402 & ~a2236;
assign a2406 = ~a2404 & ~a2340;
assign a2408 = ~a2406 & ~a2224;
assign a2410 = ~a2408 & ~a2334;
assign a2412 = ~a2410 & l1012;
assign a2414 = a2412 & ~a2208;
assign a2416 = l1012 & ~l1008;
assign a2418 = a2416 & ~l1006;
assign a2420 = a2418 & ~l1004;
assign a2422 = l1012 & l1008;
assign a2424 = a2422 & ~l1006;
assign a2426 = a2424 & ~l1004;
assign a2428 = a2416 & l1006;
assign a2430 = a2428 & ~l1004;
assign a2432 = a2422 & l1006;
assign a2434 = a2432 & ~l1004;
assign a2436 = ~l1008 & ~l1006;
assign a2438 = a2436 & l1004;
assign a2440 = ~a2438 & ~a2434;
assign a2442 = ~l1012 & l1008;
assign a2444 = a2442 & l1006;
assign a2446 = a2444 & ~l1004;
assign a2448 = ~a2446 & a2440;
assign a2450 = ~a2448 & ~a2300;
assign a2452 = a2450 & ~a2296;
assign a2454 = ~a2452 & ~a2430;
assign a2456 = ~l1012 & ~l1008;
assign a2458 = a2456 & l1006;
assign a2460 = a2458 & ~l1004;
assign a2462 = ~a2460 & a2454;
assign a2464 = ~a2462 & ~a2254;
assign a2466 = a2464 & ~a2248;
assign a2468 = ~a2466 & ~a2426;
assign a2470 = a2442 & ~l1006;
assign a2472 = a2470 & ~l1004;
assign a2474 = ~a2472 & a2468;
assign a2476 = ~a2474 & ~a2230;
assign a2478 = a2476 & ~a2224;
assign a2480 = ~a2478 & ~a2420;
assign a2482 = a2456 & ~l1006;
assign a2484 = a2482 & ~l1004;
assign a2486 = ~a2484 & a2480;
assign a2488 = ~a2486 & ~l1010;
assign a2490 = ~a2488 & a2414;
assign a2492 = a2490 & ~a2332;
assign a2494 = a2492 & ~a2280;
assign a2496 = ~a2262 & l1006;
assign a2498 = ~a2496 & ~a2252;
assign a2500 = a2498 & ~a2246;
assign a2502 = a2500 & ~a2240;
assign a2504 = a2502 & ~a2234;
assign a2506 = a2504 & ~a2228;
assign a2508 = a2506 & ~a2222;
assign a2510 = a2508 & ~a2214;
assign a2512 = a2510 & ~a2206;
assign a2514 = ~a2512 & ~l1004;
assign a2516 = ~a2514 & a2494;
assign a2518 = ~a2516 & l1004;
assign a2520 = ~a2518 & a1758;
assign a2522 = ~a1758 & ~l1004;
assign a2524 = ~a2522 & ~a2520;
assign a2528 = ~a2516 & l1006;
assign a2530 = ~a2528 & a1758;
assign a2532 = ~a1758 & ~l1006;
assign a2534 = ~a2532 & ~a2530;
assign a2538 = ~a2516 & l1008;
assign a2540 = ~a2538 & a1758;
assign a2542 = ~a1758 & ~l1008;
assign a2544 = ~a2542 & ~a2540;
assign a2548 = ~a2516 & l1010;
assign a2550 = ~a2548 & a1758;
assign a2552 = ~a1758 & ~l1010;
assign a2554 = ~a2552 & ~a2550;
assign a2558 = a1758 & l1012;
assign a2560 = ~a1758 & ~l1012;
assign a2562 = ~a2560 & ~a2558;
assign a2566 = l1026 & ~l1024;
assign a2568 = l1074 & l1072;
assign a2570 = a2568 & ~l1070;
assign a2572 = a2570 & a2566;
assign a2574 = ~l1026 & l1024;
assign a2576 = a2574 & a2570;
assign a2578 = l1074 & ~l1072;
assign a2580 = a2578 & l1070;
assign a2582 = a2580 & a2574;
assign a2584 = l1016 & ~l1014;
assign a2586 = a2568 & l1070;
assign a2588 = a2586 & a2574;
assign a2590 = a2588 & a2584;
assign a2592 = ~l1016 & ~l1014;
assign a2594 = l1026 & l1024;
assign a2596 = a2578 & ~l1070;
assign a2598 = a2596 & a2594;
assign a2600 = a2598 & a2592;
assign a2602 = a2596 & a2566;
assign a2604 = a2602 & a2584;
assign a2606 = a2596 & l1076;
assign a2608 = ~a2606 & l1018;
assign a2610 = a2608 & ~a2604;
assign a2612 = a2610 & ~a2600;
assign a2614 = ~a2612 & ~a2590;
assign a2616 = ~a2614 & ~a2582;
assign a2618 = ~a2616 & ~a2576;
assign a2620 = ~a2618 & ~a2572;
assign a2624 = ~a2606 & l1020;
assign a2626 = a2624 & ~a2604;
assign a2628 = a2626 & ~a2600;
assign a2630 = ~a2628 & ~a2590;
assign a2632 = ~a2630 & ~a2582;
assign a2634 = ~a2632 & ~a2576;
assign a2636 = a2634 & ~a2572;
assign a2640 = ~l1016 & l1014;
assign a2642 = ~l1074 & ~l1072;
assign a2644 = a2642 & ~l1070;
assign a2646 = a2644 & a2574;
assign a2648 = a2646 & a2640;
assign a2650 = ~l1074 & l1072;
assign a2652 = a2650 & ~l1070;
assign a2654 = a2652 & a2574;
assign a2656 = a2654 & a2592;
assign a2658 = a2640 & a2588;
assign a2660 = ~a2658 & ~l1026;
assign a2662 = a2660 & ~a2656;
assign a2664 = a2662 & ~a2648;
assign a2668 = l1040 & ~l1038;
assign a2670 = a2668 & a2570;
assign a2672 = ~l1040 & l1038;
assign a2674 = a2672 & a2570;
assign a2676 = a2672 & a2580;
assign a2678 = l1030 & ~l1028;
assign a2680 = a2672 & a2586;
assign a2682 = a2680 & a2678;
assign a2684 = ~l1030 & ~l1028;
assign a2686 = l1040 & l1038;
assign a2688 = a2686 & a2596;
assign a2690 = a2688 & a2684;
assign a2692 = a2668 & a2596;
assign a2694 = a2692 & a2678;
assign a2696 = ~a2606 & l1032;
assign a2698 = a2696 & ~a2694;
assign a2700 = a2698 & ~a2690;
assign a2702 = ~a2700 & ~a2682;
assign a2704 = ~a2702 & ~a2676;
assign a2706 = ~a2704 & ~a2674;
assign a2708 = ~a2706 & ~a2670;
assign a2712 = ~a2606 & l1034;
assign a2714 = a2712 & ~a2694;
assign a2716 = a2714 & ~a2690;
assign a2718 = ~a2716 & ~a2682;
assign a2720 = ~a2718 & ~a2676;
assign a2722 = ~a2720 & ~a2674;
assign a2724 = a2722 & ~a2670;
assign a2728 = ~l1030 & l1028;
assign a2730 = a2672 & a2644;
assign a2732 = a2730 & a2728;
assign a2734 = a2672 & a2652;
assign a2736 = a2734 & a2684;
assign a2738 = a2728 & a2680;
assign a2740 = ~a2738 & ~l1040;
assign a2742 = a2740 & ~a2736;
assign a2744 = a2742 & ~a2732;
assign a2748 = l1054 & ~l1052;
assign a2750 = a2748 & a2570;
assign a2752 = ~l1054 & l1052;
assign a2754 = a2752 & a2570;
assign a2756 = a2752 & a2580;
assign a2758 = l1044 & ~l1042;
assign a2760 = a2752 & a2586;
assign a2762 = a2760 & a2758;
assign a2764 = ~l1044 & ~l1042;
assign a2766 = l1054 & l1052;
assign a2768 = a2766 & a2596;
assign a2770 = a2768 & a2764;
assign a2772 = a2748 & a2596;
assign a2774 = a2772 & a2758;
assign a2776 = ~a2606 & l1046;
assign a2778 = a2776 & ~a2774;
assign a2780 = a2778 & ~a2770;
assign a2782 = ~a2780 & ~a2762;
assign a2784 = ~a2782 & ~a2756;
assign a2786 = ~a2784 & ~a2754;
assign a2788 = ~a2786 & ~a2750;
assign a2792 = ~a2606 & l1048;
assign a2794 = a2792 & ~a2774;
assign a2796 = a2794 & ~a2770;
assign a2798 = ~a2796 & ~a2762;
assign a2800 = ~a2798 & ~a2756;
assign a2802 = ~a2800 & ~a2754;
assign a2804 = a2802 & ~a2750;
assign a2808 = ~l1044 & l1042;
assign a2810 = a2752 & a2644;
assign a2812 = a2810 & a2808;
assign a2814 = a2752 & a2652;
assign a2816 = a2814 & a2764;
assign a2818 = a2808 & a2760;
assign a2820 = ~a2818 & ~l1054;
assign a2822 = a2820 & ~a2816;
assign a2824 = a2822 & ~a2812;
assign a2828 = l1068 & ~l1066;
assign a2830 = a2828 & a2570;
assign a2832 = ~l1068 & l1066;
assign a2834 = a2832 & a2570;
assign a2836 = a2832 & a2580;
assign a2838 = l1058 & ~l1056;
assign a2840 = a2832 & a2586;
assign a2842 = a2840 & a2838;
assign a2844 = ~l1058 & ~l1056;
assign a2846 = l1068 & l1066;
assign a2848 = a2846 & a2596;
assign a2850 = a2848 & a2844;
assign a2852 = a2828 & a2596;
assign a2854 = a2852 & a2838;
assign a2856 = ~a2606 & l1060;
assign a2858 = a2856 & ~a2854;
assign a2860 = a2858 & ~a2850;
assign a2862 = ~a2860 & ~a2842;
assign a2864 = ~a2862 & ~a2836;
assign a2866 = ~a2864 & ~a2834;
assign a2868 = ~a2866 & ~a2830;
assign a2872 = ~a2606 & l1062;
assign a2874 = a2872 & ~a2854;
assign a2876 = a2874 & ~a2850;
assign a2878 = ~a2876 & ~a2842;
assign a2880 = ~a2878 & ~a2836;
assign a2882 = ~a2880 & ~a2834;
assign a2884 = a2882 & ~a2830;
assign a2888 = ~l1058 & l1056;
assign a2890 = a2832 & a2644;
assign a2892 = a2890 & a2888;
assign a2894 = a2832 & a2652;
assign a2896 = a2894 & a2844;
assign a2898 = a2888 & a2840;
assign a2900 = ~a2898 & ~l1068;
assign a2902 = a2900 & ~a2896;
assign a2904 = a2902 & ~a2892;
assign a2908 = l1096 & l1094;
assign a2910 = ~a2908 & ~l1092;
assign a2912 = ~a2910 & l1090;
assign a2914 = ~a2912 & ~l1088;
assign a2916 = a2914 & l1082;
assign a2918 = ~a2672 & ~a2574;
assign a2920 = a2918 & ~a2752;
assign a2922 = a2672 & a2574;
assign a2924 = ~a2922 & ~a2752;
assign a2926 = ~a2924 & ~a2918;
assign a2928 = ~a2926 & ~a2832;
assign a2930 = ~a2928 & ~a2920;
assign a2932 = ~a2930 & a2644;
assign a2934 = a2932 & ~a2916;
assign a2936 = ~a2584 & a2566;
assign a2938 = ~a2936 & a2570;
assign a2940 = ~a2678 & a2668;
assign a2942 = ~a2940 & a2938;
assign a2944 = ~a2758 & a2748;
assign a2946 = ~a2944 & a2942;
assign a2948 = ~a2838 & a2828;
assign a2950 = ~a2948 & a2946;
assign a2952 = ~a2592 & a2574;
assign a2954 = ~a2952 & a2652;
assign a2956 = ~a2684 & a2672;
assign a2958 = ~a2956 & a2954;
assign a2960 = ~a2764 & a2752;
assign a2962 = ~a2960 & a2958;
assign a2964 = ~a2844 & a2832;
assign a2966 = ~a2964 & a2962;
assign a2968 = ~a2888 & a2832;
assign a2970 = ~a2808 & a2752;
assign a2972 = ~a2728 & a2672;
assign a2974 = ~a2640 & a2574;
assign a2976 = ~a2974 & a2652;
assign a2978 = a2976 & ~a2972;
assign a2980 = a2978 & ~a2970;
assign a2982 = a2980 & ~a2968;
assign a2984 = ~a2838 & a2832;
assign a2986 = ~a2758 & a2752;
assign a2988 = ~a2584 & a2574;
assign a2990 = ~a2678 & a2672;
assign a2992 = ~a2990 & ~a2988;
assign a2994 = a2992 & ~a2986;
assign a2996 = a2994 & ~a2984;
assign a2998 = ~a2974 & ~a2972;
assign a3000 = a2998 & ~a2970;
assign a3002 = a3000 & ~a2968;
assign a3004 = ~a3002 & ~a2996;
assign a3006 = ~a3004 & ~a2578;
assign a3008 = a3006 & a2586;
assign a3010 = a3008 & ~a2642;
assign a3012 = ~a3010 & l1070;
assign a3014 = ~a3012 & ~a2982;
assign a3016 = ~a3014 & ~a2966;
assign a3018 = a3016 & ~a2950;
assign a3020 = a3018 & ~a2934;
assign a3024 = a2580 & ~l1084;
assign a3026 = a2642 & l1070;
assign a3028 = l1074 & l1070;
assign a3030 = a3028 & l1084;
assign a3032 = ~a3030 & a3026;
assign a3034 = ~a3032 & ~l1072;
assign a3036 = a3034 & ~a3024;
assign a3038 = ~a3036 & ~a2982;
assign a3040 = a3038 & ~a2966;
assign a3042 = ~a3040 & ~a2950;
assign a3044 = a3042 & ~a2934;
assign a3048 = a2580 & l1084;
assign a3050 = ~a2986 & ~a2984;
assign a3052 = a3050 & ~a2990;
assign a3054 = a3052 & ~a2988;
assign a3056 = a3054 & a2586;
assign a3058 = ~a3056 & l1074;
assign a3060 = ~a3058 & ~a3026;
assign a3062 = ~a3060 & ~a3048;
assign a3064 = ~a3062 & ~a3024;
assign a3066 = a3064 & ~a2982;
assign a3068 = a3066 & ~a2966;
assign a3070 = ~a3068 & ~a2950;
assign a3072 = ~a3070 & ~a2934;
assign a3076 = ~l1094 & ~l1092;
assign a3078 = a3076 & ~l1090;
assign a3080 = ~a3078 & l1088;
assign a3082 = a3080 & a2644;
assign a3084 = ~a3082 & ~l1086;
assign a3088 = ~l1096 & ~l1094;
assign a3090 = a3088 & ~l1092;
assign a3092 = a3090 & ~l1090;
assign a3094 = a3092 & ~l1088;
assign a3096 = l1096 & ~l1094;
assign a3098 = a3096 & ~l1092;
assign a3100 = a3098 & ~l1090;
assign a3102 = a3100 & ~l1088;
assign a3104 = ~l1096 & l1094;
assign a3106 = a3104 & ~l1092;
assign a3108 = a3106 & ~l1090;
assign a3110 = a3108 & ~l1088;
assign a3112 = a2908 & ~l1092;
assign a3114 = a3112 & ~l1090;
assign a3116 = a3114 & ~l1088;
assign a3118 = a3088 & l1092;
assign a3120 = a3118 & ~l1090;
assign a3122 = a3120 & ~l1088;
assign a3124 = a3096 & l1092;
assign a3126 = a3124 & ~l1090;
assign a3128 = a3126 & ~l1088;
assign a3130 = a3104 & l1092;
assign a3132 = a3130 & ~l1090;
assign a3134 = a3132 & ~l1088;
assign a3136 = a2908 & l1092;
assign a3138 = a3136 & ~l1090;
assign a3140 = a3138 & ~l1088;
assign a3142 = l1090 & ~l1088;
assign a3144 = ~a3104 & a2910;
assign a3146 = a3144 & ~a3098;
assign a3148 = a3146 & ~a3090;
assign a3150 = ~a3148 & a3142;
assign a3152 = a3150 & ~a3140;
assign a3154 = a3152 & ~a3134;
assign a3156 = a3154 & ~a3128;
assign a3158 = a3156 & ~a3122;
assign a3160 = a3158 & ~a3116;
assign a3162 = a3160 & ~a3110;
assign a3164 = a3162 & ~a3102;
assign a3166 = a3164 & ~a3094;
assign a3168 = l1092 & ~l1088;
assign a3170 = a2908 & ~l1090;
assign a3172 = a3090 & l1090;
assign a3174 = a3172 & ~l1088;
assign a3176 = a3098 & l1090;
assign a3178 = a3176 & ~l1088;
assign a3180 = a3106 & l1090;
assign a3182 = a3180 & ~l1088;
assign a3184 = a3112 & l1090;
assign a3186 = a3184 & ~l1088;
assign a3188 = ~a3186 & l1090;
assign a3190 = a3188 & ~a3182;
assign a3192 = a3190 & ~a3178;
assign a3194 = a3192 & ~a3174;
assign a3196 = ~a3194 & ~a3170;
assign a3198 = a3104 & ~l1090;
assign a3200 = ~a3198 & a3196;
assign a3202 = a3096 & ~l1090;
assign a3204 = ~a3202 & a3200;
assign a3206 = a3088 & ~l1090;
assign a3208 = ~a3206 & a3204;
assign a3210 = ~a3208 & a3168;
assign a3212 = a3210 & ~a3116;
assign a3214 = a3212 & ~a3110;
assign a3216 = a3214 & ~a3102;
assign a3218 = a3216 & ~a3094;
assign a3220 = a3078 & ~l1088;
assign a3222 = l1094 & ~l1092;
assign a3224 = a3222 & ~l1090;
assign a3226 = a3224 & ~l1088;
assign a3228 = ~l1094 & l1092;
assign a3230 = a3228 & ~l1090;
assign a3232 = a3230 & ~l1088;
assign a3234 = l1094 & l1092;
assign a3236 = a3234 & ~l1090;
assign a3238 = a3236 & ~l1088;
assign a3240 = a3076 & l1090;
assign a3242 = a3240 & ~l1088;
assign a3244 = a3222 & l1090;
assign a3246 = a3244 & ~l1088;
assign a3248 = a3118 & l1090;
assign a3250 = a3248 & ~l1088;
assign a3252 = a3228 & l1090;
assign a3254 = a3252 & ~l1088;
assign a3256 = a3130 & l1090;
assign a3258 = a3256 & ~l1088;
assign a3260 = a3234 & l1090;
assign a3262 = a3260 & ~l1088;
assign a3264 = a3078 & l1088;
assign a3266 = a3264 & ~a3092;
assign a3268 = ~a3266 & ~a3262;
assign a3270 = ~a3268 & ~a3258;
assign a3272 = ~a3270 & ~a3254;
assign a3274 = ~a3272 & ~a3250;
assign a3276 = ~a3274 & ~a3246;
assign a3278 = ~a3276 & ~a3182;
assign a3280 = ~a3278 & ~a3242;
assign a3282 = ~a3280 & ~a3174;
assign a3284 = ~a3282 & ~a3238;
assign a3286 = ~a3284 & ~a3134;
assign a3288 = ~a3286 & ~a3232;
assign a3290 = ~a3288 & ~a3122;
assign a3292 = ~a3290 & ~a3226;
assign a3294 = ~a3292 & ~a3110;
assign a3296 = ~a3294 & ~a3220;
assign a3298 = ~a3296 & l1096;
assign a3300 = a3298 & ~a3094;
assign a3302 = l1096 & ~l1092;
assign a3304 = a3302 & ~l1090;
assign a3306 = a3304 & ~l1088;
assign a3308 = l1096 & l1092;
assign a3310 = a3308 & ~l1090;
assign a3312 = a3310 & ~l1088;
assign a3314 = a3302 & l1090;
assign a3316 = a3314 & ~l1088;
assign a3318 = a3308 & l1090;
assign a3320 = a3318 & ~l1088;
assign a3322 = ~l1092 & ~l1090;
assign a3324 = a3322 & l1088;
assign a3326 = ~a3324 & ~a3320;
assign a3328 = ~l1096 & l1092;
assign a3330 = a3328 & l1090;
assign a3332 = a3330 & ~l1088;
assign a3334 = ~a3332 & a3326;
assign a3336 = ~a3334 & ~a3186;
assign a3338 = a3336 & ~a3182;
assign a3340 = ~a3338 & ~a3316;
assign a3342 = ~l1096 & ~l1092;
assign a3344 = a3342 & l1090;
assign a3346 = a3344 & ~l1088;
assign a3348 = ~a3346 & a3340;
assign a3350 = ~a3348 & ~a3140;
assign a3352 = a3350 & ~a3134;
assign a3354 = ~a3352 & ~a3312;
assign a3356 = a3328 & ~l1090;
assign a3358 = a3356 & ~l1088;
assign a3360 = ~a3358 & a3354;
assign a3362 = ~a3360 & ~a3116;
assign a3364 = a3362 & ~a3110;
assign a3366 = ~a3364 & ~a3306;
assign a3368 = a3342 & ~l1090;
assign a3370 = a3368 & ~l1088;
assign a3372 = ~a3370 & a3366;
assign a3374 = ~a3372 & ~l1094;
assign a3376 = ~a3374 & a3300;
assign a3378 = a3376 & ~a3218;
assign a3380 = a3378 & ~a3166;
assign a3382 = ~a3148 & l1090;
assign a3384 = ~a3382 & ~a3138;
assign a3386 = a3384 & ~a3132;
assign a3388 = a3386 & ~a3126;
assign a3390 = a3388 & ~a3120;
assign a3392 = a3390 & ~a3114;
assign a3394 = a3392 & ~a3108;
assign a3396 = a3394 & ~a3100;
assign a3398 = a3396 & ~a3092;
assign a3400 = ~a3398 & ~l1088;
assign a3402 = ~a3400 & a3380;
assign a3404 = ~a3402 & l1088;
assign a3406 = ~a3404 & a2644;
assign a3408 = ~a2644 & ~l1088;
assign a3410 = ~a3408 & ~a3406;
assign a3414 = ~a3402 & l1090;
assign a3416 = ~a3414 & a2644;
assign a3418 = ~a2644 & ~l1090;
assign a3420 = ~a3418 & ~a3416;
assign a3424 = ~a3402 & l1092;
assign a3426 = ~a3424 & a2644;
assign a3428 = ~a2644 & ~l1092;
assign a3430 = ~a3428 & ~a3426;
assign a3434 = ~a3402 & l1094;
assign a3436 = ~a3434 & a2644;
assign a3438 = ~a2644 & ~l1094;
assign a3440 = ~a3438 & ~a3436;
assign a3444 = a2644 & l1096;
assign a3446 = ~a2644 & ~l1096;
assign a3448 = ~a3446 & ~a3444;
assign a3452 = l1110 & ~l1108;
assign a3454 = l1158 & l1156;
assign a3456 = a3454 & ~l1154;
assign a3458 = a3456 & a3452;
assign a3460 = ~l1110 & l1108;
assign a3462 = a3460 & a3456;
assign a3464 = l1158 & ~l1156;
assign a3466 = a3464 & l1154;
assign a3468 = a3466 & a3460;
assign a3470 = l1100 & ~l1098;
assign a3472 = a3454 & l1154;
assign a3474 = a3472 & a3460;
assign a3476 = a3474 & a3470;
assign a3478 = ~l1100 & ~l1098;
assign a3480 = l1110 & l1108;
assign a3482 = a3464 & ~l1154;
assign a3484 = a3482 & a3480;
assign a3486 = a3484 & a3478;
assign a3488 = a3482 & a3452;
assign a3490 = a3488 & a3470;
assign a3492 = a3482 & l1160;
assign a3494 = ~a3492 & l1102;
assign a3496 = a3494 & ~a3490;
assign a3498 = a3496 & ~a3486;
assign a3500 = ~a3498 & ~a3476;
assign a3502 = ~a3500 & ~a3468;
assign a3504 = ~a3502 & ~a3462;
assign a3506 = ~a3504 & ~a3458;
assign a3510 = ~a3492 & l1104;
assign a3512 = a3510 & ~a3490;
assign a3514 = a3512 & ~a3486;
assign a3516 = ~a3514 & ~a3476;
assign a3518 = ~a3516 & ~a3468;
assign a3520 = ~a3518 & ~a3462;
assign a3522 = a3520 & ~a3458;
assign a3526 = ~l1100 & l1098;
assign a3528 = ~l1158 & ~l1156;
assign a3530 = a3528 & ~l1154;
assign a3532 = a3530 & a3460;
assign a3534 = a3532 & a3526;
assign a3536 = ~l1158 & l1156;
assign a3538 = a3536 & ~l1154;
assign a3540 = a3538 & a3460;
assign a3542 = a3540 & a3478;
assign a3544 = a3526 & a3474;
assign a3546 = ~a3544 & ~l1110;
assign a3548 = a3546 & ~a3542;
assign a3550 = a3548 & ~a3534;
assign a3554 = l1124 & ~l1122;
assign a3556 = a3554 & a3456;
assign a3558 = ~l1124 & l1122;
assign a3560 = a3558 & a3456;
assign a3562 = a3558 & a3466;
assign a3564 = l1114 & ~l1112;
assign a3566 = a3558 & a3472;
assign a3568 = a3566 & a3564;
assign a3570 = ~l1114 & ~l1112;
assign a3572 = l1124 & l1122;
assign a3574 = a3572 & a3482;
assign a3576 = a3574 & a3570;
assign a3578 = a3554 & a3482;
assign a3580 = a3578 & a3564;
assign a3582 = ~a3492 & l1116;
assign a3584 = a3582 & ~a3580;
assign a3586 = a3584 & ~a3576;
assign a3588 = ~a3586 & ~a3568;
assign a3590 = ~a3588 & ~a3562;
assign a3592 = ~a3590 & ~a3560;
assign a3594 = ~a3592 & ~a3556;
assign a3598 = ~a3492 & l1118;
assign a3600 = a3598 & ~a3580;
assign a3602 = a3600 & ~a3576;
assign a3604 = ~a3602 & ~a3568;
assign a3606 = ~a3604 & ~a3562;
assign a3608 = ~a3606 & ~a3560;
assign a3610 = a3608 & ~a3556;
assign a3614 = ~l1114 & l1112;
assign a3616 = a3558 & a3530;
assign a3618 = a3616 & a3614;
assign a3620 = a3558 & a3538;
assign a3622 = a3620 & a3570;
assign a3624 = a3614 & a3566;
assign a3626 = ~a3624 & ~l1124;
assign a3628 = a3626 & ~a3622;
assign a3630 = a3628 & ~a3618;
assign a3634 = l1138 & ~l1136;
assign a3636 = a3634 & a3456;
assign a3638 = ~l1138 & l1136;
assign a3640 = a3638 & a3456;
assign a3642 = a3638 & a3466;
assign a3644 = l1128 & ~l1126;
assign a3646 = a3638 & a3472;
assign a3648 = a3646 & a3644;
assign a3650 = ~l1128 & ~l1126;
assign a3652 = l1138 & l1136;
assign a3654 = a3652 & a3482;
assign a3656 = a3654 & a3650;
assign a3658 = a3634 & a3482;
assign a3660 = a3658 & a3644;
assign a3662 = ~a3492 & l1130;
assign a3664 = a3662 & ~a3660;
assign a3666 = a3664 & ~a3656;
assign a3668 = ~a3666 & ~a3648;
assign a3670 = ~a3668 & ~a3642;
assign a3672 = ~a3670 & ~a3640;
assign a3674 = ~a3672 & ~a3636;
assign a3678 = ~a3492 & l1132;
assign a3680 = a3678 & ~a3660;
assign a3682 = a3680 & ~a3656;
assign a3684 = ~a3682 & ~a3648;
assign a3686 = ~a3684 & ~a3642;
assign a3688 = ~a3686 & ~a3640;
assign a3690 = a3688 & ~a3636;
assign a3694 = ~l1128 & l1126;
assign a3696 = a3638 & a3530;
assign a3698 = a3696 & a3694;
assign a3700 = a3638 & a3538;
assign a3702 = a3700 & a3650;
assign a3704 = a3694 & a3646;
assign a3706 = ~a3704 & ~l1138;
assign a3708 = a3706 & ~a3702;
assign a3710 = a3708 & ~a3698;
assign a3714 = l1152 & ~l1150;
assign a3716 = a3714 & a3456;
assign a3718 = ~l1152 & l1150;
assign a3720 = a3718 & a3456;
assign a3722 = a3718 & a3466;
assign a3724 = l1142 & ~l1140;
assign a3726 = a3718 & a3472;
assign a3728 = a3726 & a3724;
assign a3730 = ~l1142 & ~l1140;
assign a3732 = l1152 & l1150;
assign a3734 = a3732 & a3482;
assign a3736 = a3734 & a3730;
assign a3738 = a3714 & a3482;
assign a3740 = a3738 & a3724;
assign a3742 = ~a3492 & l1144;
assign a3744 = a3742 & ~a3740;
assign a3746 = a3744 & ~a3736;
assign a3748 = ~a3746 & ~a3728;
assign a3750 = ~a3748 & ~a3722;
assign a3752 = ~a3750 & ~a3720;
assign a3754 = ~a3752 & ~a3716;
assign a3758 = ~a3492 & l1146;
assign a3760 = a3758 & ~a3740;
assign a3762 = a3760 & ~a3736;
assign a3764 = ~a3762 & ~a3728;
assign a3766 = ~a3764 & ~a3722;
assign a3768 = ~a3766 & ~a3720;
assign a3770 = a3768 & ~a3716;
assign a3774 = ~l1142 & l1140;
assign a3776 = a3718 & a3530;
assign a3778 = a3776 & a3774;
assign a3780 = a3718 & a3538;
assign a3782 = a3780 & a3730;
assign a3784 = a3774 & a3726;
assign a3786 = ~a3784 & ~l1152;
assign a3788 = a3786 & ~a3782;
assign a3790 = a3788 & ~a3778;
assign a3794 = l1180 & l1178;
assign a3796 = ~a3794 & ~l1176;
assign a3798 = ~a3796 & l1174;
assign a3800 = ~a3798 & ~l1172;
assign a3802 = a3800 & l1166;
assign a3804 = ~a3558 & ~a3460;
assign a3806 = a3804 & ~a3638;
assign a3808 = a3558 & a3460;
assign a3810 = ~a3808 & ~a3638;
assign a3812 = ~a3810 & ~a3804;
assign a3814 = ~a3812 & ~a3718;
assign a3816 = ~a3814 & ~a3806;
assign a3818 = ~a3816 & a3530;
assign a3820 = a3818 & ~a3802;
assign a3822 = ~a3470 & a3452;
assign a3824 = ~a3822 & a3456;
assign a3826 = ~a3564 & a3554;
assign a3828 = ~a3826 & a3824;
assign a3830 = ~a3644 & a3634;
assign a3832 = ~a3830 & a3828;
assign a3834 = ~a3724 & a3714;
assign a3836 = ~a3834 & a3832;
assign a3838 = ~a3478 & a3460;
assign a3840 = ~a3838 & a3538;
assign a3842 = ~a3570 & a3558;
assign a3844 = ~a3842 & a3840;
assign a3846 = ~a3650 & a3638;
assign a3848 = ~a3846 & a3844;
assign a3850 = ~a3730 & a3718;
assign a3852 = ~a3850 & a3848;
assign a3854 = ~a3774 & a3718;
assign a3856 = ~a3694 & a3638;
assign a3858 = ~a3614 & a3558;
assign a3860 = ~a3526 & a3460;
assign a3862 = ~a3860 & a3538;
assign a3864 = a3862 & ~a3858;
assign a3866 = a3864 & ~a3856;
assign a3868 = a3866 & ~a3854;
assign a3870 = ~a3724 & a3718;
assign a3872 = ~a3644 & a3638;
assign a3874 = ~a3470 & a3460;
assign a3876 = ~a3564 & a3558;
assign a3878 = ~a3876 & ~a3874;
assign a3880 = a3878 & ~a3872;
assign a3882 = a3880 & ~a3870;
assign a3884 = ~a3860 & ~a3858;
assign a3886 = a3884 & ~a3856;
assign a3888 = a3886 & ~a3854;
assign a3890 = ~a3888 & ~a3882;
assign a3892 = ~a3890 & ~a3464;
assign a3894 = a3892 & a3472;
assign a3896 = a3894 & ~a3528;
assign a3898 = ~a3896 & l1154;
assign a3900 = ~a3898 & ~a3868;
assign a3902 = ~a3900 & ~a3852;
assign a3904 = a3902 & ~a3836;
assign a3906 = a3904 & ~a3820;
assign a3910 = a3466 & ~l1168;
assign a3912 = a3528 & l1154;
assign a3914 = l1158 & l1154;
assign a3916 = a3914 & l1168;
assign a3918 = ~a3916 & a3912;
assign a3920 = ~a3918 & ~l1156;
assign a3922 = a3920 & ~a3910;
assign a3924 = ~a3922 & ~a3868;
assign a3926 = a3924 & ~a3852;
assign a3928 = ~a3926 & ~a3836;
assign a3930 = a3928 & ~a3820;
assign a3934 = a3466 & l1168;
assign a3936 = ~a3872 & ~a3870;
assign a3938 = a3936 & ~a3876;
assign a3940 = a3938 & ~a3874;
assign a3942 = a3940 & a3472;
assign a3944 = ~a3942 & l1158;
assign a3946 = ~a3944 & ~a3912;
assign a3948 = ~a3946 & ~a3934;
assign a3950 = ~a3948 & ~a3910;
assign a3952 = a3950 & ~a3868;
assign a3954 = a3952 & ~a3852;
assign a3956 = ~a3954 & ~a3836;
assign a3958 = ~a3956 & ~a3820;
assign a3962 = ~l1178 & ~l1176;
assign a3964 = a3962 & ~l1174;
assign a3966 = ~a3964 & l1172;
assign a3968 = a3966 & a3530;
assign a3970 = ~a3968 & ~l1170;
assign a3974 = ~l1180 & ~l1178;
assign a3976 = a3974 & ~l1176;
assign a3978 = a3976 & ~l1174;
assign a3980 = a3978 & ~l1172;
assign a3982 = l1180 & ~l1178;
assign a3984 = a3982 & ~l1176;
assign a3986 = a3984 & ~l1174;
assign a3988 = a3986 & ~l1172;
assign a3990 = ~l1180 & l1178;
assign a3992 = a3990 & ~l1176;
assign a3994 = a3992 & ~l1174;
assign a3996 = a3994 & ~l1172;
assign a3998 = a3794 & ~l1176;
assign a4000 = a3998 & ~l1174;
assign a4002 = a4000 & ~l1172;
assign a4004 = a3974 & l1176;
assign a4006 = a4004 & ~l1174;
assign a4008 = a4006 & ~l1172;
assign a4010 = a3982 & l1176;
assign a4012 = a4010 & ~l1174;
assign a4014 = a4012 & ~l1172;
assign a4016 = a3990 & l1176;
assign a4018 = a4016 & ~l1174;
assign a4020 = a4018 & ~l1172;
assign a4022 = a3794 & l1176;
assign a4024 = a4022 & ~l1174;
assign a4026 = a4024 & ~l1172;
assign a4028 = l1174 & ~l1172;
assign a4030 = ~a3990 & a3796;
assign a4032 = a4030 & ~a3984;
assign a4034 = a4032 & ~a3976;
assign a4036 = ~a4034 & a4028;
assign a4038 = a4036 & ~a4026;
assign a4040 = a4038 & ~a4020;
assign a4042 = a4040 & ~a4014;
assign a4044 = a4042 & ~a4008;
assign a4046 = a4044 & ~a4002;
assign a4048 = a4046 & ~a3996;
assign a4050 = a4048 & ~a3988;
assign a4052 = a4050 & ~a3980;
assign a4054 = l1176 & ~l1172;
assign a4056 = a3794 & ~l1174;
assign a4058 = a3976 & l1174;
assign a4060 = a4058 & ~l1172;
assign a4062 = a3984 & l1174;
assign a4064 = a4062 & ~l1172;
assign a4066 = a3992 & l1174;
assign a4068 = a4066 & ~l1172;
assign a4070 = a3998 & l1174;
assign a4072 = a4070 & ~l1172;
assign a4074 = ~a4072 & l1174;
assign a4076 = a4074 & ~a4068;
assign a4078 = a4076 & ~a4064;
assign a4080 = a4078 & ~a4060;
assign a4082 = ~a4080 & ~a4056;
assign a4084 = a3990 & ~l1174;
assign a4086 = ~a4084 & a4082;
assign a4088 = a3982 & ~l1174;
assign a4090 = ~a4088 & a4086;
assign a4092 = a3974 & ~l1174;
assign a4094 = ~a4092 & a4090;
assign a4096 = ~a4094 & a4054;
assign a4098 = a4096 & ~a4002;
assign a4100 = a4098 & ~a3996;
assign a4102 = a4100 & ~a3988;
assign a4104 = a4102 & ~a3980;
assign a4106 = a3964 & ~l1172;
assign a4108 = l1178 & ~l1176;
assign a4110 = a4108 & ~l1174;
assign a4112 = a4110 & ~l1172;
assign a4114 = ~l1178 & l1176;
assign a4116 = a4114 & ~l1174;
assign a4118 = a4116 & ~l1172;
assign a4120 = l1178 & l1176;
assign a4122 = a4120 & ~l1174;
assign a4124 = a4122 & ~l1172;
assign a4126 = a3962 & l1174;
assign a4128 = a4126 & ~l1172;
assign a4130 = a4108 & l1174;
assign a4132 = a4130 & ~l1172;
assign a4134 = a4004 & l1174;
assign a4136 = a4134 & ~l1172;
assign a4138 = a4114 & l1174;
assign a4140 = a4138 & ~l1172;
assign a4142 = a4016 & l1174;
assign a4144 = a4142 & ~l1172;
assign a4146 = a4120 & l1174;
assign a4148 = a4146 & ~l1172;
assign a4150 = a3964 & l1172;
assign a4152 = a4150 & ~a3978;
assign a4154 = ~a4152 & ~a4148;
assign a4156 = ~a4154 & ~a4144;
assign a4158 = ~a4156 & ~a4140;
assign a4160 = ~a4158 & ~a4136;
assign a4162 = ~a4160 & ~a4132;
assign a4164 = ~a4162 & ~a4068;
assign a4166 = ~a4164 & ~a4128;
assign a4168 = ~a4166 & ~a4060;
assign a4170 = ~a4168 & ~a4124;
assign a4172 = ~a4170 & ~a4020;
assign a4174 = ~a4172 & ~a4118;
assign a4176 = ~a4174 & ~a4008;
assign a4178 = ~a4176 & ~a4112;
assign a4180 = ~a4178 & ~a3996;
assign a4182 = ~a4180 & ~a4106;
assign a4184 = ~a4182 & l1180;
assign a4186 = a4184 & ~a3980;
assign a4188 = l1180 & ~l1176;
assign a4190 = a4188 & ~l1174;
assign a4192 = a4190 & ~l1172;
assign a4194 = l1180 & l1176;
assign a4196 = a4194 & ~l1174;
assign a4198 = a4196 & ~l1172;
assign a4200 = a4188 & l1174;
assign a4202 = a4200 & ~l1172;
assign a4204 = a4194 & l1174;
assign a4206 = a4204 & ~l1172;
assign a4208 = ~l1176 & ~l1174;
assign a4210 = a4208 & l1172;
assign a4212 = ~a4210 & ~a4206;
assign a4214 = ~l1180 & l1176;
assign a4216 = a4214 & l1174;
assign a4218 = a4216 & ~l1172;
assign a4220 = ~a4218 & a4212;
assign a4222 = ~a4220 & ~a4072;
assign a4224 = a4222 & ~a4068;
assign a4226 = ~a4224 & ~a4202;
assign a4228 = ~l1180 & ~l1176;
assign a4230 = a4228 & l1174;
assign a4232 = a4230 & ~l1172;
assign a4234 = ~a4232 & a4226;
assign a4236 = ~a4234 & ~a4026;
assign a4238 = a4236 & ~a4020;
assign a4240 = ~a4238 & ~a4198;
assign a4242 = a4214 & ~l1174;
assign a4244 = a4242 & ~l1172;
assign a4246 = ~a4244 & a4240;
assign a4248 = ~a4246 & ~a4002;
assign a4250 = a4248 & ~a3996;
assign a4252 = ~a4250 & ~a4192;
assign a4254 = a4228 & ~l1174;
assign a4256 = a4254 & ~l1172;
assign a4258 = ~a4256 & a4252;
assign a4260 = ~a4258 & ~l1178;
assign a4262 = ~a4260 & a4186;
assign a4264 = a4262 & ~a4104;
assign a4266 = a4264 & ~a4052;
assign a4268 = ~a4034 & l1174;
assign a4270 = ~a4268 & ~a4024;
assign a4272 = a4270 & ~a4018;
assign a4274 = a4272 & ~a4012;
assign a4276 = a4274 & ~a4006;
assign a4278 = a4276 & ~a4000;
assign a4280 = a4278 & ~a3994;
assign a4282 = a4280 & ~a3986;
assign a4284 = a4282 & ~a3978;
assign a4286 = ~a4284 & ~l1172;
assign a4288 = ~a4286 & a4266;
assign a4290 = ~a4288 & l1172;
assign a4292 = ~a4290 & a3530;
assign a4294 = ~a3530 & ~l1172;
assign a4296 = ~a4294 & ~a4292;
assign a4300 = ~a4288 & l1174;
assign a4302 = ~a4300 & a3530;
assign a4304 = ~a3530 & ~l1174;
assign a4306 = ~a4304 & ~a4302;
assign a4310 = ~a4288 & l1176;
assign a4312 = ~a4310 & a3530;
assign a4314 = ~a3530 & ~l1176;
assign a4316 = ~a4314 & ~a4312;
assign a4320 = ~a4288 & l1178;
assign a4322 = ~a4320 & a3530;
assign a4324 = ~a3530 & ~l1178;
assign a4326 = ~a4324 & ~a4322;
assign a4330 = a3530 & l1180;
assign a4332 = ~a3530 & ~l1180;
assign a4334 = ~a4332 & ~a4330;
assign a4338 = l1194 & ~l1192;
assign a4340 = l1242 & l1240;
assign a4342 = a4340 & ~l1238;
assign a4344 = a4342 & a4338;
assign a4346 = ~l1194 & l1192;
assign a4348 = a4346 & a4342;
assign a4350 = l1242 & ~l1240;
assign a4352 = a4350 & l1238;
assign a4354 = a4352 & a4346;
assign a4356 = l1184 & ~l1182;
assign a4358 = a4340 & l1238;
assign a4360 = a4358 & a4346;
assign a4362 = a4360 & a4356;
assign a4364 = ~l1184 & ~l1182;
assign a4366 = l1194 & l1192;
assign a4368 = a4350 & ~l1238;
assign a4370 = a4368 & a4366;
assign a4372 = a4370 & a4364;
assign a4374 = a4368 & a4338;
assign a4376 = a4374 & a4356;
assign a4378 = a4368 & l1244;
assign a4380 = ~a4378 & l1186;
assign a4382 = a4380 & ~a4376;
assign a4384 = a4382 & ~a4372;
assign a4386 = ~a4384 & ~a4362;
assign a4388 = ~a4386 & ~a4354;
assign a4390 = ~a4388 & ~a4348;
assign a4392 = ~a4390 & ~a4344;
assign a4396 = ~a4378 & l1188;
assign a4398 = a4396 & ~a4376;
assign a4400 = a4398 & ~a4372;
assign a4402 = ~a4400 & ~a4362;
assign a4404 = ~a4402 & ~a4354;
assign a4406 = ~a4404 & ~a4348;
assign a4408 = a4406 & ~a4344;
assign a4412 = ~l1184 & l1182;
assign a4414 = ~l1242 & ~l1240;
assign a4416 = a4414 & ~l1238;
assign a4418 = a4416 & a4346;
assign a4420 = a4418 & a4412;
assign a4422 = ~l1242 & l1240;
assign a4424 = a4422 & ~l1238;
assign a4426 = a4424 & a4346;
assign a4428 = a4426 & a4364;
assign a4430 = a4412 & a4360;
assign a4432 = ~a4430 & ~l1194;
assign a4434 = a4432 & ~a4428;
assign a4436 = a4434 & ~a4420;
assign a4440 = l1208 & ~l1206;
assign a4442 = a4440 & a4342;
assign a4444 = ~l1208 & l1206;
assign a4446 = a4444 & a4342;
assign a4448 = a4444 & a4352;
assign a4450 = l1198 & ~l1196;
assign a4452 = a4444 & a4358;
assign a4454 = a4452 & a4450;
assign a4456 = ~l1198 & ~l1196;
assign a4458 = l1208 & l1206;
assign a4460 = a4458 & a4368;
assign a4462 = a4460 & a4456;
assign a4464 = a4440 & a4368;
assign a4466 = a4464 & a4450;
assign a4468 = ~a4378 & l1200;
assign a4470 = a4468 & ~a4466;
assign a4472 = a4470 & ~a4462;
assign a4474 = ~a4472 & ~a4454;
assign a4476 = ~a4474 & ~a4448;
assign a4478 = ~a4476 & ~a4446;
assign a4480 = ~a4478 & ~a4442;
assign a4484 = ~a4378 & l1202;
assign a4486 = a4484 & ~a4466;
assign a4488 = a4486 & ~a4462;
assign a4490 = ~a4488 & ~a4454;
assign a4492 = ~a4490 & ~a4448;
assign a4494 = ~a4492 & ~a4446;
assign a4496 = a4494 & ~a4442;
assign a4500 = ~l1198 & l1196;
assign a4502 = a4444 & a4416;
assign a4504 = a4502 & a4500;
assign a4506 = a4444 & a4424;
assign a4508 = a4506 & a4456;
assign a4510 = a4500 & a4452;
assign a4512 = ~a4510 & ~l1208;
assign a4514 = a4512 & ~a4508;
assign a4516 = a4514 & ~a4504;
assign a4520 = l1222 & ~l1220;
assign a4522 = a4520 & a4342;
assign a4524 = ~l1222 & l1220;
assign a4526 = a4524 & a4342;
assign a4528 = a4524 & a4352;
assign a4530 = l1212 & ~l1210;
assign a4532 = a4524 & a4358;
assign a4534 = a4532 & a4530;
assign a4536 = ~l1212 & ~l1210;
assign a4538 = l1222 & l1220;
assign a4540 = a4538 & a4368;
assign a4542 = a4540 & a4536;
assign a4544 = a4520 & a4368;
assign a4546 = a4544 & a4530;
assign a4548 = ~a4378 & l1214;
assign a4550 = a4548 & ~a4546;
assign a4552 = a4550 & ~a4542;
assign a4554 = ~a4552 & ~a4534;
assign a4556 = ~a4554 & ~a4528;
assign a4558 = ~a4556 & ~a4526;
assign a4560 = ~a4558 & ~a4522;
assign a4564 = ~a4378 & l1216;
assign a4566 = a4564 & ~a4546;
assign a4568 = a4566 & ~a4542;
assign a4570 = ~a4568 & ~a4534;
assign a4572 = ~a4570 & ~a4528;
assign a4574 = ~a4572 & ~a4526;
assign a4576 = a4574 & ~a4522;
assign a4580 = ~l1212 & l1210;
assign a4582 = a4524 & a4416;
assign a4584 = a4582 & a4580;
assign a4586 = a4524 & a4424;
assign a4588 = a4586 & a4536;
assign a4590 = a4580 & a4532;
assign a4592 = ~a4590 & ~l1222;
assign a4594 = a4592 & ~a4588;
assign a4596 = a4594 & ~a4584;
assign a4600 = l1236 & ~l1234;
assign a4602 = a4600 & a4342;
assign a4604 = ~l1236 & l1234;
assign a4606 = a4604 & a4342;
assign a4608 = a4604 & a4352;
assign a4610 = l1226 & ~l1224;
assign a4612 = a4604 & a4358;
assign a4614 = a4612 & a4610;
assign a4616 = ~l1226 & ~l1224;
assign a4618 = l1236 & l1234;
assign a4620 = a4618 & a4368;
assign a4622 = a4620 & a4616;
assign a4624 = a4600 & a4368;
assign a4626 = a4624 & a4610;
assign a4628 = ~a4378 & l1228;
assign a4630 = a4628 & ~a4626;
assign a4632 = a4630 & ~a4622;
assign a4634 = ~a4632 & ~a4614;
assign a4636 = ~a4634 & ~a4608;
assign a4638 = ~a4636 & ~a4606;
assign a4640 = ~a4638 & ~a4602;
assign a4644 = ~a4378 & l1230;
assign a4646 = a4644 & ~a4626;
assign a4648 = a4646 & ~a4622;
assign a4650 = ~a4648 & ~a4614;
assign a4652 = ~a4650 & ~a4608;
assign a4654 = ~a4652 & ~a4606;
assign a4656 = a4654 & ~a4602;
assign a4660 = ~l1226 & l1224;
assign a4662 = a4604 & a4416;
assign a4664 = a4662 & a4660;
assign a4666 = a4604 & a4424;
assign a4668 = a4666 & a4616;
assign a4670 = a4660 & a4612;
assign a4672 = ~a4670 & ~l1236;
assign a4674 = a4672 & ~a4668;
assign a4676 = a4674 & ~a4664;
assign a4680 = l1264 & l1262;
assign a4682 = ~a4680 & ~l1260;
assign a4684 = ~a4682 & l1258;
assign a4686 = ~a4684 & ~l1256;
assign a4688 = a4686 & l1250;
assign a4690 = ~a4444 & ~a4346;
assign a4692 = a4690 & ~a4524;
assign a4694 = a4444 & a4346;
assign a4696 = ~a4694 & ~a4524;
assign a4698 = ~a4696 & ~a4690;
assign a4700 = ~a4698 & ~a4604;
assign a4702 = ~a4700 & ~a4692;
assign a4704 = ~a4702 & a4416;
assign a4706 = a4704 & ~a4688;
assign a4708 = ~a4356 & a4338;
assign a4710 = ~a4708 & a4342;
assign a4712 = ~a4450 & a4440;
assign a4714 = ~a4712 & a4710;
assign a4716 = ~a4530 & a4520;
assign a4718 = ~a4716 & a4714;
assign a4720 = ~a4610 & a4600;
assign a4722 = ~a4720 & a4718;
assign a4724 = ~a4364 & a4346;
assign a4726 = ~a4724 & a4424;
assign a4728 = ~a4456 & a4444;
assign a4730 = ~a4728 & a4726;
assign a4732 = ~a4536 & a4524;
assign a4734 = ~a4732 & a4730;
assign a4736 = ~a4616 & a4604;
assign a4738 = ~a4736 & a4734;
assign a4740 = ~a4660 & a4604;
assign a4742 = ~a4580 & a4524;
assign a4744 = ~a4500 & a4444;
assign a4746 = ~a4412 & a4346;
assign a4748 = ~a4746 & a4424;
assign a4750 = a4748 & ~a4744;
assign a4752 = a4750 & ~a4742;
assign a4754 = a4752 & ~a4740;
assign a4756 = ~a4610 & a4604;
assign a4758 = ~a4530 & a4524;
assign a4760 = ~a4356 & a4346;
assign a4762 = ~a4450 & a4444;
assign a4764 = ~a4762 & ~a4760;
assign a4766 = a4764 & ~a4758;
assign a4768 = a4766 & ~a4756;
assign a4770 = ~a4746 & ~a4744;
assign a4772 = a4770 & ~a4742;
assign a4774 = a4772 & ~a4740;
assign a4776 = ~a4774 & ~a4768;
assign a4778 = ~a4776 & ~a4350;
assign a4780 = a4778 & a4358;
assign a4782 = a4780 & ~a4414;
assign a4784 = ~a4782 & l1238;
assign a4786 = ~a4784 & ~a4754;
assign a4788 = ~a4786 & ~a4738;
assign a4790 = a4788 & ~a4722;
assign a4792 = a4790 & ~a4706;
assign a4796 = a4352 & ~l1252;
assign a4798 = a4414 & l1238;
assign a4800 = l1242 & l1238;
assign a4802 = a4800 & l1252;
assign a4804 = ~a4802 & a4798;
assign a4806 = ~a4804 & ~l1240;
assign a4808 = a4806 & ~a4796;
assign a4810 = ~a4808 & ~a4754;
assign a4812 = a4810 & ~a4738;
assign a4814 = ~a4812 & ~a4722;
assign a4816 = a4814 & ~a4706;
assign a4820 = a4352 & l1252;
assign a4822 = ~a4758 & ~a4756;
assign a4824 = a4822 & ~a4762;
assign a4826 = a4824 & ~a4760;
assign a4828 = a4826 & a4358;
assign a4830 = ~a4828 & l1242;
assign a4832 = ~a4830 & ~a4798;
assign a4834 = ~a4832 & ~a4820;
assign a4836 = ~a4834 & ~a4796;
assign a4838 = a4836 & ~a4754;
assign a4840 = a4838 & ~a4738;
assign a4842 = ~a4840 & ~a4722;
assign a4844 = ~a4842 & ~a4706;
assign a4848 = ~l1262 & ~l1260;
assign a4850 = a4848 & ~l1258;
assign a4852 = ~a4850 & l1256;
assign a4854 = a4852 & a4416;
assign a4856 = ~a4854 & ~l1254;
assign a4860 = ~l1264 & ~l1262;
assign a4862 = a4860 & ~l1260;
assign a4864 = a4862 & ~l1258;
assign a4866 = a4864 & ~l1256;
assign a4868 = l1264 & ~l1262;
assign a4870 = a4868 & ~l1260;
assign a4872 = a4870 & ~l1258;
assign a4874 = a4872 & ~l1256;
assign a4876 = ~l1264 & l1262;
assign a4878 = a4876 & ~l1260;
assign a4880 = a4878 & ~l1258;
assign a4882 = a4880 & ~l1256;
assign a4884 = a4680 & ~l1260;
assign a4886 = a4884 & ~l1258;
assign a4888 = a4886 & ~l1256;
assign a4890 = a4860 & l1260;
assign a4892 = a4890 & ~l1258;
assign a4894 = a4892 & ~l1256;
assign a4896 = a4868 & l1260;
assign a4898 = a4896 & ~l1258;
assign a4900 = a4898 & ~l1256;
assign a4902 = a4876 & l1260;
assign a4904 = a4902 & ~l1258;
assign a4906 = a4904 & ~l1256;
assign a4908 = a4680 & l1260;
assign a4910 = a4908 & ~l1258;
assign a4912 = a4910 & ~l1256;
assign a4914 = l1258 & ~l1256;
assign a4916 = ~a4876 & a4682;
assign a4918 = a4916 & ~a4870;
assign a4920 = a4918 & ~a4862;
assign a4922 = ~a4920 & a4914;
assign a4924 = a4922 & ~a4912;
assign a4926 = a4924 & ~a4906;
assign a4928 = a4926 & ~a4900;
assign a4930 = a4928 & ~a4894;
assign a4932 = a4930 & ~a4888;
assign a4934 = a4932 & ~a4882;
assign a4936 = a4934 & ~a4874;
assign a4938 = a4936 & ~a4866;
assign a4940 = l1260 & ~l1256;
assign a4942 = a4680 & ~l1258;
assign a4944 = a4862 & l1258;
assign a4946 = a4944 & ~l1256;
assign a4948 = a4870 & l1258;
assign a4950 = a4948 & ~l1256;
assign a4952 = a4878 & l1258;
assign a4954 = a4952 & ~l1256;
assign a4956 = a4884 & l1258;
assign a4958 = a4956 & ~l1256;
assign a4960 = ~a4958 & l1258;
assign a4962 = a4960 & ~a4954;
assign a4964 = a4962 & ~a4950;
assign a4966 = a4964 & ~a4946;
assign a4968 = ~a4966 & ~a4942;
assign a4970 = a4876 & ~l1258;
assign a4972 = ~a4970 & a4968;
assign a4974 = a4868 & ~l1258;
assign a4976 = ~a4974 & a4972;
assign a4978 = a4860 & ~l1258;
assign a4980 = ~a4978 & a4976;
assign a4982 = ~a4980 & a4940;
assign a4984 = a4982 & ~a4888;
assign a4986 = a4984 & ~a4882;
assign a4988 = a4986 & ~a4874;
assign a4990 = a4988 & ~a4866;
assign a4992 = a4850 & ~l1256;
assign a4994 = l1262 & ~l1260;
assign a4996 = a4994 & ~l1258;
assign a4998 = a4996 & ~l1256;
assign a5000 = ~l1262 & l1260;
assign a5002 = a5000 & ~l1258;
assign a5004 = a5002 & ~l1256;
assign a5006 = l1262 & l1260;
assign a5008 = a5006 & ~l1258;
assign a5010 = a5008 & ~l1256;
assign a5012 = a4848 & l1258;
assign a5014 = a5012 & ~l1256;
assign a5016 = a4994 & l1258;
assign a5018 = a5016 & ~l1256;
assign a5020 = a4890 & l1258;
assign a5022 = a5020 & ~l1256;
assign a5024 = a5000 & l1258;
assign a5026 = a5024 & ~l1256;
assign a5028 = a4902 & l1258;
assign a5030 = a5028 & ~l1256;
assign a5032 = a5006 & l1258;
assign a5034 = a5032 & ~l1256;
assign a5036 = a4850 & l1256;
assign a5038 = a5036 & ~a4864;
assign a5040 = ~a5038 & ~a5034;
assign a5042 = ~a5040 & ~a5030;
assign a5044 = ~a5042 & ~a5026;
assign a5046 = ~a5044 & ~a5022;
assign a5048 = ~a5046 & ~a5018;
assign a5050 = ~a5048 & ~a4954;
assign a5052 = ~a5050 & ~a5014;
assign a5054 = ~a5052 & ~a4946;
assign a5056 = ~a5054 & ~a5010;
assign a5058 = ~a5056 & ~a4906;
assign a5060 = ~a5058 & ~a5004;
assign a5062 = ~a5060 & ~a4894;
assign a5064 = ~a5062 & ~a4998;
assign a5066 = ~a5064 & ~a4882;
assign a5068 = ~a5066 & ~a4992;
assign a5070 = ~a5068 & l1264;
assign a5072 = a5070 & ~a4866;
assign a5074 = l1264 & ~l1260;
assign a5076 = a5074 & ~l1258;
assign a5078 = a5076 & ~l1256;
assign a5080 = l1264 & l1260;
assign a5082 = a5080 & ~l1258;
assign a5084 = a5082 & ~l1256;
assign a5086 = a5074 & l1258;
assign a5088 = a5086 & ~l1256;
assign a5090 = a5080 & l1258;
assign a5092 = a5090 & ~l1256;
assign a5094 = ~l1260 & ~l1258;
assign a5096 = a5094 & l1256;
assign a5098 = ~a5096 & ~a5092;
assign a5100 = ~l1264 & l1260;
assign a5102 = a5100 & l1258;
assign a5104 = a5102 & ~l1256;
assign a5106 = ~a5104 & a5098;
assign a5108 = ~a5106 & ~a4958;
assign a5110 = a5108 & ~a4954;
assign a5112 = ~a5110 & ~a5088;
assign a5114 = ~l1264 & ~l1260;
assign a5116 = a5114 & l1258;
assign a5118 = a5116 & ~l1256;
assign a5120 = ~a5118 & a5112;
assign a5122 = ~a5120 & ~a4912;
assign a5124 = a5122 & ~a4906;
assign a5126 = ~a5124 & ~a5084;
assign a5128 = a5100 & ~l1258;
assign a5130 = a5128 & ~l1256;
assign a5132 = ~a5130 & a5126;
assign a5134 = ~a5132 & ~a4888;
assign a5136 = a5134 & ~a4882;
assign a5138 = ~a5136 & ~a5078;
assign a5140 = a5114 & ~l1258;
assign a5142 = a5140 & ~l1256;
assign a5144 = ~a5142 & a5138;
assign a5146 = ~a5144 & ~l1262;
assign a5148 = ~a5146 & a5072;
assign a5150 = a5148 & ~a4990;
assign a5152 = a5150 & ~a4938;
assign a5154 = ~a4920 & l1258;
assign a5156 = ~a5154 & ~a4910;
assign a5158 = a5156 & ~a4904;
assign a5160 = a5158 & ~a4898;
assign a5162 = a5160 & ~a4892;
assign a5164 = a5162 & ~a4886;
assign a5166 = a5164 & ~a4880;
assign a5168 = a5166 & ~a4872;
assign a5170 = a5168 & ~a4864;
assign a5172 = ~a5170 & ~l1256;
assign a5174 = ~a5172 & a5152;
assign a5176 = ~a5174 & l1256;
assign a5178 = ~a5176 & a4416;
assign a5180 = ~a4416 & ~l1256;
assign a5182 = ~a5180 & ~a5178;
assign a5186 = ~a5174 & l1258;
assign a5188 = ~a5186 & a4416;
assign a5190 = ~a4416 & ~l1258;
assign a5192 = ~a5190 & ~a5188;
assign a5196 = ~a5174 & l1260;
assign a5198 = ~a5196 & a4416;
assign a5200 = ~a4416 & ~l1260;
assign a5202 = ~a5200 & ~a5198;
assign a5206 = ~a5174 & l1262;
assign a5208 = ~a5206 & a4416;
assign a5210 = ~a4416 & ~l1262;
assign a5212 = ~a5210 & ~a5208;
assign a5216 = a4416 & l1264;
assign a5218 = ~a4416 & ~l1264;
assign a5220 = ~a5218 & ~a5216;
assign a5224 = l1278 & ~l1276;
assign a5226 = l1326 & l1324;
assign a5228 = a5226 & ~l1322;
assign a5230 = a5228 & a5224;
assign a5232 = ~l1278 & l1276;
assign a5234 = a5232 & a5228;
assign a5236 = l1326 & ~l1324;
assign a5238 = a5236 & l1322;
assign a5240 = a5238 & a5232;
assign a5242 = l1268 & ~l1266;
assign a5244 = a5226 & l1322;
assign a5246 = a5244 & a5232;
assign a5248 = a5246 & a5242;
assign a5250 = ~l1268 & ~l1266;
assign a5252 = l1278 & l1276;
assign a5254 = a5236 & ~l1322;
assign a5256 = a5254 & a5252;
assign a5258 = a5256 & a5250;
assign a5260 = a5254 & a5224;
assign a5262 = a5260 & a5242;
assign a5264 = a5254 & l1328;
assign a5266 = ~a5264 & l1270;
assign a5268 = a5266 & ~a5262;
assign a5270 = a5268 & ~a5258;
assign a5272 = ~a5270 & ~a5248;
assign a5274 = ~a5272 & ~a5240;
assign a5276 = ~a5274 & ~a5234;
assign a5278 = ~a5276 & ~a5230;
assign a5282 = ~a5264 & l1272;
assign a5284 = a5282 & ~a5262;
assign a5286 = a5284 & ~a5258;
assign a5288 = ~a5286 & ~a5248;
assign a5290 = ~a5288 & ~a5240;
assign a5292 = ~a5290 & ~a5234;
assign a5294 = a5292 & ~a5230;
assign a5298 = ~l1268 & l1266;
assign a5300 = ~l1326 & ~l1324;
assign a5302 = a5300 & ~l1322;
assign a5304 = a5302 & a5232;
assign a5306 = a5304 & a5298;
assign a5308 = ~l1326 & l1324;
assign a5310 = a5308 & ~l1322;
assign a5312 = a5310 & a5232;
assign a5314 = a5312 & a5250;
assign a5316 = a5298 & a5246;
assign a5318 = ~a5316 & ~l1278;
assign a5320 = a5318 & ~a5314;
assign a5322 = a5320 & ~a5306;
assign a5326 = l1292 & ~l1290;
assign a5328 = a5326 & a5228;
assign a5330 = ~l1292 & l1290;
assign a5332 = a5330 & a5228;
assign a5334 = a5330 & a5238;
assign a5336 = l1282 & ~l1280;
assign a5338 = a5330 & a5244;
assign a5340 = a5338 & a5336;
assign a5342 = ~l1282 & ~l1280;
assign a5344 = l1292 & l1290;
assign a5346 = a5344 & a5254;
assign a5348 = a5346 & a5342;
assign a5350 = a5326 & a5254;
assign a5352 = a5350 & a5336;
assign a5354 = ~a5264 & l1284;
assign a5356 = a5354 & ~a5352;
assign a5358 = a5356 & ~a5348;
assign a5360 = ~a5358 & ~a5340;
assign a5362 = ~a5360 & ~a5334;
assign a5364 = ~a5362 & ~a5332;
assign a5366 = ~a5364 & ~a5328;
assign a5370 = ~a5264 & l1286;
assign a5372 = a5370 & ~a5352;
assign a5374 = a5372 & ~a5348;
assign a5376 = ~a5374 & ~a5340;
assign a5378 = ~a5376 & ~a5334;
assign a5380 = ~a5378 & ~a5332;
assign a5382 = a5380 & ~a5328;
assign a5386 = ~l1282 & l1280;
assign a5388 = a5330 & a5302;
assign a5390 = a5388 & a5386;
assign a5392 = a5330 & a5310;
assign a5394 = a5392 & a5342;
assign a5396 = a5386 & a5338;
assign a5398 = ~a5396 & ~l1292;
assign a5400 = a5398 & ~a5394;
assign a5402 = a5400 & ~a5390;
assign a5406 = l1306 & ~l1304;
assign a5408 = a5406 & a5228;
assign a5410 = ~l1306 & l1304;
assign a5412 = a5410 & a5228;
assign a5414 = a5410 & a5238;
assign a5416 = l1296 & ~l1294;
assign a5418 = a5410 & a5244;
assign a5420 = a5418 & a5416;
assign a5422 = ~l1296 & ~l1294;
assign a5424 = l1306 & l1304;
assign a5426 = a5424 & a5254;
assign a5428 = a5426 & a5422;
assign a5430 = a5406 & a5254;
assign a5432 = a5430 & a5416;
assign a5434 = ~a5264 & l1298;
assign a5436 = a5434 & ~a5432;
assign a5438 = a5436 & ~a5428;
assign a5440 = ~a5438 & ~a5420;
assign a5442 = ~a5440 & ~a5414;
assign a5444 = ~a5442 & ~a5412;
assign a5446 = ~a5444 & ~a5408;
assign a5450 = ~a5264 & l1300;
assign a5452 = a5450 & ~a5432;
assign a5454 = a5452 & ~a5428;
assign a5456 = ~a5454 & ~a5420;
assign a5458 = ~a5456 & ~a5414;
assign a5460 = ~a5458 & ~a5412;
assign a5462 = a5460 & ~a5408;
assign a5466 = ~l1296 & l1294;
assign a5468 = a5410 & a5302;
assign a5470 = a5468 & a5466;
assign a5472 = a5410 & a5310;
assign a5474 = a5472 & a5422;
assign a5476 = a5466 & a5418;
assign a5478 = ~a5476 & ~l1306;
assign a5480 = a5478 & ~a5474;
assign a5482 = a5480 & ~a5470;
assign a5486 = l1320 & ~l1318;
assign a5488 = a5486 & a5228;
assign a5490 = ~l1320 & l1318;
assign a5492 = a5490 & a5228;
assign a5494 = a5490 & a5238;
assign a5496 = l1310 & ~l1308;
assign a5498 = a5490 & a5244;
assign a5500 = a5498 & a5496;
assign a5502 = ~l1310 & ~l1308;
assign a5504 = l1320 & l1318;
assign a5506 = a5504 & a5254;
assign a5508 = a5506 & a5502;
assign a5510 = a5486 & a5254;
assign a5512 = a5510 & a5496;
assign a5514 = ~a5264 & l1312;
assign a5516 = a5514 & ~a5512;
assign a5518 = a5516 & ~a5508;
assign a5520 = ~a5518 & ~a5500;
assign a5522 = ~a5520 & ~a5494;
assign a5524 = ~a5522 & ~a5492;
assign a5526 = ~a5524 & ~a5488;
assign a5530 = ~a5264 & l1314;
assign a5532 = a5530 & ~a5512;
assign a5534 = a5532 & ~a5508;
assign a5536 = ~a5534 & ~a5500;
assign a5538 = ~a5536 & ~a5494;
assign a5540 = ~a5538 & ~a5492;
assign a5542 = a5540 & ~a5488;
assign a5546 = ~l1310 & l1308;
assign a5548 = a5490 & a5302;
assign a5550 = a5548 & a5546;
assign a5552 = a5490 & a5310;
assign a5554 = a5552 & a5502;
assign a5556 = a5546 & a5498;
assign a5558 = ~a5556 & ~l1320;
assign a5560 = a5558 & ~a5554;
assign a5562 = a5560 & ~a5550;
assign a5566 = l1348 & l1346;
assign a5568 = ~a5566 & ~l1344;
assign a5570 = ~a5568 & l1342;
assign a5572 = ~a5570 & ~l1340;
assign a5574 = a5572 & l1334;
assign a5576 = ~a5330 & ~a5232;
assign a5578 = a5576 & ~a5410;
assign a5580 = a5330 & a5232;
assign a5582 = ~a5580 & ~a5410;
assign a5584 = ~a5582 & ~a5576;
assign a5586 = ~a5584 & ~a5490;
assign a5588 = ~a5586 & ~a5578;
assign a5590 = ~a5588 & a5302;
assign a5592 = a5590 & ~a5574;
assign a5594 = ~a5242 & a5224;
assign a5596 = ~a5594 & a5228;
assign a5598 = ~a5336 & a5326;
assign a5600 = ~a5598 & a5596;
assign a5602 = ~a5416 & a5406;
assign a5604 = ~a5602 & a5600;
assign a5606 = ~a5496 & a5486;
assign a5608 = ~a5606 & a5604;
assign a5610 = ~a5250 & a5232;
assign a5612 = ~a5610 & a5310;
assign a5614 = ~a5342 & a5330;
assign a5616 = ~a5614 & a5612;
assign a5618 = ~a5422 & a5410;
assign a5620 = ~a5618 & a5616;
assign a5622 = ~a5502 & a5490;
assign a5624 = ~a5622 & a5620;
assign a5626 = ~a5546 & a5490;
assign a5628 = ~a5466 & a5410;
assign a5630 = ~a5386 & a5330;
assign a5632 = ~a5298 & a5232;
assign a5634 = ~a5632 & a5310;
assign a5636 = a5634 & ~a5630;
assign a5638 = a5636 & ~a5628;
assign a5640 = a5638 & ~a5626;
assign a5642 = ~a5496 & a5490;
assign a5644 = ~a5416 & a5410;
assign a5646 = ~a5242 & a5232;
assign a5648 = ~a5336 & a5330;
assign a5650 = ~a5648 & ~a5646;
assign a5652 = a5650 & ~a5644;
assign a5654 = a5652 & ~a5642;
assign a5656 = ~a5632 & ~a5630;
assign a5658 = a5656 & ~a5628;
assign a5660 = a5658 & ~a5626;
assign a5662 = ~a5660 & ~a5654;
assign a5664 = ~a5662 & ~a5236;
assign a5666 = a5664 & a5244;
assign a5668 = a5666 & ~a5300;
assign a5670 = ~a5668 & l1322;
assign a5672 = ~a5670 & ~a5640;
assign a5674 = ~a5672 & ~a5624;
assign a5676 = a5674 & ~a5608;
assign a5678 = a5676 & ~a5592;
assign a5682 = a5238 & ~l1336;
assign a5684 = a5300 & l1322;
assign a5686 = l1326 & l1322;
assign a5688 = a5686 & l1336;
assign a5690 = ~a5688 & a5684;
assign a5692 = ~a5690 & ~l1324;
assign a5694 = a5692 & ~a5682;
assign a5696 = ~a5694 & ~a5640;
assign a5698 = a5696 & ~a5624;
assign a5700 = ~a5698 & ~a5608;
assign a5702 = a5700 & ~a5592;
assign a5706 = a5238 & l1336;
assign a5708 = ~a5644 & ~a5642;
assign a5710 = a5708 & ~a5648;
assign a5712 = a5710 & ~a5646;
assign a5714 = a5712 & a5244;
assign a5716 = ~a5714 & l1326;
assign a5718 = ~a5716 & ~a5684;
assign a5720 = ~a5718 & ~a5706;
assign a5722 = ~a5720 & ~a5682;
assign a5724 = a5722 & ~a5640;
assign a5726 = a5724 & ~a5624;
assign a5728 = ~a5726 & ~a5608;
assign a5730 = ~a5728 & ~a5592;
assign a5734 = ~l1346 & ~l1344;
assign a5736 = a5734 & ~l1342;
assign a5738 = ~a5736 & l1340;
assign a5740 = a5738 & a5302;
assign a5742 = ~a5740 & ~l1338;
assign a5746 = ~l1348 & ~l1346;
assign a5748 = a5746 & ~l1344;
assign a5750 = a5748 & ~l1342;
assign a5752 = a5750 & ~l1340;
assign a5754 = l1348 & ~l1346;
assign a5756 = a5754 & ~l1344;
assign a5758 = a5756 & ~l1342;
assign a5760 = a5758 & ~l1340;
assign a5762 = ~l1348 & l1346;
assign a5764 = a5762 & ~l1344;
assign a5766 = a5764 & ~l1342;
assign a5768 = a5766 & ~l1340;
assign a5770 = a5566 & ~l1344;
assign a5772 = a5770 & ~l1342;
assign a5774 = a5772 & ~l1340;
assign a5776 = a5746 & l1344;
assign a5778 = a5776 & ~l1342;
assign a5780 = a5778 & ~l1340;
assign a5782 = a5754 & l1344;
assign a5784 = a5782 & ~l1342;
assign a5786 = a5784 & ~l1340;
assign a5788 = a5762 & l1344;
assign a5790 = a5788 & ~l1342;
assign a5792 = a5790 & ~l1340;
assign a5794 = a5566 & l1344;
assign a5796 = a5794 & ~l1342;
assign a5798 = a5796 & ~l1340;
assign a5800 = l1342 & ~l1340;
assign a5802 = ~a5762 & a5568;
assign a5804 = a5802 & ~a5756;
assign a5806 = a5804 & ~a5748;
assign a5808 = ~a5806 & a5800;
assign a5810 = a5808 & ~a5798;
assign a5812 = a5810 & ~a5792;
assign a5814 = a5812 & ~a5786;
assign a5816 = a5814 & ~a5780;
assign a5818 = a5816 & ~a5774;
assign a5820 = a5818 & ~a5768;
assign a5822 = a5820 & ~a5760;
assign a5824 = a5822 & ~a5752;
assign a5826 = l1344 & ~l1340;
assign a5828 = a5566 & ~l1342;
assign a5830 = a5748 & l1342;
assign a5832 = a5830 & ~l1340;
assign a5834 = a5756 & l1342;
assign a5836 = a5834 & ~l1340;
assign a5838 = a5764 & l1342;
assign a5840 = a5838 & ~l1340;
assign a5842 = a5770 & l1342;
assign a5844 = a5842 & ~l1340;
assign a5846 = ~a5844 & l1342;
assign a5848 = a5846 & ~a5840;
assign a5850 = a5848 & ~a5836;
assign a5852 = a5850 & ~a5832;
assign a5854 = ~a5852 & ~a5828;
assign a5856 = a5762 & ~l1342;
assign a5858 = ~a5856 & a5854;
assign a5860 = a5754 & ~l1342;
assign a5862 = ~a5860 & a5858;
assign a5864 = a5746 & ~l1342;
assign a5866 = ~a5864 & a5862;
assign a5868 = ~a5866 & a5826;
assign a5870 = a5868 & ~a5774;
assign a5872 = a5870 & ~a5768;
assign a5874 = a5872 & ~a5760;
assign a5876 = a5874 & ~a5752;
assign a5878 = a5736 & ~l1340;
assign a5880 = l1346 & ~l1344;
assign a5882 = a5880 & ~l1342;
assign a5884 = a5882 & ~l1340;
assign a5886 = ~l1346 & l1344;
assign a5888 = a5886 & ~l1342;
assign a5890 = a5888 & ~l1340;
assign a5892 = l1346 & l1344;
assign a5894 = a5892 & ~l1342;
assign a5896 = a5894 & ~l1340;
assign a5898 = a5734 & l1342;
assign a5900 = a5898 & ~l1340;
assign a5902 = a5880 & l1342;
assign a5904 = a5902 & ~l1340;
assign a5906 = a5776 & l1342;
assign a5908 = a5906 & ~l1340;
assign a5910 = a5886 & l1342;
assign a5912 = a5910 & ~l1340;
assign a5914 = a5788 & l1342;
assign a5916 = a5914 & ~l1340;
assign a5918 = a5892 & l1342;
assign a5920 = a5918 & ~l1340;
assign a5922 = a5736 & l1340;
assign a5924 = a5922 & ~a5750;
assign a5926 = ~a5924 & ~a5920;
assign a5928 = ~a5926 & ~a5916;
assign a5930 = ~a5928 & ~a5912;
assign a5932 = ~a5930 & ~a5908;
assign a5934 = ~a5932 & ~a5904;
assign a5936 = ~a5934 & ~a5840;
assign a5938 = ~a5936 & ~a5900;
assign a5940 = ~a5938 & ~a5832;
assign a5942 = ~a5940 & ~a5896;
assign a5944 = ~a5942 & ~a5792;
assign a5946 = ~a5944 & ~a5890;
assign a5948 = ~a5946 & ~a5780;
assign a5950 = ~a5948 & ~a5884;
assign a5952 = ~a5950 & ~a5768;
assign a5954 = ~a5952 & ~a5878;
assign a5956 = ~a5954 & l1348;
assign a5958 = a5956 & ~a5752;
assign a5960 = l1348 & ~l1344;
assign a5962 = a5960 & ~l1342;
assign a5964 = a5962 & ~l1340;
assign a5966 = l1348 & l1344;
assign a5968 = a5966 & ~l1342;
assign a5970 = a5968 & ~l1340;
assign a5972 = a5960 & l1342;
assign a5974 = a5972 & ~l1340;
assign a5976 = a5966 & l1342;
assign a5978 = a5976 & ~l1340;
assign a5980 = ~l1344 & ~l1342;
assign a5982 = a5980 & l1340;
assign a5984 = ~a5982 & ~a5978;
assign a5986 = ~l1348 & l1344;
assign a5988 = a5986 & l1342;
assign a5990 = a5988 & ~l1340;
assign a5992 = ~a5990 & a5984;
assign a5994 = ~a5992 & ~a5844;
assign a5996 = a5994 & ~a5840;
assign a5998 = ~a5996 & ~a5974;
assign a6000 = ~l1348 & ~l1344;
assign a6002 = a6000 & l1342;
assign a6004 = a6002 & ~l1340;
assign a6006 = ~a6004 & a5998;
assign a6008 = ~a6006 & ~a5798;
assign a6010 = a6008 & ~a5792;
assign a6012 = ~a6010 & ~a5970;
assign a6014 = a5986 & ~l1342;
assign a6016 = a6014 & ~l1340;
assign a6018 = ~a6016 & a6012;
assign a6020 = ~a6018 & ~a5774;
assign a6022 = a6020 & ~a5768;
assign a6024 = ~a6022 & ~a5964;
assign a6026 = a6000 & ~l1342;
assign a6028 = a6026 & ~l1340;
assign a6030 = ~a6028 & a6024;
assign a6032 = ~a6030 & ~l1346;
assign a6034 = ~a6032 & a5958;
assign a6036 = a6034 & ~a5876;
assign a6038 = a6036 & ~a5824;
assign a6040 = ~a5806 & l1342;
assign a6042 = ~a6040 & ~a5796;
assign a6044 = a6042 & ~a5790;
assign a6046 = a6044 & ~a5784;
assign a6048 = a6046 & ~a5778;
assign a6050 = a6048 & ~a5772;
assign a6052 = a6050 & ~a5766;
assign a6054 = a6052 & ~a5758;
assign a6056 = a6054 & ~a5750;
assign a6058 = ~a6056 & ~l1340;
assign a6060 = ~a6058 & a6038;
assign a6062 = ~a6060 & l1340;
assign a6064 = ~a6062 & a5302;
assign a6066 = ~a5302 & ~l1340;
assign a6068 = ~a6066 & ~a6064;
assign a6072 = ~a6060 & l1342;
assign a6074 = ~a6072 & a5302;
assign a6076 = ~a5302 & ~l1342;
assign a6078 = ~a6076 & ~a6074;
assign a6082 = ~a6060 & l1344;
assign a6084 = ~a6082 & a5302;
assign a6086 = ~a5302 & ~l1344;
assign a6088 = ~a6086 & ~a6084;
assign a6092 = ~a6060 & l1346;
assign a6094 = ~a6092 & a5302;
assign a6096 = ~a5302 & ~l1346;
assign a6098 = ~a6096 & ~a6094;
assign a6102 = a5302 & l1348;
assign a6104 = ~a5302 & ~l1348;
assign a6106 = ~a6104 & ~a6102;
assign a6110 = ~a3026 & l1352;
assign a6112 = ~a6110 & ~a2140;
assign a6116 = ~l1664 & ~l1662;
assign a6118 = ~a6116 & l1350;
assign a6120 = ~a6118 & ~l1656;
assign a6124 = ~l1354 & l1076;
assign a6126 = ~a6124 & l1356;
assign a6128 = ~a6126 & ~a6116;
assign a6130 = ~a6128 & ~l1658;
assign a6134 = l1354 & l1076;
assign a6136 = ~a6134 & ~a6116;
assign a6138 = ~a6136 & ~l1660;
assign a6144 = ~l1354 & ~l1076;
assign a6146 = l1350 & ~i412;
assign a6148 = a6124 & ~l1356;
assign a6150 = ~a6148 & ~a6146;
assign a6152 = a6150 & ~a6144;
assign a6154 = l730 & ~i2;
assign a6156 = ~l730 & i2;
assign a6158 = ~a6156 & ~a6154;
assign a6160 = a6158 & a6152;
assign a6162 = l732 & ~i4;
assign a6164 = ~l732 & i4;
assign a6166 = ~a6164 & ~a6162;
assign a6168 = a6166 & a6160;
assign a6170 = l734 & ~i6;
assign a6172 = ~l734 & i6;
assign a6174 = ~a6172 & ~a6170;
assign a6176 = a6174 & a6168;
assign a6178 = l736 & ~i8;
assign a6180 = ~l736 & i8;
assign a6182 = ~a6180 & ~a6178;
assign a6184 = a6182 & a6176;
assign a6186 = l738 & ~i10;
assign a6188 = ~l738 & i10;
assign a6190 = ~a6188 & ~a6186;
assign a6192 = a6190 & a6184;
assign a6194 = l740 & ~i12;
assign a6196 = ~l740 & i12;
assign a6198 = ~a6196 & ~a6194;
assign a6200 = a6198 & a6192;
assign a6202 = l742 & ~i14;
assign a6204 = ~l742 & i14;
assign a6206 = ~a6204 & ~a6202;
assign a6208 = a6206 & a6200;
assign a6210 = l744 & ~i16;
assign a6212 = ~l744 & i16;
assign a6214 = ~a6212 & ~a6210;
assign a6216 = a6214 & a6208;
assign a6218 = l746 & ~i18;
assign a6220 = ~l746 & i18;
assign a6222 = ~a6220 & ~a6218;
assign a6224 = a6222 & a6216;
assign a6226 = l748 & ~i20;
assign a6228 = ~l748 & i20;
assign a6230 = ~a6228 & ~a6226;
assign a6232 = a6230 & a6224;
assign a6234 = l750 & ~i22;
assign a6236 = ~l750 & i22;
assign a6238 = ~a6236 & ~a6234;
assign a6240 = a6238 & a6232;
assign a6242 = l752 & ~i24;
assign a6244 = ~l752 & i24;
assign a6246 = ~a6244 & ~a6242;
assign a6248 = a6246 & a6240;
assign a6250 = l754 & ~i26;
assign a6252 = ~l754 & i26;
assign a6254 = ~a6252 & ~a6250;
assign a6256 = a6254 & a6248;
assign a6258 = l756 & ~i28;
assign a6260 = ~l756 & i28;
assign a6262 = ~a6260 & ~a6258;
assign a6264 = a6262 & a6256;
assign a6266 = l758 & ~i30;
assign a6268 = ~l758 & i30;
assign a6270 = ~a6268 & ~a6266;
assign a6272 = a6270 & a6264;
assign a6274 = l760 & ~i32;
assign a6276 = ~l760 & i32;
assign a6278 = ~a6276 & ~a6274;
assign a6280 = a6278 & a6272;
assign a6282 = l762 & ~i34;
assign a6284 = ~l762 & i34;
assign a6286 = ~a6284 & ~a6282;
assign a6288 = a6286 & a6280;
assign a6290 = l764 & ~i36;
assign a6292 = ~l764 & i36;
assign a6294 = ~a6292 & ~a6290;
assign a6296 = a6294 & a6288;
assign a6298 = l766 & ~i38;
assign a6300 = ~l766 & i38;
assign a6302 = ~a6300 & ~a6298;
assign a6304 = a6302 & a6296;
assign a6306 = l768 & ~i40;
assign a6308 = ~l768 & i40;
assign a6310 = ~a6308 & ~a6306;
assign a6312 = a6310 & a6304;
assign a6314 = l770 & ~i42;
assign a6316 = ~l770 & i42;
assign a6318 = ~a6316 & ~a6314;
assign a6320 = a6318 & a6312;
assign a6322 = l772 & ~i44;
assign a6324 = ~l772 & i44;
assign a6326 = ~a6324 & ~a6322;
assign a6328 = a6326 & a6320;
assign a6330 = l774 & ~i46;
assign a6332 = ~l774 & i46;
assign a6334 = ~a6332 & ~a6330;
assign a6336 = a6334 & a6328;
assign a6338 = l776 & ~i48;
assign a6340 = ~l776 & i48;
assign a6342 = ~a6340 & ~a6338;
assign a6344 = a6342 & a6336;
assign a6346 = l778 & ~i50;
assign a6348 = ~l778 & i50;
assign a6350 = ~a6348 & ~a6346;
assign a6352 = a6350 & a6344;
assign a6354 = l780 & ~i52;
assign a6356 = ~l780 & i52;
assign a6358 = ~a6356 & ~a6354;
assign a6360 = a6358 & a6352;
assign a6362 = l782 & ~i54;
assign a6364 = ~l782 & i54;
assign a6366 = ~a6364 & ~a6362;
assign a6368 = a6366 & a6360;
assign a6370 = l784 & ~i56;
assign a6372 = ~l784 & i56;
assign a6374 = ~a6372 & ~a6370;
assign a6376 = a6374 & a6368;
assign a6378 = l786 & ~i58;
assign a6380 = ~l786 & i58;
assign a6382 = ~a6380 & ~a6378;
assign a6384 = a6382 & a6376;
assign a6386 = l788 & ~i60;
assign a6388 = ~l788 & i60;
assign a6390 = ~a6388 & ~a6386;
assign a6392 = a6390 & a6384;
assign a6394 = l790 & ~i62;
assign a6396 = ~l790 & i62;
assign a6398 = ~a6396 & ~a6394;
assign a6400 = a6398 & a6392;
assign a6402 = l792 & ~i64;
assign a6404 = ~l792 & i64;
assign a6406 = ~a6404 & ~a6402;
assign a6408 = a6406 & a6400;
assign a6410 = l794 & ~i66;
assign a6412 = ~l794 & i66;
assign a6414 = ~a6412 & ~a6410;
assign a6416 = a6414 & a6408;
assign a6418 = l796 & ~i68;
assign a6420 = ~l796 & i68;
assign a6422 = ~a6420 & ~a6418;
assign a6424 = a6422 & a6416;
assign a6426 = l798 & ~i70;
assign a6428 = ~l798 & i70;
assign a6430 = ~a6428 & ~a6426;
assign a6432 = a6430 & a6424;
assign a6434 = l800 & ~i72;
assign a6436 = ~l800 & i72;
assign a6438 = ~a6436 & ~a6434;
assign a6440 = a6438 & a6432;
assign a6442 = l802 & ~i74;
assign a6444 = ~l802 & i74;
assign a6446 = ~a6444 & ~a6442;
assign a6448 = a6446 & a6440;
assign a6450 = l804 & ~i76;
assign a6452 = ~l804 & i76;
assign a6454 = ~a6452 & ~a6450;
assign a6456 = a6454 & a6448;
assign a6458 = l806 & ~i78;
assign a6460 = ~l806 & i78;
assign a6462 = ~a6460 & ~a6458;
assign a6464 = a6462 & a6456;
assign a6466 = l808 & ~i80;
assign a6468 = ~l808 & i80;
assign a6470 = ~a6468 & ~a6466;
assign a6472 = a6470 & a6464;
assign a6474 = l810 & ~i82;
assign a6476 = ~l810 & i82;
assign a6478 = ~a6476 & ~a6474;
assign a6480 = a6478 & a6472;
assign a6482 = l812 & ~i84;
assign a6484 = ~l812 & i84;
assign a6486 = ~a6484 & ~a6482;
assign a6488 = a6486 & a6480;
assign a6490 = l814 & ~i86;
assign a6492 = ~l814 & i86;
assign a6494 = ~a6492 & ~a6490;
assign a6496 = a6494 & a6488;
assign a6498 = l816 & ~i88;
assign a6500 = ~l816 & i88;
assign a6502 = ~a6500 & ~a6498;
assign a6504 = a6502 & a6496;
assign a6506 = l818 & ~i90;
assign a6508 = ~l818 & i90;
assign a6510 = ~a6508 & ~a6506;
assign a6512 = a6510 & a6504;
assign a6514 = l820 & ~i92;
assign a6516 = ~l820 & i92;
assign a6518 = ~a6516 & ~a6514;
assign a6520 = a6518 & a6512;
assign a6522 = l822 & ~i94;
assign a6524 = ~l822 & i94;
assign a6526 = ~a6524 & ~a6522;
assign a6528 = a6526 & a6520;
assign a6530 = l824 & ~i96;
assign a6532 = ~l824 & i96;
assign a6534 = ~a6532 & ~a6530;
assign a6536 = a6534 & a6528;
assign a6538 = l826 & ~i98;
assign a6540 = ~l826 & i98;
assign a6542 = ~a6540 & ~a6538;
assign a6544 = a6542 & a6536;
assign a6546 = l828 & ~i100;
assign a6548 = ~l828 & i100;
assign a6550 = ~a6548 & ~a6546;
assign a6552 = a6550 & a6544;
assign a6554 = l830 & ~i102;
assign a6556 = ~l830 & i102;
assign a6558 = ~a6556 & ~a6554;
assign a6560 = a6558 & a6552;
assign a6562 = l832 & ~i104;
assign a6564 = ~l832 & i104;
assign a6566 = ~a6564 & ~a6562;
assign a6568 = a6566 & a6560;
assign a6570 = l834 & ~i106;
assign a6572 = ~l834 & i106;
assign a6574 = ~a6572 & ~a6570;
assign a6576 = a6574 & a6568;
assign a6578 = l836 & ~i108;
assign a6580 = ~l836 & i108;
assign a6582 = ~a6580 & ~a6578;
assign a6584 = a6582 & a6576;
assign a6586 = l838 & ~i110;
assign a6588 = ~l838 & i110;
assign a6590 = ~a6588 & ~a6586;
assign a6592 = a6590 & a6584;
assign a6594 = l840 & ~i112;
assign a6596 = ~l840 & i112;
assign a6598 = ~a6596 & ~a6594;
assign a6600 = a6598 & a6592;
assign a6602 = l842 & ~i114;
assign a6604 = ~l842 & i114;
assign a6606 = ~a6604 & ~a6602;
assign a6608 = a6606 & a6600;
assign a6610 = l844 & ~i116;
assign a6612 = ~l844 & i116;
assign a6614 = ~a6612 & ~a6610;
assign a6616 = a6614 & a6608;
assign a6618 = l846 & ~i118;
assign a6620 = ~l846 & i118;
assign a6622 = ~a6620 & ~a6618;
assign a6624 = a6622 & a6616;
assign a6626 = l848 & ~i120;
assign a6628 = ~l848 & i120;
assign a6630 = ~a6628 & ~a6626;
assign a6632 = a6630 & a6624;
assign a6634 = l850 & ~i122;
assign a6636 = ~l850 & i122;
assign a6638 = ~a6636 & ~a6634;
assign a6640 = a6638 & a6632;
assign a6642 = l852 & ~i124;
assign a6644 = ~l852 & i124;
assign a6646 = ~a6644 & ~a6642;
assign a6648 = a6646 & a6640;
assign a6650 = l854 & ~i126;
assign a6652 = ~l854 & i126;
assign a6654 = ~a6652 & ~a6650;
assign a6656 = a6654 & a6648;
assign a6658 = l856 & ~i128;
assign a6660 = ~l856 & i128;
assign a6662 = ~a6660 & ~a6658;
assign a6664 = a6662 & a6656;
assign a6666 = l858 & ~i130;
assign a6668 = ~l858 & i130;
assign a6670 = ~a6668 & ~a6666;
assign a6672 = a6670 & a6664;
assign a6674 = l860 & ~i132;
assign a6676 = ~l860 & i132;
assign a6678 = ~a6676 & ~a6674;
assign a6680 = a6678 & a6672;
assign a6682 = l862 & ~i134;
assign a6684 = ~l862 & i134;
assign a6686 = ~a6684 & ~a6682;
assign a6688 = a6686 & a6680;
assign a6690 = l864 & ~i136;
assign a6692 = ~l864 & i136;
assign a6694 = ~a6692 & ~a6690;
assign a6696 = a6694 & a6688;
assign a6698 = l866 & ~i138;
assign a6700 = ~l866 & i138;
assign a6702 = ~a6700 & ~a6698;
assign a6704 = a6702 & a6696;
assign a6706 = l868 & ~i140;
assign a6708 = ~l868 & i140;
assign a6710 = ~a6708 & ~a6706;
assign a6712 = a6710 & a6704;
assign a6714 = l870 & ~i142;
assign a6716 = ~l870 & i142;
assign a6718 = ~a6716 & ~a6714;
assign a6720 = a6718 & a6712;
assign a6722 = l872 & ~i144;
assign a6724 = ~l872 & i144;
assign a6726 = ~a6724 & ~a6722;
assign a6728 = a6726 & a6720;
assign a6730 = l874 & ~i146;
assign a6732 = ~l874 & i146;
assign a6734 = ~a6732 & ~a6730;
assign a6736 = a6734 & a6728;
assign a6738 = l876 & ~i148;
assign a6740 = ~l876 & i148;
assign a6742 = ~a6740 & ~a6738;
assign a6744 = a6742 & a6736;
assign a6746 = l878 & ~i150;
assign a6748 = ~l878 & i150;
assign a6750 = ~a6748 & ~a6746;
assign a6752 = a6750 & a6744;
assign a6754 = l880 & ~i152;
assign a6756 = ~l880 & i152;
assign a6758 = ~a6756 & ~a6754;
assign a6760 = a6758 & a6752;
assign a6762 = l882 & ~i154;
assign a6764 = ~l882 & i154;
assign a6766 = ~a6764 & ~a6762;
assign a6768 = a6766 & a6760;
assign a6770 = l884 & ~i156;
assign a6772 = ~l884 & i156;
assign a6774 = ~a6772 & ~a6770;
assign a6776 = a6774 & a6768;
assign a6778 = l886 & ~i158;
assign a6780 = ~l886 & i158;
assign a6782 = ~a6780 & ~a6778;
assign a6784 = a6782 & a6776;
assign a6786 = l888 & ~i160;
assign a6788 = ~l888 & i160;
assign a6790 = ~a6788 & ~a6786;
assign a6792 = a6790 & a6784;
assign a6794 = l890 & ~i162;
assign a6796 = ~l890 & i162;
assign a6798 = ~a6796 & ~a6794;
assign a6800 = a6798 & a6792;
assign a6802 = l892 & ~i164;
assign a6804 = ~l892 & i164;
assign a6806 = ~a6804 & ~a6802;
assign a6808 = a6806 & a6800;
assign a6810 = l894 & ~i166;
assign a6812 = ~l894 & i166;
assign a6814 = ~a6812 & ~a6810;
assign a6816 = a6814 & a6808;
assign a6818 = l896 & ~i168;
assign a6820 = ~l896 & i168;
assign a6822 = ~a6820 & ~a6818;
assign a6824 = a6822 & a6816;
assign a6826 = l898 & ~i170;
assign a6828 = ~l898 & i170;
assign a6830 = ~a6828 & ~a6826;
assign a6832 = a6830 & a6824;
assign a6834 = l900 & ~i172;
assign a6836 = ~l900 & i172;
assign a6838 = ~a6836 & ~a6834;
assign a6840 = a6838 & a6832;
assign a6842 = l902 & ~i174;
assign a6844 = ~l902 & i174;
assign a6846 = ~a6844 & ~a6842;
assign a6848 = a6846 & a6840;
assign a6850 = l904 & ~i176;
assign a6852 = ~l904 & i176;
assign a6854 = ~a6852 & ~a6850;
assign a6856 = a6854 & a6848;
assign a6858 = l906 & ~i178;
assign a6860 = ~l906 & i178;
assign a6862 = ~a6860 & ~a6858;
assign a6864 = a6862 & a6856;
assign a6866 = l908 & ~i180;
assign a6868 = ~l908 & i180;
assign a6870 = ~a6868 & ~a6866;
assign a6872 = a6870 & a6864;
assign a6874 = l910 & ~i182;
assign a6876 = ~l910 & i182;
assign a6878 = ~a6876 & ~a6874;
assign a6880 = a6878 & a6872;
assign a6882 = l912 & ~i184;
assign a6884 = ~l912 & i184;
assign a6886 = ~a6884 & ~a6882;
assign a6888 = a6886 & a6880;
assign a6890 = l914 & ~i186;
assign a6892 = ~l914 & i186;
assign a6894 = ~a6892 & ~a6890;
assign a6896 = a6894 & a6888;
assign a6898 = l916 & ~i188;
assign a6900 = ~l916 & i188;
assign a6902 = ~a6900 & ~a6898;
assign a6904 = a6902 & a6896;
assign a6906 = l918 & ~i190;
assign a6908 = ~l918 & i190;
assign a6910 = ~a6908 & ~a6906;
assign a6912 = a6910 & a6904;
assign a6914 = l920 & ~i192;
assign a6916 = ~l920 & i192;
assign a6918 = ~a6916 & ~a6914;
assign a6920 = a6918 & a6912;
assign a6922 = l922 & ~i194;
assign a6924 = ~l922 & i194;
assign a6926 = ~a6924 & ~a6922;
assign a6928 = a6926 & a6920;
assign a6930 = l924 & ~i196;
assign a6932 = ~l924 & i196;
assign a6934 = ~a6932 & ~a6930;
assign a6936 = a6934 & a6928;
assign a6938 = l926 & ~i198;
assign a6940 = ~l926 & i198;
assign a6942 = ~a6940 & ~a6938;
assign a6944 = a6942 & a6936;
assign a6946 = l928 & ~i200;
assign a6948 = ~l928 & i200;
assign a6950 = ~a6948 & ~a6946;
assign a6952 = a6950 & a6944;
assign a6954 = l938 & ~i206;
assign a6956 = ~l938 & i206;
assign a6958 = ~a6956 & ~a6954;
assign a6960 = a6958 & a6952;
assign a6962 = a1766 & ~l942;
assign a6964 = a6962 & a1706;
assign a6966 = ~a6964 & a1772;
assign a6968 = ~a6966 & l940;
assign a6970 = a6968 & ~a1762;
assign a6972 = a6970 & ~i208;
assign a6974 = ~a6970 & i208;
assign a6976 = ~a6974 & ~a6972;
assign a6978 = a6976 & a6960;
assign a6980 = l952 & ~i214;
assign a6982 = ~l952 & i214;
assign a6984 = ~a6982 & ~a6980;
assign a6986 = a6984 & a6978;
assign a6988 = a1766 & ~l956;
assign a6990 = a6988 & a1798;
assign a6992 = ~a6990 & a1852;
assign a6994 = ~a6992 & l954;
assign a6996 = a6994 & ~a1846;
assign a6998 = a6996 & ~i216;
assign a7000 = ~a6996 & i216;
assign a7002 = ~a7000 & ~a6998;
assign a7004 = a7002 & a6986;
assign a7006 = l966 & ~i222;
assign a7008 = ~l966 & i222;
assign a7010 = ~a7008 & ~a7006;
assign a7012 = a7010 & a7004;
assign a7014 = a1766 & ~l970;
assign a7016 = a7014 & a1878;
assign a7018 = ~a7016 & a1932;
assign a7020 = ~a7018 & l968;
assign a7022 = a7020 & ~a1926;
assign a7024 = a7022 & ~i224;
assign a7026 = ~a7022 & i224;
assign a7028 = ~a7026 & ~a7024;
assign a7030 = a7028 & a7012;
assign a7032 = l980 & ~i230;
assign a7034 = ~l980 & i230;
assign a7036 = ~a7034 & ~a7032;
assign a7038 = a7036 & a7030;
assign a7040 = a1766 & ~l984;
assign a7042 = a7040 & a1958;
assign a7044 = ~a7042 & a2012;
assign a7046 = ~a7044 & l982;
assign a7048 = a7046 & ~a2006;
assign a7050 = a7048 & ~i232;
assign a7052 = ~a7048 & i232;
assign a7054 = ~a7052 & ~a7050;
assign a7056 = a7054 & a7038;
assign a7058 = a2034 & ~a1946;
assign a7060 = ~a7058 & a1684;
assign a7062 = ~a1684 & ~l992;
assign a7064 = ~a7062 & ~a7060;
assign a7066 = a7064 & ~i234;
assign a7068 = ~a7064 & i234;
assign a7070 = ~a7068 & ~a7066;
assign a7072 = a7070 & a7056;
assign a7074 = ~a1948 & ~l994;
assign a7076 = a7074 & ~a1868;
assign a7078 = ~a7076 & ~a1788;
assign a7080 = a7078 & ~a1690;
assign a7082 = a7080 & ~i236;
assign a7084 = ~a7080 & i236;
assign a7086 = ~a7084 & ~a7082;
assign a7088 = a7086 & a7072;
assign a7090 = ~a1948 & ~l996;
assign a7092 = ~a7090 & ~a1868;
assign a7094 = ~a7092 & ~a1788;
assign a7096 = ~a7094 & ~a1690;
assign a7098 = a7096 & ~i238;
assign a7100 = ~a7096 & i238;
assign a7102 = ~a7100 & ~a7098;
assign a7104 = a7102 & a7088;
assign a7106 = l998 & ~i240;
assign a7108 = ~l998 & i240;
assign a7110 = ~a7108 & ~a7106;
assign a7112 = a7110 & a7104;
assign a7114 = a1766 & l1666;
assign a7116 = ~a1766 & ~l1000;
assign a7118 = ~a7116 & ~a7114;
assign a7120 = a7118 & ~i242;
assign a7122 = ~a7118 & i242;
assign a7124 = ~a7122 & ~a7120;
assign a7126 = a7124 & a7112;
assign a7128 = l1022 & ~i248;
assign a7130 = ~l1022 & i248;
assign a7132 = ~a7130 & ~a7128;
assign a7134 = a7132 & a7126;
assign a7136 = a2652 & ~l1026;
assign a7138 = a7136 & a2592;
assign a7140 = ~a7138 & a2658;
assign a7142 = ~a7140 & l1024;
assign a7144 = a7142 & ~a2648;
assign a7146 = a7144 & ~i250;
assign a7148 = ~a7144 & i250;
assign a7150 = ~a7148 & ~a7146;
assign a7152 = a7150 & a7134;
assign a7154 = l1036 & ~i256;
assign a7156 = ~l1036 & i256;
assign a7158 = ~a7156 & ~a7154;
assign a7160 = a7158 & a7152;
assign a7162 = a2652 & ~l1040;
assign a7164 = a7162 & a2684;
assign a7166 = ~a7164 & a2738;
assign a7168 = ~a7166 & l1038;
assign a7170 = a7168 & ~a2732;
assign a7172 = a7170 & ~i258;
assign a7174 = ~a7170 & i258;
assign a7176 = ~a7174 & ~a7172;
assign a7178 = a7176 & a7160;
assign a7180 = l1050 & ~i264;
assign a7182 = ~l1050 & i264;
assign a7184 = ~a7182 & ~a7180;
assign a7186 = a7184 & a7178;
assign a7188 = a2652 & ~l1054;
assign a7190 = a7188 & a2764;
assign a7192 = ~a7190 & a2818;
assign a7194 = ~a7192 & l1052;
assign a7196 = a7194 & ~a2812;
assign a7198 = a7196 & ~i266;
assign a7200 = ~a7196 & i266;
assign a7202 = ~a7200 & ~a7198;
assign a7204 = a7202 & a7186;
assign a7206 = l1064 & ~i272;
assign a7208 = ~l1064 & i272;
assign a7210 = ~a7208 & ~a7206;
assign a7212 = a7210 & a7204;
assign a7214 = a2652 & ~l1068;
assign a7216 = a7214 & a2844;
assign a7218 = ~a7216 & a2898;
assign a7220 = ~a7218 & l1066;
assign a7222 = a7220 & ~a2892;
assign a7224 = a7222 & ~i274;
assign a7226 = ~a7222 & i274;
assign a7228 = ~a7226 & ~a7224;
assign a7230 = a7228 & a7212;
assign a7232 = a2920 & ~a2832;
assign a7234 = ~a7232 & a2570;
assign a7236 = ~a2570 & ~l1076;
assign a7238 = ~a7236 & ~a7234;
assign a7240 = a7238 & ~i276;
assign a7242 = ~a7238 & i276;
assign a7244 = ~a7242 & ~a7240;
assign a7246 = a7244 & a7230;
assign a7248 = ~a2834 & ~l1078;
assign a7250 = a7248 & ~a2754;
assign a7252 = ~a7250 & ~a2674;
assign a7254 = a7252 & ~a2576;
assign a7256 = a7254 & ~i278;
assign a7258 = ~a7254 & i278;
assign a7260 = ~a7258 & ~a7256;
assign a7262 = a7260 & a7246;
assign a7264 = ~a2834 & ~l1080;
assign a7266 = ~a7264 & ~a2754;
assign a7268 = ~a7266 & ~a2674;
assign a7270 = ~a7268 & ~a2576;
assign a7272 = a7270 & ~i280;
assign a7274 = ~a7270 & i280;
assign a7276 = ~a7274 & ~a7272;
assign a7278 = a7276 & a7262;
assign a7280 = l1082 & ~i282;
assign a7282 = ~l1082 & i282;
assign a7284 = ~a7282 & ~a7280;
assign a7286 = a7284 & a7278;
assign a7288 = a2652 & l1668;
assign a7290 = ~a2652 & ~l1084;
assign a7292 = ~a7290 & ~a7288;
assign a7294 = a7292 & ~i284;
assign a7296 = ~a7292 & i284;
assign a7298 = ~a7296 & ~a7294;
assign a7300 = a7298 & a7286;
assign a7302 = l1106 & ~i290;
assign a7304 = ~l1106 & i290;
assign a7306 = ~a7304 & ~a7302;
assign a7308 = a7306 & a7300;
assign a7310 = a3538 & ~l1110;
assign a7312 = a7310 & a3478;
assign a7314 = ~a7312 & a3544;
assign a7316 = ~a7314 & l1108;
assign a7318 = a7316 & ~a3534;
assign a7320 = a7318 & ~i292;
assign a7322 = ~a7318 & i292;
assign a7324 = ~a7322 & ~a7320;
assign a7326 = a7324 & a7308;
assign a7328 = l1120 & ~i298;
assign a7330 = ~l1120 & i298;
assign a7332 = ~a7330 & ~a7328;
assign a7334 = a7332 & a7326;
assign a7336 = a3538 & ~l1124;
assign a7338 = a7336 & a3570;
assign a7340 = ~a7338 & a3624;
assign a7342 = ~a7340 & l1122;
assign a7344 = a7342 & ~a3618;
assign a7346 = a7344 & ~i300;
assign a7348 = ~a7344 & i300;
assign a7350 = ~a7348 & ~a7346;
assign a7352 = a7350 & a7334;
assign a7354 = l1134 & ~i306;
assign a7356 = ~l1134 & i306;
assign a7358 = ~a7356 & ~a7354;
assign a7360 = a7358 & a7352;
assign a7362 = a3538 & ~l1138;
assign a7364 = a7362 & a3650;
assign a7366 = ~a7364 & a3704;
assign a7368 = ~a7366 & l1136;
assign a7370 = a7368 & ~a3698;
assign a7372 = a7370 & ~i308;
assign a7374 = ~a7370 & i308;
assign a7376 = ~a7374 & ~a7372;
assign a7378 = a7376 & a7360;
assign a7380 = l1148 & ~i314;
assign a7382 = ~l1148 & i314;
assign a7384 = ~a7382 & ~a7380;
assign a7386 = a7384 & a7378;
assign a7388 = a3538 & ~l1152;
assign a7390 = a7388 & a3730;
assign a7392 = ~a7390 & a3784;
assign a7394 = ~a7392 & l1150;
assign a7396 = a7394 & ~a3778;
assign a7398 = a7396 & ~i316;
assign a7400 = ~a7396 & i316;
assign a7402 = ~a7400 & ~a7398;
assign a7404 = a7402 & a7386;
assign a7406 = a3806 & ~a3718;
assign a7408 = ~a7406 & a3456;
assign a7410 = ~a3456 & ~l1160;
assign a7412 = ~a7410 & ~a7408;
assign a7414 = a7412 & ~i318;
assign a7416 = ~a7412 & i318;
assign a7418 = ~a7416 & ~a7414;
assign a7420 = a7418 & a7404;
assign a7422 = ~a3720 & ~l1162;
assign a7424 = a7422 & ~a3640;
assign a7426 = ~a7424 & ~a3560;
assign a7428 = a7426 & ~a3462;
assign a7430 = a7428 & ~i320;
assign a7432 = ~a7428 & i320;
assign a7434 = ~a7432 & ~a7430;
assign a7436 = a7434 & a7420;
assign a7438 = ~a3720 & ~l1164;
assign a7440 = ~a7438 & ~a3640;
assign a7442 = ~a7440 & ~a3560;
assign a7444 = ~a7442 & ~a3462;
assign a7446 = a7444 & ~i322;
assign a7448 = ~a7444 & i322;
assign a7450 = ~a7448 & ~a7446;
assign a7452 = a7450 & a7436;
assign a7454 = l1166 & ~i324;
assign a7456 = ~l1166 & i324;
assign a7458 = ~a7456 & ~a7454;
assign a7460 = a7458 & a7452;
assign a7462 = a3538 & l1670;
assign a7464 = ~a3538 & ~l1168;
assign a7466 = ~a7464 & ~a7462;
assign a7468 = a7466 & ~i326;
assign a7470 = ~a7466 & i326;
assign a7472 = ~a7470 & ~a7468;
assign a7474 = a7472 & a7460;
assign a7476 = l1190 & ~i332;
assign a7478 = ~l1190 & i332;
assign a7480 = ~a7478 & ~a7476;
assign a7482 = a7480 & a7474;
assign a7484 = a4424 & ~l1194;
assign a7486 = a7484 & a4364;
assign a7488 = ~a7486 & a4430;
assign a7490 = ~a7488 & l1192;
assign a7492 = a7490 & ~a4420;
assign a7494 = a7492 & ~i334;
assign a7496 = ~a7492 & i334;
assign a7498 = ~a7496 & ~a7494;
assign a7500 = a7498 & a7482;
assign a7502 = l1204 & ~i340;
assign a7504 = ~l1204 & i340;
assign a7506 = ~a7504 & ~a7502;
assign a7508 = a7506 & a7500;
assign a7510 = a4424 & ~l1208;
assign a7512 = a7510 & a4456;
assign a7514 = ~a7512 & a4510;
assign a7516 = ~a7514 & l1206;
assign a7518 = a7516 & ~a4504;
assign a7520 = a7518 & ~i342;
assign a7522 = ~a7518 & i342;
assign a7524 = ~a7522 & ~a7520;
assign a7526 = a7524 & a7508;
assign a7528 = l1218 & ~i348;
assign a7530 = ~l1218 & i348;
assign a7532 = ~a7530 & ~a7528;
assign a7534 = a7532 & a7526;
assign a7536 = a4424 & ~l1222;
assign a7538 = a7536 & a4536;
assign a7540 = ~a7538 & a4590;
assign a7542 = ~a7540 & l1220;
assign a7544 = a7542 & ~a4584;
assign a7546 = a7544 & ~i350;
assign a7548 = ~a7544 & i350;
assign a7550 = ~a7548 & ~a7546;
assign a7552 = a7550 & a7534;
assign a7554 = l1232 & ~i356;
assign a7556 = ~l1232 & i356;
assign a7558 = ~a7556 & ~a7554;
assign a7560 = a7558 & a7552;
assign a7562 = a4424 & ~l1236;
assign a7564 = a7562 & a4616;
assign a7566 = ~a7564 & a4670;
assign a7568 = ~a7566 & l1234;
assign a7570 = a7568 & ~a4664;
assign a7572 = a7570 & ~i358;
assign a7574 = ~a7570 & i358;
assign a7576 = ~a7574 & ~a7572;
assign a7578 = a7576 & a7560;
assign a7580 = a4692 & ~a4604;
assign a7582 = ~a7580 & a4342;
assign a7584 = ~a4342 & ~l1244;
assign a7586 = ~a7584 & ~a7582;
assign a7588 = a7586 & ~i360;
assign a7590 = ~a7586 & i360;
assign a7592 = ~a7590 & ~a7588;
assign a7594 = a7592 & a7578;
assign a7596 = ~a4606 & ~l1246;
assign a7598 = a7596 & ~a4526;
assign a7600 = ~a7598 & ~a4446;
assign a7602 = a7600 & ~a4348;
assign a7604 = a7602 & ~i362;
assign a7606 = ~a7602 & i362;
assign a7608 = ~a7606 & ~a7604;
assign a7610 = a7608 & a7594;
assign a7612 = ~a4606 & ~l1248;
assign a7614 = ~a7612 & ~a4526;
assign a7616 = ~a7614 & ~a4446;
assign a7618 = ~a7616 & ~a4348;
assign a7620 = a7618 & ~i364;
assign a7622 = ~a7618 & i364;
assign a7624 = ~a7622 & ~a7620;
assign a7626 = a7624 & a7610;
assign a7628 = l1250 & ~i366;
assign a7630 = ~l1250 & i366;
assign a7632 = ~a7630 & ~a7628;
assign a7634 = a7632 & a7626;
assign a7636 = a4424 & l1672;
assign a7638 = ~a4424 & ~l1252;
assign a7640 = ~a7638 & ~a7636;
assign a7642 = a7640 & ~i368;
assign a7644 = ~a7640 & i368;
assign a7646 = ~a7644 & ~a7642;
assign a7648 = a7646 & a7634;
assign a7650 = l1274 & ~i374;
assign a7652 = ~l1274 & i374;
assign a7654 = ~a7652 & ~a7650;
assign a7656 = a7654 & a7648;
assign a7658 = a5310 & ~l1278;
assign a7660 = a7658 & a5250;
assign a7662 = ~a7660 & a5316;
assign a7664 = ~a7662 & l1276;
assign a7666 = a7664 & ~a5306;
assign a7668 = a7666 & ~i376;
assign a7670 = ~a7666 & i376;
assign a7672 = ~a7670 & ~a7668;
assign a7674 = a7672 & a7656;
assign a7676 = l1288 & ~i382;
assign a7678 = ~l1288 & i382;
assign a7680 = ~a7678 & ~a7676;
assign a7682 = a7680 & a7674;
assign a7684 = a5310 & ~l1292;
assign a7686 = a7684 & a5342;
assign a7688 = ~a7686 & a5396;
assign a7690 = ~a7688 & l1290;
assign a7692 = a7690 & ~a5390;
assign a7694 = a7692 & ~i384;
assign a7696 = ~a7692 & i384;
assign a7698 = ~a7696 & ~a7694;
assign a7700 = a7698 & a7682;
assign a7702 = l1302 & ~i390;
assign a7704 = ~l1302 & i390;
assign a7706 = ~a7704 & ~a7702;
assign a7708 = a7706 & a7700;
assign a7710 = a5310 & ~l1306;
assign a7712 = a7710 & a5422;
assign a7714 = ~a7712 & a5476;
assign a7716 = ~a7714 & l1304;
assign a7718 = a7716 & ~a5470;
assign a7720 = a7718 & ~i392;
assign a7722 = ~a7718 & i392;
assign a7724 = ~a7722 & ~a7720;
assign a7726 = a7724 & a7708;
assign a7728 = l1316 & ~i398;
assign a7730 = ~l1316 & i398;
assign a7732 = ~a7730 & ~a7728;
assign a7734 = a7732 & a7726;
assign a7736 = a5310 & ~l1320;
assign a7738 = a7736 & a5502;
assign a7740 = ~a7738 & a5556;
assign a7742 = ~a7740 & l1318;
assign a7744 = a7742 & ~a5550;
assign a7746 = a7744 & ~i400;
assign a7748 = ~a7744 & i400;
assign a7750 = ~a7748 & ~a7746;
assign a7752 = a7750 & a7734;
assign a7754 = a5578 & ~a5490;
assign a7756 = ~a7754 & a5228;
assign a7758 = ~a5228 & ~l1328;
assign a7760 = ~a7758 & ~a7756;
assign a7762 = a7760 & ~i402;
assign a7764 = ~a7760 & i402;
assign a7766 = ~a7764 & ~a7762;
assign a7768 = a7766 & a7752;
assign a7770 = ~a5492 & ~l1330;
assign a7772 = a7770 & ~a5412;
assign a7774 = ~a7772 & ~a5332;
assign a7776 = a7774 & ~a5234;
assign a7778 = a7776 & ~i404;
assign a7780 = ~a7776 & i404;
assign a7782 = ~a7780 & ~a7778;
assign a7784 = a7782 & a7768;
assign a7786 = ~a5492 & ~l1332;
assign a7788 = ~a7786 & ~a5412;
assign a7790 = ~a7788 & ~a5332;
assign a7792 = ~a7790 & ~a5234;
assign a7794 = a7792 & ~i406;
assign a7796 = ~a7792 & i406;
assign a7798 = ~a7796 & ~a7794;
assign a7800 = a7798 & a7784;
assign a7802 = l1334 & ~i408;
assign a7804 = ~l1334 & i408;
assign a7806 = ~a7804 & ~a7802;
assign a7808 = a7806 & a7800;
assign a7810 = a5310 & l1674;
assign a7812 = ~a5310 & ~l1336;
assign a7814 = ~a7812 & ~a7810;
assign a7816 = a7814 & ~i410;
assign a7818 = ~a7814 & i410;
assign a7820 = ~a7818 & ~a7816;
assign a7822 = a7820 & a7808;
assign a7824 = ~l1664 & l1662;
assign a7826 = a7824 & ~l934;
assign a7828 = ~a7824 & ~l1358;
assign a7830 = ~a7828 & ~a7826;
assign a7832 = a7830 & ~i418;
assign a7834 = ~a7830 & i418;
assign a7836 = ~a7834 & ~a7832;
assign a7838 = a7836 & a7822;
assign a7840 = ~a7824 & ~l1360;
assign a7842 = a7824 & l936;
assign a7844 = ~a7842 & ~a7840;
assign a7846 = a7844 & ~i420;
assign a7848 = ~a7844 & i420;
assign a7850 = ~a7848 & ~a7846;
assign a7852 = a7850 & a7838;
assign a7854 = a7824 & ~l940;
assign a7856 = ~a7824 & ~l1362;
assign a7858 = ~a7856 & ~a7854;
assign a7860 = a7858 & ~i422;
assign a7862 = ~a7858 & i422;
assign a7864 = ~a7862 & ~a7860;
assign a7866 = a7864 & a7852;
assign a7868 = ~a7824 & ~l1364;
assign a7870 = a7824 & l942;
assign a7872 = ~a7870 & ~a7868;
assign a7874 = a7872 & ~i424;
assign a7876 = ~a7872 & i424;
assign a7878 = ~a7876 & ~a7874;
assign a7880 = a7878 & a7866;
assign a7882 = a7824 & ~l948;
assign a7884 = ~a7824 & ~l1366;
assign a7886 = ~a7884 & ~a7882;
assign a7888 = a7886 & ~i426;
assign a7890 = ~a7886 & i426;
assign a7892 = ~a7890 & ~a7888;
assign a7894 = a7892 & a7880;
assign a7896 = ~a7824 & ~l1368;
assign a7898 = a7824 & l950;
assign a7900 = ~a7898 & ~a7896;
assign a7902 = a7900 & ~i428;
assign a7904 = ~a7900 & i428;
assign a7906 = ~a7904 & ~a7902;
assign a7908 = a7906 & a7894;
assign a7910 = a7824 & ~l954;
assign a7912 = ~a7824 & ~l1370;
assign a7914 = ~a7912 & ~a7910;
assign a7916 = a7914 & ~i430;
assign a7918 = ~a7914 & i430;
assign a7920 = ~a7918 & ~a7916;
assign a7922 = a7920 & a7908;
assign a7924 = ~a7824 & ~l1372;
assign a7926 = a7824 & l956;
assign a7928 = ~a7926 & ~a7924;
assign a7930 = a7928 & ~i432;
assign a7932 = ~a7928 & i432;
assign a7934 = ~a7932 & ~a7930;
assign a7936 = a7934 & a7922;
assign a7938 = a7824 & ~l962;
assign a7940 = ~a7824 & ~l1374;
assign a7942 = ~a7940 & ~a7938;
assign a7944 = a7942 & ~i434;
assign a7946 = ~a7942 & i434;
assign a7948 = ~a7946 & ~a7944;
assign a7950 = a7948 & a7936;
assign a7952 = ~a7824 & ~l1376;
assign a7954 = a7824 & l964;
assign a7956 = ~a7954 & ~a7952;
assign a7958 = a7956 & ~i436;
assign a7960 = ~a7956 & i436;
assign a7962 = ~a7960 & ~a7958;
assign a7964 = a7962 & a7950;
assign a7966 = a7824 & ~l968;
assign a7968 = ~a7824 & ~l1378;
assign a7970 = ~a7968 & ~a7966;
assign a7972 = a7970 & ~i438;
assign a7974 = ~a7970 & i438;
assign a7976 = ~a7974 & ~a7972;
assign a7978 = a7976 & a7964;
assign a7980 = ~a7824 & ~l1380;
assign a7982 = a7824 & l970;
assign a7984 = ~a7982 & ~a7980;
assign a7986 = a7984 & ~i440;
assign a7988 = ~a7984 & i440;
assign a7990 = ~a7988 & ~a7986;
assign a7992 = a7990 & a7978;
assign a7994 = a7824 & ~l976;
assign a7996 = ~a7824 & ~l1382;
assign a7998 = ~a7996 & ~a7994;
assign a8000 = a7998 & ~i442;
assign a8002 = ~a7998 & i442;
assign a8004 = ~a8002 & ~a8000;
assign a8006 = a8004 & a7992;
assign a8008 = ~a7824 & ~l1384;
assign a8010 = a7824 & l978;
assign a8012 = ~a8010 & ~a8008;
assign a8014 = a8012 & ~i444;
assign a8016 = ~a8012 & i444;
assign a8018 = ~a8016 & ~a8014;
assign a8020 = a8018 & a8006;
assign a8022 = a7824 & ~l982;
assign a8024 = ~a7824 & ~l1386;
assign a8026 = ~a8024 & ~a8022;
assign a8028 = a8026 & ~i446;
assign a8030 = ~a8026 & i446;
assign a8032 = ~a8030 & ~a8028;
assign a8034 = a8032 & a8020;
assign a8036 = ~a7824 & ~l1388;
assign a8038 = a7824 & l984;
assign a8040 = ~a8038 & ~a8036;
assign a8042 = a8040 & ~i448;
assign a8044 = ~a8040 & i448;
assign a8046 = ~a8044 & ~a8042;
assign a8048 = a8046 & a8034;
assign a8050 = a7824 & ~l986;
assign a8052 = ~a7824 & ~l1390;
assign a8054 = ~a8052 & ~a8050;
assign a8056 = a8054 & ~i450;
assign a8058 = ~a8054 & i450;
assign a8060 = ~a8058 & ~a8056;
assign a8062 = a8060 & a8048;
assign a8064 = a7824 & ~l988;
assign a8066 = ~a7824 & ~l1392;
assign a8068 = ~a8066 & ~a8064;
assign a8070 = a8068 & ~i452;
assign a8072 = ~a8068 & i452;
assign a8074 = ~a8072 & ~a8070;
assign a8076 = a8074 & a8062;
assign a8078 = ~a7824 & ~l1394;
assign a8080 = a7824 & l990;
assign a8082 = ~a8080 & ~a8078;
assign a8084 = a8082 & ~i454;
assign a8086 = ~a8082 & i454;
assign a8088 = ~a8086 & ~a8084;
assign a8090 = a8088 & a8076;
assign a8092 = a7824 & ~l992;
assign a8094 = ~a7824 & ~l1396;
assign a8096 = ~a8094 & ~a8092;
assign a8098 = a8096 & ~i456;
assign a8100 = ~a8096 & i456;
assign a8102 = ~a8100 & ~a8098;
assign a8104 = a8102 & a8090;
assign a8106 = a7824 & ~l994;
assign a8108 = ~a7824 & ~l1398;
assign a8110 = ~a8108 & ~a8106;
assign a8112 = a8110 & ~i458;
assign a8114 = ~a8110 & i458;
assign a8116 = ~a8114 & ~a8112;
assign a8118 = a8116 & a8104;
assign a8120 = a7824 & ~l996;
assign a8122 = ~a7824 & ~l1400;
assign a8124 = ~a8122 & ~a8120;
assign a8126 = a8124 & ~i460;
assign a8128 = ~a8124 & i460;
assign a8130 = ~a8128 & ~a8126;
assign a8132 = a8130 & a8118;
assign a8134 = a7824 & ~l1000;
assign a8136 = ~a7824 & ~l1402;
assign a8138 = ~a8136 & ~a8134;
assign a8140 = a8138 & ~i462;
assign a8142 = ~a8138 & i462;
assign a8144 = ~a8142 & ~a8140;
assign a8146 = a8144 & a8132;
assign a8148 = a7824 & ~l1002;
assign a8150 = ~a7824 & ~l1404;
assign a8152 = ~a8150 & ~a8148;
assign a8154 = a8152 & ~i464;
assign a8156 = ~a8152 & i464;
assign a8158 = ~a8156 & ~a8154;
assign a8160 = a8158 & a8146;
assign a8162 = a7824 & ~l1004;
assign a8164 = ~a7824 & ~l1406;
assign a8166 = ~a8164 & ~a8162;
assign a8168 = a8166 & ~i466;
assign a8170 = ~a8166 & i466;
assign a8172 = ~a8170 & ~a8168;
assign a8174 = a8172 & a8160;
assign a8176 = a7824 & ~l1006;
assign a8178 = ~a7824 & ~l1408;
assign a8180 = ~a8178 & ~a8176;
assign a8182 = a8180 & ~i468;
assign a8184 = ~a8180 & i468;
assign a8186 = ~a8184 & ~a8182;
assign a8188 = a8186 & a8174;
assign a8190 = a7824 & ~l1008;
assign a8192 = ~a7824 & ~l1410;
assign a8194 = ~a8192 & ~a8190;
assign a8196 = a8194 & ~i470;
assign a8198 = ~a8194 & i470;
assign a8200 = ~a8198 & ~a8196;
assign a8202 = a8200 & a8188;
assign a8204 = a7824 & ~l1010;
assign a8206 = ~a7824 & ~l1412;
assign a8208 = ~a8206 & ~a8204;
assign a8210 = a8208 & ~i472;
assign a8212 = ~a8208 & i472;
assign a8214 = ~a8212 & ~a8210;
assign a8216 = a8214 & a8202;
assign a8218 = a7824 & ~l1012;
assign a8220 = ~a7824 & ~l1414;
assign a8222 = ~a8220 & ~a8218;
assign a8224 = a8222 & ~i474;
assign a8226 = ~a8222 & i474;
assign a8228 = ~a8226 & ~a8224;
assign a8230 = a8228 & a8216;
assign a8232 = a7824 & ~l1018;
assign a8234 = ~a7824 & ~l1416;
assign a8236 = ~a8234 & ~a8232;
assign a8238 = a8236 & ~i476;
assign a8240 = ~a8236 & i476;
assign a8242 = ~a8240 & ~a8238;
assign a8244 = a8242 & a8230;
assign a8246 = ~a7824 & ~l1418;
assign a8248 = a7824 & l1020;
assign a8250 = ~a8248 & ~a8246;
assign a8252 = a8250 & ~i478;
assign a8254 = ~a8250 & i478;
assign a8256 = ~a8254 & ~a8252;
assign a8258 = a8256 & a8244;
assign a8260 = a7824 & ~l1024;
assign a8262 = ~a7824 & ~l1420;
assign a8264 = ~a8262 & ~a8260;
assign a8266 = a8264 & ~i480;
assign a8268 = ~a8264 & i480;
assign a8270 = ~a8268 & ~a8266;
assign a8272 = a8270 & a8258;
assign a8274 = ~a7824 & ~l1422;
assign a8276 = a7824 & l1026;
assign a8278 = ~a8276 & ~a8274;
assign a8280 = a8278 & ~i482;
assign a8282 = ~a8278 & i482;
assign a8284 = ~a8282 & ~a8280;
assign a8286 = a8284 & a8272;
assign a8288 = a7824 & ~l1032;
assign a8290 = ~a7824 & ~l1424;
assign a8292 = ~a8290 & ~a8288;
assign a8294 = a8292 & ~i484;
assign a8296 = ~a8292 & i484;
assign a8298 = ~a8296 & ~a8294;
assign a8300 = a8298 & a8286;
assign a8302 = ~a7824 & ~l1426;
assign a8304 = a7824 & l1034;
assign a8306 = ~a8304 & ~a8302;
assign a8308 = a8306 & ~i486;
assign a8310 = ~a8306 & i486;
assign a8312 = ~a8310 & ~a8308;
assign a8314 = a8312 & a8300;
assign a8316 = a7824 & ~l1038;
assign a8318 = ~a7824 & ~l1428;
assign a8320 = ~a8318 & ~a8316;
assign a8322 = a8320 & ~i488;
assign a8324 = ~a8320 & i488;
assign a8326 = ~a8324 & ~a8322;
assign a8328 = a8326 & a8314;
assign a8330 = ~a7824 & ~l1430;
assign a8332 = a7824 & l1040;
assign a8334 = ~a8332 & ~a8330;
assign a8336 = a8334 & ~i490;
assign a8338 = ~a8334 & i490;
assign a8340 = ~a8338 & ~a8336;
assign a8342 = a8340 & a8328;
assign a8344 = a7824 & ~l1046;
assign a8346 = ~a7824 & ~l1432;
assign a8348 = ~a8346 & ~a8344;
assign a8350 = a8348 & ~i492;
assign a8352 = ~a8348 & i492;
assign a8354 = ~a8352 & ~a8350;
assign a8356 = a8354 & a8342;
assign a8358 = ~a7824 & ~l1434;
assign a8360 = a7824 & l1048;
assign a8362 = ~a8360 & ~a8358;
assign a8364 = a8362 & ~i494;
assign a8366 = ~a8362 & i494;
assign a8368 = ~a8366 & ~a8364;
assign a8370 = a8368 & a8356;
assign a8372 = a7824 & ~l1052;
assign a8374 = ~a7824 & ~l1436;
assign a8376 = ~a8374 & ~a8372;
assign a8378 = a8376 & ~i496;
assign a8380 = ~a8376 & i496;
assign a8382 = ~a8380 & ~a8378;
assign a8384 = a8382 & a8370;
assign a8386 = ~a7824 & ~l1438;
assign a8388 = a7824 & l1054;
assign a8390 = ~a8388 & ~a8386;
assign a8392 = a8390 & ~i498;
assign a8394 = ~a8390 & i498;
assign a8396 = ~a8394 & ~a8392;
assign a8398 = a8396 & a8384;
assign a8400 = a7824 & ~l1060;
assign a8402 = ~a7824 & ~l1440;
assign a8404 = ~a8402 & ~a8400;
assign a8406 = a8404 & ~i500;
assign a8408 = ~a8404 & i500;
assign a8410 = ~a8408 & ~a8406;
assign a8412 = a8410 & a8398;
assign a8414 = ~a7824 & ~l1442;
assign a8416 = a7824 & l1062;
assign a8418 = ~a8416 & ~a8414;
assign a8420 = a8418 & ~i502;
assign a8422 = ~a8418 & i502;
assign a8424 = ~a8422 & ~a8420;
assign a8426 = a8424 & a8412;
assign a8428 = a7824 & ~l1066;
assign a8430 = ~a7824 & ~l1444;
assign a8432 = ~a8430 & ~a8428;
assign a8434 = a8432 & ~i504;
assign a8436 = ~a8432 & i504;
assign a8438 = ~a8436 & ~a8434;
assign a8440 = a8438 & a8426;
assign a8442 = ~a7824 & ~l1446;
assign a8444 = a7824 & l1068;
assign a8446 = ~a8444 & ~a8442;
assign a8448 = a8446 & ~i506;
assign a8450 = ~a8446 & i506;
assign a8452 = ~a8450 & ~a8448;
assign a8454 = a8452 & a8440;
assign a8456 = a7824 & ~l1070;
assign a8458 = ~a7824 & ~l1448;
assign a8460 = ~a8458 & ~a8456;
assign a8462 = a8460 & ~i508;
assign a8464 = ~a8460 & i508;
assign a8466 = ~a8464 & ~a8462;
assign a8468 = a8466 & a8454;
assign a8470 = a7824 & ~l1072;
assign a8472 = ~a7824 & ~l1450;
assign a8474 = ~a8472 & ~a8470;
assign a8476 = a8474 & ~i510;
assign a8478 = ~a8474 & i510;
assign a8480 = ~a8478 & ~a8476;
assign a8482 = a8480 & a8468;
assign a8484 = ~a7824 & ~l1452;
assign a8486 = a7824 & l1074;
assign a8488 = ~a8486 & ~a8484;
assign a8490 = a8488 & ~i512;
assign a8492 = ~a8488 & i512;
assign a8494 = ~a8492 & ~a8490;
assign a8496 = a8494 & a8482;
assign a8498 = a7824 & ~l1076;
assign a8500 = ~a7824 & ~l1454;
assign a8502 = ~a8500 & ~a8498;
assign a8504 = a8502 & ~i514;
assign a8506 = ~a8502 & i514;
assign a8508 = ~a8506 & ~a8504;
assign a8510 = a8508 & a8496;
assign a8512 = a7824 & ~l1078;
assign a8514 = ~a7824 & ~l1456;
assign a8516 = ~a8514 & ~a8512;
assign a8518 = a8516 & ~i516;
assign a8520 = ~a8516 & i516;
assign a8522 = ~a8520 & ~a8518;
assign a8524 = a8522 & a8510;
assign a8526 = a7824 & ~l1080;
assign a8528 = ~a7824 & ~l1458;
assign a8530 = ~a8528 & ~a8526;
assign a8532 = a8530 & ~i518;
assign a8534 = ~a8530 & i518;
assign a8536 = ~a8534 & ~a8532;
assign a8538 = a8536 & a8524;
assign a8540 = a7824 & ~l1084;
assign a8542 = ~a7824 & ~l1460;
assign a8544 = ~a8542 & ~a8540;
assign a8546 = a8544 & ~i520;
assign a8548 = ~a8544 & i520;
assign a8550 = ~a8548 & ~a8546;
assign a8552 = a8550 & a8538;
assign a8554 = a7824 & ~l1086;
assign a8556 = ~a7824 & ~l1462;
assign a8558 = ~a8556 & ~a8554;
assign a8560 = a8558 & ~i522;
assign a8562 = ~a8558 & i522;
assign a8564 = ~a8562 & ~a8560;
assign a8566 = a8564 & a8552;
assign a8568 = a7824 & ~l1088;
assign a8570 = ~a7824 & ~l1464;
assign a8572 = ~a8570 & ~a8568;
assign a8574 = a8572 & ~i524;
assign a8576 = ~a8572 & i524;
assign a8578 = ~a8576 & ~a8574;
assign a8580 = a8578 & a8566;
assign a8582 = a7824 & ~l1090;
assign a8584 = ~a7824 & ~l1466;
assign a8586 = ~a8584 & ~a8582;
assign a8588 = a8586 & ~i526;
assign a8590 = ~a8586 & i526;
assign a8592 = ~a8590 & ~a8588;
assign a8594 = a8592 & a8580;
assign a8596 = a7824 & ~l1092;
assign a8598 = ~a7824 & ~l1468;
assign a8600 = ~a8598 & ~a8596;
assign a8602 = a8600 & ~i528;
assign a8604 = ~a8600 & i528;
assign a8606 = ~a8604 & ~a8602;
assign a8608 = a8606 & a8594;
assign a8610 = a7824 & ~l1094;
assign a8612 = ~a7824 & ~l1470;
assign a8614 = ~a8612 & ~a8610;
assign a8616 = a8614 & ~i530;
assign a8618 = ~a8614 & i530;
assign a8620 = ~a8618 & ~a8616;
assign a8622 = a8620 & a8608;
assign a8624 = a7824 & ~l1096;
assign a8626 = ~a7824 & ~l1472;
assign a8628 = ~a8626 & ~a8624;
assign a8630 = a8628 & ~i532;
assign a8632 = ~a8628 & i532;
assign a8634 = ~a8632 & ~a8630;
assign a8636 = a8634 & a8622;
assign a8638 = a7824 & ~l1102;
assign a8640 = ~a7824 & ~l1474;
assign a8642 = ~a8640 & ~a8638;
assign a8644 = a8642 & ~i534;
assign a8646 = ~a8642 & i534;
assign a8648 = ~a8646 & ~a8644;
assign a8650 = a8648 & a8636;
assign a8652 = ~a7824 & ~l1476;
assign a8654 = a7824 & l1104;
assign a8656 = ~a8654 & ~a8652;
assign a8658 = a8656 & ~i536;
assign a8660 = ~a8656 & i536;
assign a8662 = ~a8660 & ~a8658;
assign a8664 = a8662 & a8650;
assign a8666 = a7824 & ~l1108;
assign a8668 = ~a7824 & ~l1478;
assign a8670 = ~a8668 & ~a8666;
assign a8672 = a8670 & ~i538;
assign a8674 = ~a8670 & i538;
assign a8676 = ~a8674 & ~a8672;
assign a8678 = a8676 & a8664;
assign a8680 = ~a7824 & ~l1480;
assign a8682 = a7824 & l1110;
assign a8684 = ~a8682 & ~a8680;
assign a8686 = a8684 & ~i540;
assign a8688 = ~a8684 & i540;
assign a8690 = ~a8688 & ~a8686;
assign a8692 = a8690 & a8678;
assign a8694 = a7824 & ~l1116;
assign a8696 = ~a7824 & ~l1482;
assign a8698 = ~a8696 & ~a8694;
assign a8700 = a8698 & ~i542;
assign a8702 = ~a8698 & i542;
assign a8704 = ~a8702 & ~a8700;
assign a8706 = a8704 & a8692;
assign a8708 = ~a7824 & ~l1484;
assign a8710 = a7824 & l1118;
assign a8712 = ~a8710 & ~a8708;
assign a8714 = a8712 & ~i544;
assign a8716 = ~a8712 & i544;
assign a8718 = ~a8716 & ~a8714;
assign a8720 = a8718 & a8706;
assign a8722 = a7824 & ~l1122;
assign a8724 = ~a7824 & ~l1486;
assign a8726 = ~a8724 & ~a8722;
assign a8728 = a8726 & ~i546;
assign a8730 = ~a8726 & i546;
assign a8732 = ~a8730 & ~a8728;
assign a8734 = a8732 & a8720;
assign a8736 = ~a7824 & ~l1488;
assign a8738 = a7824 & l1124;
assign a8740 = ~a8738 & ~a8736;
assign a8742 = a8740 & ~i548;
assign a8744 = ~a8740 & i548;
assign a8746 = ~a8744 & ~a8742;
assign a8748 = a8746 & a8734;
assign a8750 = a7824 & ~l1130;
assign a8752 = ~a7824 & ~l1490;
assign a8754 = ~a8752 & ~a8750;
assign a8756 = a8754 & ~i550;
assign a8758 = ~a8754 & i550;
assign a8760 = ~a8758 & ~a8756;
assign a8762 = a8760 & a8748;
assign a8764 = ~a7824 & ~l1492;
assign a8766 = a7824 & l1132;
assign a8768 = ~a8766 & ~a8764;
assign a8770 = a8768 & ~i552;
assign a8772 = ~a8768 & i552;
assign a8774 = ~a8772 & ~a8770;
assign a8776 = a8774 & a8762;
assign a8778 = a7824 & ~l1136;
assign a8780 = ~a7824 & ~l1494;
assign a8782 = ~a8780 & ~a8778;
assign a8784 = a8782 & ~i554;
assign a8786 = ~a8782 & i554;
assign a8788 = ~a8786 & ~a8784;
assign a8790 = a8788 & a8776;
assign a8792 = ~a7824 & ~l1496;
assign a8794 = a7824 & l1138;
assign a8796 = ~a8794 & ~a8792;
assign a8798 = a8796 & ~i556;
assign a8800 = ~a8796 & i556;
assign a8802 = ~a8800 & ~a8798;
assign a8804 = a8802 & a8790;
assign a8806 = a7824 & ~l1144;
assign a8808 = ~a7824 & ~l1498;
assign a8810 = ~a8808 & ~a8806;
assign a8812 = a8810 & ~i558;
assign a8814 = ~a8810 & i558;
assign a8816 = ~a8814 & ~a8812;
assign a8818 = a8816 & a8804;
assign a8820 = ~a7824 & ~l1500;
assign a8822 = a7824 & l1146;
assign a8824 = ~a8822 & ~a8820;
assign a8826 = a8824 & ~i560;
assign a8828 = ~a8824 & i560;
assign a8830 = ~a8828 & ~a8826;
assign a8832 = a8830 & a8818;
assign a8834 = a7824 & ~l1150;
assign a8836 = ~a7824 & ~l1502;
assign a8838 = ~a8836 & ~a8834;
assign a8840 = a8838 & ~i562;
assign a8842 = ~a8838 & i562;
assign a8844 = ~a8842 & ~a8840;
assign a8846 = a8844 & a8832;
assign a8848 = ~a7824 & ~l1504;
assign a8850 = a7824 & l1152;
assign a8852 = ~a8850 & ~a8848;
assign a8854 = a8852 & ~i564;
assign a8856 = ~a8852 & i564;
assign a8858 = ~a8856 & ~a8854;
assign a8860 = a8858 & a8846;
assign a8862 = a7824 & ~l1154;
assign a8864 = ~a7824 & ~l1506;
assign a8866 = ~a8864 & ~a8862;
assign a8868 = a8866 & ~i566;
assign a8870 = ~a8866 & i566;
assign a8872 = ~a8870 & ~a8868;
assign a8874 = a8872 & a8860;
assign a8876 = a7824 & ~l1156;
assign a8878 = ~a7824 & ~l1508;
assign a8880 = ~a8878 & ~a8876;
assign a8882 = a8880 & ~i568;
assign a8884 = ~a8880 & i568;
assign a8886 = ~a8884 & ~a8882;
assign a8888 = a8886 & a8874;
assign a8890 = ~a7824 & ~l1510;
assign a8892 = a7824 & l1158;
assign a8894 = ~a8892 & ~a8890;
assign a8896 = a8894 & ~i570;
assign a8898 = ~a8894 & i570;
assign a8900 = ~a8898 & ~a8896;
assign a8902 = a8900 & a8888;
assign a8904 = a7824 & ~l1160;
assign a8906 = ~a7824 & ~l1512;
assign a8908 = ~a8906 & ~a8904;
assign a8910 = a8908 & ~i572;
assign a8912 = ~a8908 & i572;
assign a8914 = ~a8912 & ~a8910;
assign a8916 = a8914 & a8902;
assign a8918 = a7824 & ~l1162;
assign a8920 = ~a7824 & ~l1514;
assign a8922 = ~a8920 & ~a8918;
assign a8924 = a8922 & ~i574;
assign a8926 = ~a8922 & i574;
assign a8928 = ~a8926 & ~a8924;
assign a8930 = a8928 & a8916;
assign a8932 = a7824 & ~l1164;
assign a8934 = ~a7824 & ~l1516;
assign a8936 = ~a8934 & ~a8932;
assign a8938 = a8936 & ~i576;
assign a8940 = ~a8936 & i576;
assign a8942 = ~a8940 & ~a8938;
assign a8944 = a8942 & a8930;
assign a8946 = a7824 & ~l1168;
assign a8948 = ~a7824 & ~l1518;
assign a8950 = ~a8948 & ~a8946;
assign a8952 = a8950 & ~i578;
assign a8954 = ~a8950 & i578;
assign a8956 = ~a8954 & ~a8952;
assign a8958 = a8956 & a8944;
assign a8960 = a7824 & ~l1170;
assign a8962 = ~a7824 & ~l1520;
assign a8964 = ~a8962 & ~a8960;
assign a8966 = a8964 & ~i580;
assign a8968 = ~a8964 & i580;
assign a8970 = ~a8968 & ~a8966;
assign a8972 = a8970 & a8958;
assign a8974 = a7824 & ~l1172;
assign a8976 = ~a7824 & ~l1522;
assign a8978 = ~a8976 & ~a8974;
assign a8980 = a8978 & ~i582;
assign a8982 = ~a8978 & i582;
assign a8984 = ~a8982 & ~a8980;
assign a8986 = a8984 & a8972;
assign a8988 = a7824 & ~l1174;
assign a8990 = ~a7824 & ~l1524;
assign a8992 = ~a8990 & ~a8988;
assign a8994 = a8992 & ~i584;
assign a8996 = ~a8992 & i584;
assign a8998 = ~a8996 & ~a8994;
assign a9000 = a8998 & a8986;
assign a9002 = a7824 & ~l1176;
assign a9004 = ~a7824 & ~l1526;
assign a9006 = ~a9004 & ~a9002;
assign a9008 = a9006 & ~i586;
assign a9010 = ~a9006 & i586;
assign a9012 = ~a9010 & ~a9008;
assign a9014 = a9012 & a9000;
assign a9016 = a7824 & ~l1178;
assign a9018 = ~a7824 & ~l1528;
assign a9020 = ~a9018 & ~a9016;
assign a9022 = a9020 & ~i588;
assign a9024 = ~a9020 & i588;
assign a9026 = ~a9024 & ~a9022;
assign a9028 = a9026 & a9014;
assign a9030 = a7824 & ~l1180;
assign a9032 = ~a7824 & ~l1530;
assign a9034 = ~a9032 & ~a9030;
assign a9036 = a9034 & ~i590;
assign a9038 = ~a9034 & i590;
assign a9040 = ~a9038 & ~a9036;
assign a9042 = a9040 & a9028;
assign a9044 = a7824 & ~l1186;
assign a9046 = ~a7824 & ~l1532;
assign a9048 = ~a9046 & ~a9044;
assign a9050 = a9048 & ~i592;
assign a9052 = ~a9048 & i592;
assign a9054 = ~a9052 & ~a9050;
assign a9056 = a9054 & a9042;
assign a9058 = ~a7824 & ~l1534;
assign a9060 = a7824 & l1188;
assign a9062 = ~a9060 & ~a9058;
assign a9064 = a9062 & ~i594;
assign a9066 = ~a9062 & i594;
assign a9068 = ~a9066 & ~a9064;
assign a9070 = a9068 & a9056;
assign a9072 = a7824 & ~l1192;
assign a9074 = ~a7824 & ~l1536;
assign a9076 = ~a9074 & ~a9072;
assign a9078 = a9076 & ~i596;
assign a9080 = ~a9076 & i596;
assign a9082 = ~a9080 & ~a9078;
assign a9084 = a9082 & a9070;
assign a9086 = ~a7824 & ~l1538;
assign a9088 = a7824 & l1194;
assign a9090 = ~a9088 & ~a9086;
assign a9092 = a9090 & ~i598;
assign a9094 = ~a9090 & i598;
assign a9096 = ~a9094 & ~a9092;
assign a9098 = a9096 & a9084;
assign a9100 = a7824 & ~l1200;
assign a9102 = ~a7824 & ~l1540;
assign a9104 = ~a9102 & ~a9100;
assign a9106 = a9104 & ~i600;
assign a9108 = ~a9104 & i600;
assign a9110 = ~a9108 & ~a9106;
assign a9112 = a9110 & a9098;
assign a9114 = ~a7824 & ~l1542;
assign a9116 = a7824 & l1202;
assign a9118 = ~a9116 & ~a9114;
assign a9120 = a9118 & ~i602;
assign a9122 = ~a9118 & i602;
assign a9124 = ~a9122 & ~a9120;
assign a9126 = a9124 & a9112;
assign a9128 = a7824 & ~l1206;
assign a9130 = ~a7824 & ~l1544;
assign a9132 = ~a9130 & ~a9128;
assign a9134 = a9132 & ~i604;
assign a9136 = ~a9132 & i604;
assign a9138 = ~a9136 & ~a9134;
assign a9140 = a9138 & a9126;
assign a9142 = ~a7824 & ~l1546;
assign a9144 = a7824 & l1208;
assign a9146 = ~a9144 & ~a9142;
assign a9148 = a9146 & ~i606;
assign a9150 = ~a9146 & i606;
assign a9152 = ~a9150 & ~a9148;
assign a9154 = a9152 & a9140;
assign a9156 = a7824 & ~l1214;
assign a9158 = ~a7824 & ~l1548;
assign a9160 = ~a9158 & ~a9156;
assign a9162 = a9160 & ~i608;
assign a9164 = ~a9160 & i608;
assign a9166 = ~a9164 & ~a9162;
assign a9168 = a9166 & a9154;
assign a9170 = ~a7824 & ~l1550;
assign a9172 = a7824 & l1216;
assign a9174 = ~a9172 & ~a9170;
assign a9176 = a9174 & ~i610;
assign a9178 = ~a9174 & i610;
assign a9180 = ~a9178 & ~a9176;
assign a9182 = a9180 & a9168;
assign a9184 = a7824 & ~l1220;
assign a9186 = ~a7824 & ~l1552;
assign a9188 = ~a9186 & ~a9184;
assign a9190 = a9188 & ~i612;
assign a9192 = ~a9188 & i612;
assign a9194 = ~a9192 & ~a9190;
assign a9196 = a9194 & a9182;
assign a9198 = ~a7824 & ~l1554;
assign a9200 = a7824 & l1222;
assign a9202 = ~a9200 & ~a9198;
assign a9204 = a9202 & ~i614;
assign a9206 = ~a9202 & i614;
assign a9208 = ~a9206 & ~a9204;
assign a9210 = a9208 & a9196;
assign a9212 = a7824 & ~l1228;
assign a9214 = ~a7824 & ~l1556;
assign a9216 = ~a9214 & ~a9212;
assign a9218 = a9216 & ~i616;
assign a9220 = ~a9216 & i616;
assign a9222 = ~a9220 & ~a9218;
assign a9224 = a9222 & a9210;
assign a9226 = ~a7824 & ~l1558;
assign a9228 = a7824 & l1230;
assign a9230 = ~a9228 & ~a9226;
assign a9232 = a9230 & ~i618;
assign a9234 = ~a9230 & i618;
assign a9236 = ~a9234 & ~a9232;
assign a9238 = a9236 & a9224;
assign a9240 = a7824 & ~l1234;
assign a9242 = ~a7824 & ~l1560;
assign a9244 = ~a9242 & ~a9240;
assign a9246 = a9244 & ~i620;
assign a9248 = ~a9244 & i620;
assign a9250 = ~a9248 & ~a9246;
assign a9252 = a9250 & a9238;
assign a9254 = ~a7824 & ~l1562;
assign a9256 = a7824 & l1236;
assign a9258 = ~a9256 & ~a9254;
assign a9260 = a9258 & ~i622;
assign a9262 = ~a9258 & i622;
assign a9264 = ~a9262 & ~a9260;
assign a9266 = a9264 & a9252;
assign a9268 = a7824 & ~l1238;
assign a9270 = ~a7824 & ~l1564;
assign a9272 = ~a9270 & ~a9268;
assign a9274 = a9272 & ~i624;
assign a9276 = ~a9272 & i624;
assign a9278 = ~a9276 & ~a9274;
assign a9280 = a9278 & a9266;
assign a9282 = a7824 & ~l1240;
assign a9284 = ~a7824 & ~l1566;
assign a9286 = ~a9284 & ~a9282;
assign a9288 = a9286 & ~i626;
assign a9290 = ~a9286 & i626;
assign a9292 = ~a9290 & ~a9288;
assign a9294 = a9292 & a9280;
assign a9296 = ~a7824 & ~l1568;
assign a9298 = a7824 & l1242;
assign a9300 = ~a9298 & ~a9296;
assign a9302 = a9300 & ~i628;
assign a9304 = ~a9300 & i628;
assign a9306 = ~a9304 & ~a9302;
assign a9308 = a9306 & a9294;
assign a9310 = a7824 & ~l1244;
assign a9312 = ~a7824 & ~l1570;
assign a9314 = ~a9312 & ~a9310;
assign a9316 = a9314 & ~i630;
assign a9318 = ~a9314 & i630;
assign a9320 = ~a9318 & ~a9316;
assign a9322 = a9320 & a9308;
assign a9324 = a7824 & ~l1246;
assign a9326 = ~a7824 & ~l1572;
assign a9328 = ~a9326 & ~a9324;
assign a9330 = a9328 & ~i632;
assign a9332 = ~a9328 & i632;
assign a9334 = ~a9332 & ~a9330;
assign a9336 = a9334 & a9322;
assign a9338 = a7824 & ~l1248;
assign a9340 = ~a7824 & ~l1574;
assign a9342 = ~a9340 & ~a9338;
assign a9344 = a9342 & ~i634;
assign a9346 = ~a9342 & i634;
assign a9348 = ~a9346 & ~a9344;
assign a9350 = a9348 & a9336;
assign a9352 = a7824 & ~l1252;
assign a9354 = ~a7824 & ~l1576;
assign a9356 = ~a9354 & ~a9352;
assign a9358 = a9356 & ~i636;
assign a9360 = ~a9356 & i636;
assign a9362 = ~a9360 & ~a9358;
assign a9364 = a9362 & a9350;
assign a9366 = a7824 & ~l1254;
assign a9368 = ~a7824 & ~l1578;
assign a9370 = ~a9368 & ~a9366;
assign a9372 = a9370 & ~i638;
assign a9374 = ~a9370 & i638;
assign a9376 = ~a9374 & ~a9372;
assign a9378 = a9376 & a9364;
assign a9380 = a7824 & ~l1256;
assign a9382 = ~a7824 & ~l1580;
assign a9384 = ~a9382 & ~a9380;
assign a9386 = a9384 & ~i640;
assign a9388 = ~a9384 & i640;
assign a9390 = ~a9388 & ~a9386;
assign a9392 = a9390 & a9378;
assign a9394 = a7824 & ~l1258;
assign a9396 = ~a7824 & ~l1582;
assign a9398 = ~a9396 & ~a9394;
assign a9400 = a9398 & ~i642;
assign a9402 = ~a9398 & i642;
assign a9404 = ~a9402 & ~a9400;
assign a9406 = a9404 & a9392;
assign a9408 = a7824 & ~l1260;
assign a9410 = ~a7824 & ~l1584;
assign a9412 = ~a9410 & ~a9408;
assign a9414 = a9412 & ~i644;
assign a9416 = ~a9412 & i644;
assign a9418 = ~a9416 & ~a9414;
assign a9420 = a9418 & a9406;
assign a9422 = a7824 & ~l1262;
assign a9424 = ~a7824 & ~l1586;
assign a9426 = ~a9424 & ~a9422;
assign a9428 = a9426 & ~i646;
assign a9430 = ~a9426 & i646;
assign a9432 = ~a9430 & ~a9428;
assign a9434 = a9432 & a9420;
assign a9436 = a7824 & ~l1264;
assign a9438 = ~a7824 & ~l1588;
assign a9440 = ~a9438 & ~a9436;
assign a9442 = a9440 & ~i648;
assign a9444 = ~a9440 & i648;
assign a9446 = ~a9444 & ~a9442;
assign a9448 = a9446 & a9434;
assign a9450 = a7824 & ~l1270;
assign a9452 = ~a7824 & ~l1590;
assign a9454 = ~a9452 & ~a9450;
assign a9456 = a9454 & ~i650;
assign a9458 = ~a9454 & i650;
assign a9460 = ~a9458 & ~a9456;
assign a9462 = a9460 & a9448;
assign a9464 = ~a7824 & ~l1592;
assign a9466 = a7824 & l1272;
assign a9468 = ~a9466 & ~a9464;
assign a9470 = a9468 & ~i652;
assign a9472 = ~a9468 & i652;
assign a9474 = ~a9472 & ~a9470;
assign a9476 = a9474 & a9462;
assign a9478 = a7824 & ~l1276;
assign a9480 = ~a7824 & ~l1594;
assign a9482 = ~a9480 & ~a9478;
assign a9484 = a9482 & ~i654;
assign a9486 = ~a9482 & i654;
assign a9488 = ~a9486 & ~a9484;
assign a9490 = a9488 & a9476;
assign a9492 = ~a7824 & ~l1596;
assign a9494 = a7824 & l1278;
assign a9496 = ~a9494 & ~a9492;
assign a9498 = a9496 & ~i656;
assign a9500 = ~a9496 & i656;
assign a9502 = ~a9500 & ~a9498;
assign a9504 = a9502 & a9490;
assign a9506 = a7824 & ~l1284;
assign a9508 = ~a7824 & ~l1598;
assign a9510 = ~a9508 & ~a9506;
assign a9512 = a9510 & ~i658;
assign a9514 = ~a9510 & i658;
assign a9516 = ~a9514 & ~a9512;
assign a9518 = a9516 & a9504;
assign a9520 = ~a7824 & ~l1600;
assign a9522 = a7824 & l1286;
assign a9524 = ~a9522 & ~a9520;
assign a9526 = a9524 & ~i660;
assign a9528 = ~a9524 & i660;
assign a9530 = ~a9528 & ~a9526;
assign a9532 = a9530 & a9518;
assign a9534 = a7824 & ~l1290;
assign a9536 = ~a7824 & ~l1602;
assign a9538 = ~a9536 & ~a9534;
assign a9540 = a9538 & ~i662;
assign a9542 = ~a9538 & i662;
assign a9544 = ~a9542 & ~a9540;
assign a9546 = a9544 & a9532;
assign a9548 = ~a7824 & ~l1604;
assign a9550 = a7824 & l1292;
assign a9552 = ~a9550 & ~a9548;
assign a9554 = a9552 & ~i664;
assign a9556 = ~a9552 & i664;
assign a9558 = ~a9556 & ~a9554;
assign a9560 = a9558 & a9546;
assign a9562 = a7824 & ~l1298;
assign a9564 = ~a7824 & ~l1606;
assign a9566 = ~a9564 & ~a9562;
assign a9568 = a9566 & ~i666;
assign a9570 = ~a9566 & i666;
assign a9572 = ~a9570 & ~a9568;
assign a9574 = a9572 & a9560;
assign a9576 = ~a7824 & ~l1608;
assign a9578 = a7824 & l1300;
assign a9580 = ~a9578 & ~a9576;
assign a9582 = a9580 & ~i668;
assign a9584 = ~a9580 & i668;
assign a9586 = ~a9584 & ~a9582;
assign a9588 = a9586 & a9574;
assign a9590 = a7824 & ~l1304;
assign a9592 = ~a7824 & ~l1610;
assign a9594 = ~a9592 & ~a9590;
assign a9596 = a9594 & ~i670;
assign a9598 = ~a9594 & i670;
assign a9600 = ~a9598 & ~a9596;
assign a9602 = a9600 & a9588;
assign a9604 = ~a7824 & ~l1612;
assign a9606 = a7824 & l1306;
assign a9608 = ~a9606 & ~a9604;
assign a9610 = a9608 & ~i672;
assign a9612 = ~a9608 & i672;
assign a9614 = ~a9612 & ~a9610;
assign a9616 = a9614 & a9602;
assign a9618 = a7824 & ~l1312;
assign a9620 = ~a7824 & ~l1614;
assign a9622 = ~a9620 & ~a9618;
assign a9624 = a9622 & ~i674;
assign a9626 = ~a9622 & i674;
assign a9628 = ~a9626 & ~a9624;
assign a9630 = a9628 & a9616;
assign a9632 = ~a7824 & ~l1616;
assign a9634 = a7824 & l1314;
assign a9636 = ~a9634 & ~a9632;
assign a9638 = a9636 & ~i676;
assign a9640 = ~a9636 & i676;
assign a9642 = ~a9640 & ~a9638;
assign a9644 = a9642 & a9630;
assign a9646 = a7824 & ~l1318;
assign a9648 = ~a7824 & ~l1618;
assign a9650 = ~a9648 & ~a9646;
assign a9652 = a9650 & ~i678;
assign a9654 = ~a9650 & i678;
assign a9656 = ~a9654 & ~a9652;
assign a9658 = a9656 & a9644;
assign a9660 = ~a7824 & ~l1620;
assign a9662 = a7824 & l1320;
assign a9664 = ~a9662 & ~a9660;
assign a9666 = a9664 & ~i680;
assign a9668 = ~a9664 & i680;
assign a9670 = ~a9668 & ~a9666;
assign a9672 = a9670 & a9658;
assign a9674 = a7824 & ~l1322;
assign a9676 = ~a7824 & ~l1622;
assign a9678 = ~a9676 & ~a9674;
assign a9680 = a9678 & ~i682;
assign a9682 = ~a9678 & i682;
assign a9684 = ~a9682 & ~a9680;
assign a9686 = a9684 & a9672;
assign a9688 = a7824 & ~l1324;
assign a9690 = ~a7824 & ~l1624;
assign a9692 = ~a9690 & ~a9688;
assign a9694 = a9692 & ~i684;
assign a9696 = ~a9692 & i684;
assign a9698 = ~a9696 & ~a9694;
assign a9700 = a9698 & a9686;
assign a9702 = ~a7824 & ~l1626;
assign a9704 = a7824 & l1326;
assign a9706 = ~a9704 & ~a9702;
assign a9708 = a9706 & ~i686;
assign a9710 = ~a9706 & i686;
assign a9712 = ~a9710 & ~a9708;
assign a9714 = a9712 & a9700;
assign a9716 = a7824 & ~l1328;
assign a9718 = ~a7824 & ~l1628;
assign a9720 = ~a9718 & ~a9716;
assign a9722 = a9720 & ~i688;
assign a9724 = ~a9720 & i688;
assign a9726 = ~a9724 & ~a9722;
assign a9728 = a9726 & a9714;
assign a9730 = a7824 & ~l1330;
assign a9732 = ~a7824 & ~l1630;
assign a9734 = ~a9732 & ~a9730;
assign a9736 = a9734 & ~i690;
assign a9738 = ~a9734 & i690;
assign a9740 = ~a9738 & ~a9736;
assign a9742 = a9740 & a9728;
assign a9744 = a7824 & ~l1332;
assign a9746 = ~a7824 & ~l1632;
assign a9748 = ~a9746 & ~a9744;
assign a9750 = a9748 & ~i692;
assign a9752 = ~a9748 & i692;
assign a9754 = ~a9752 & ~a9750;
assign a9756 = a9754 & a9742;
assign a9758 = a7824 & ~l1336;
assign a9760 = ~a7824 & ~l1634;
assign a9762 = ~a9760 & ~a9758;
assign a9764 = a9762 & ~i694;
assign a9766 = ~a9762 & i694;
assign a9768 = ~a9766 & ~a9764;
assign a9770 = a9768 & a9756;
assign a9772 = a7824 & ~l1338;
assign a9774 = ~a7824 & ~l1636;
assign a9776 = ~a9774 & ~a9772;
assign a9778 = a9776 & ~i696;
assign a9780 = ~a9776 & i696;
assign a9782 = ~a9780 & ~a9778;
assign a9784 = a9782 & a9770;
assign a9786 = a7824 & ~l1340;
assign a9788 = ~a7824 & ~l1638;
assign a9790 = ~a9788 & ~a9786;
assign a9792 = a9790 & ~i698;
assign a9794 = ~a9790 & i698;
assign a9796 = ~a9794 & ~a9792;
assign a9798 = a9796 & a9784;
assign a9800 = a7824 & ~l1342;
assign a9802 = ~a7824 & ~l1640;
assign a9804 = ~a9802 & ~a9800;
assign a9806 = a9804 & ~i700;
assign a9808 = ~a9804 & i700;
assign a9810 = ~a9808 & ~a9806;
assign a9812 = a9810 & a9798;
assign a9814 = a7824 & ~l1344;
assign a9816 = ~a7824 & ~l1642;
assign a9818 = ~a9816 & ~a9814;
assign a9820 = a9818 & ~i702;
assign a9822 = ~a9818 & i702;
assign a9824 = ~a9822 & ~a9820;
assign a9826 = a9824 & a9812;
assign a9828 = a7824 & ~l1346;
assign a9830 = ~a7824 & ~l1644;
assign a9832 = ~a9830 & ~a9828;
assign a9834 = a9832 & ~i704;
assign a9836 = ~a9832 & i704;
assign a9838 = ~a9836 & ~a9834;
assign a9840 = a9838 & a9826;
assign a9842 = a7824 & ~l1348;
assign a9844 = ~a7824 & ~l1646;
assign a9846 = ~a9844 & ~a9842;
assign a9848 = a9846 & ~i706;
assign a9850 = ~a9846 & i706;
assign a9852 = ~a9850 & ~a9848;
assign a9854 = a9852 & a9840;
assign a9856 = a7824 & ~l1350;
assign a9858 = ~a7824 & ~l1648;
assign a9860 = ~a9858 & ~a9856;
assign a9862 = a9860 & ~i708;
assign a9864 = ~a9860 & i708;
assign a9866 = ~a9864 & ~a9862;
assign a9868 = a9866 & a9854;
assign a9870 = a7824 & ~l1352;
assign a9872 = ~a7824 & ~l1650;
assign a9874 = ~a9872 & ~a9870;
assign a9876 = a9874 & ~i710;
assign a9878 = ~a9874 & i710;
assign a9880 = ~a9878 & ~a9876;
assign a9882 = a9880 & a9868;
assign a9884 = a7824 & ~l1354;
assign a9886 = ~a7824 & ~l1652;
assign a9888 = ~a9886 & ~a9884;
assign a9890 = a9888 & ~i712;
assign a9892 = ~a9888 & i712;
assign a9894 = ~a9892 & ~a9890;
assign a9896 = a9894 & a9882;
assign a9898 = a7824 & ~l1356;
assign a9900 = ~a7824 & ~l1654;
assign a9902 = ~a9900 & ~a9898;
assign a9904 = a9902 & ~i714;
assign a9906 = ~a9902 & i714;
assign a9908 = ~a9906 & ~a9904;
assign a9910 = a9908 & a9896;
assign a9912 = l732 & l730;
assign a9914 = l742 & l740;
assign a9916 = l752 & l750;
assign a9918 = l762 & l760;
assign a9920 = l772 & l770;
assign a9922 = l782 & l780;
assign a9924 = l792 & l790;
assign a9926 = l802 & l800;
assign a9928 = l812 & l810;
assign a9930 = l822 & l820;
assign a9932 = l832 & l830;
assign a9934 = l842 & l840;
assign a9936 = l852 & l850;
assign a9938 = l862 & l860;
assign a9940 = l872 & l870;
assign a9942 = l882 & l880;
assign a9944 = l892 & l890;
assign a9946 = l902 & l900;
assign a9948 = l912 & l910;
assign a9950 = l922 & l920;
assign a9952 = l932 & l930;
assign a9954 = ~l936 & l934;
assign a9956 = l946 & l944;
assign a9958 = ~l950 & l948;
assign a9960 = l960 & l958;
assign a9962 = ~l964 & l962;
assign a9964 = l974 & l972;
assign a9966 = ~l978 & l976;
assign a9968 = a1764 & l986;
assign a9970 = a2024 & ~l1006;
assign a9972 = ~a9970 & l1004;
assign a9974 = l1016 & l1014;
assign a9976 = ~l1020 & l1018;
assign a9978 = l1030 & l1028;
assign a9980 = ~l1034 & l1032;
assign a9982 = l1044 & l1042;
assign a9984 = ~l1048 & l1046;
assign a9986 = l1058 & l1056;
assign a9988 = ~l1062 & l1060;
assign a9990 = a2650 & l1070;
assign a9992 = a2910 & ~l1090;
assign a9994 = ~a9992 & l1088;
assign a9996 = l1100 & l1098;
assign a9998 = ~l1104 & l1102;
assign a10000 = l1114 & l1112;
assign a10002 = ~l1118 & l1116;
assign a10004 = l1128 & l1126;
assign a10006 = ~l1132 & l1130;
assign a10008 = l1142 & l1140;
assign a10010 = ~l1146 & l1144;
assign a10012 = a3536 & l1154;
assign a10014 = a3796 & ~l1174;
assign a10016 = ~a10014 & l1172;
assign a10018 = l1184 & l1182;
assign a10020 = ~l1188 & l1186;
assign a10022 = l1198 & l1196;
assign a10024 = ~l1202 & l1200;
assign a10026 = l1212 & l1210;
assign a10028 = ~l1216 & l1214;
assign a10030 = l1226 & l1224;
assign a10032 = ~l1230 & l1228;
assign a10034 = a4422 & l1238;
assign a10036 = a4682 & ~l1258;
assign a10038 = ~a10036 & l1256;
assign a10040 = l1268 & l1266;
assign a10042 = ~l1272 & l1270;
assign a10044 = l1282 & l1280;
assign a10046 = ~l1286 & l1284;
assign a10048 = l1296 & l1294;
assign a10050 = ~l1300 & l1298;
assign a10052 = l1310 & l1308;
assign a10054 = ~l1314 & l1312;
assign a10056 = a5308 & l1322;
assign a10058 = a5568 & ~l1342;
assign a10060 = ~a10058 & l1340;
assign a10062 = l1360 & l1358;
assign a10064 = l1368 & l1366;
assign a10066 = l1376 & l1374;
assign a10068 = l1384 & l1382;
assign a10070 = l1394 & l1392;
assign a10072 = a10070 & l1390;
assign a10074 = l1414 & l1412;
assign a10076 = ~a10074 & ~l1410;
assign a10078 = a10076 & ~l1408;
assign a10080 = ~a10078 & l1406;
assign a10082 = l1418 & l1416;
assign a10084 = l1426 & l1424;
assign a10086 = l1434 & l1432;
assign a10088 = l1442 & l1440;
assign a10090 = l1452 & l1450;
assign a10092 = a10090 & l1448;
assign a10094 = l1472 & l1470;
assign a10096 = ~a10094 & ~l1468;
assign a10098 = a10096 & ~l1466;
assign a10100 = ~a10098 & l1464;
assign a10102 = l1476 & l1474;
assign a10104 = l1484 & l1482;
assign a10106 = l1492 & l1490;
assign a10108 = l1500 & l1498;
assign a10110 = l1510 & l1508;
assign a10112 = a10110 & l1506;
assign a10114 = l1530 & l1528;
assign a10116 = ~a10114 & ~l1526;
assign a10118 = a10116 & ~l1524;
assign a10120 = ~a10118 & l1522;
assign a10122 = l1534 & l1532;
assign a10124 = l1542 & l1540;
assign a10126 = l1550 & l1548;
assign a10128 = l1558 & l1556;
assign a10130 = l1568 & l1566;
assign a10132 = a10130 & l1564;
assign a10134 = l1588 & l1586;
assign a10136 = ~a10134 & ~l1584;
assign a10138 = a10136 & ~l1582;
assign a10140 = ~a10138 & l1580;
assign a10142 = l1592 & l1590;
assign a10144 = l1600 & l1598;
assign a10146 = l1608 & l1606;
assign a10148 = l1616 & l1614;
assign a10150 = l1626 & l1624;
assign a10152 = a10150 & l1622;
assign a10154 = l1646 & l1644;
assign a10156 = ~a10154 & ~l1642;
assign a10158 = a10156 & ~l1640;
assign a10160 = ~a10158 & l1638;
assign a10162 = ~l1168 & ~l1084;
assign a10164 = l1168 & l1084;
assign a10166 = ~a10164 & ~a10162;
assign a10168 = a3466 & a2580;
assign a10170 = a10168 & ~a10166;
assign a10172 = ~l1084 & ~l1000;
assign a10174 = l1084 & l1000;
assign a10176 = ~a10174 & ~a10172;
assign a10178 = ~a10176 & a2580;
assign a10180 = ~l1168 & ~l1000;
assign a10182 = l1168 & l1000;
assign a10184 = ~a10182 & ~a10180;
assign a10186 = ~a10184 & a3466;
assign a10188 = ~l1252 & ~l1000;
assign a10190 = l1252 & l1000;
assign a10192 = ~a10190 & ~a10188;
assign a10194 = ~a10192 & a4352;
assign a10196 = ~l1336 & ~l1000;
assign a10198 = l1336 & l1000;
assign a10200 = ~a10198 & ~a10196;
assign a10202 = ~a10200 & a5238;
assign a10204 = ~a10202 & ~a10194;
assign a10206 = a10204 & ~a10186;
assign a10208 = a10206 & ~a10178;
assign a10210 = ~a10208 & a1694;
assign a10212 = ~l1252 & ~l1084;
assign a10214 = l1252 & l1084;
assign a10216 = ~a10214 & ~a10212;
assign a10218 = a4352 & a2580;
assign a10220 = a10218 & ~a10216;
assign a10222 = ~l1336 & ~l1084;
assign a10224 = l1336 & l1084;
assign a10226 = ~a10224 & ~a10222;
assign a10228 = a5238 & a2580;
assign a10230 = a10228 & ~a10226;
assign a10232 = ~l1252 & ~l1168;
assign a10234 = l1252 & l1168;
assign a10236 = ~a10234 & ~a10232;
assign a10238 = a4352 & a3466;
assign a10240 = a10238 & ~a10236;
assign a10242 = ~l1336 & ~l1168;
assign a10244 = l1336 & l1168;
assign a10246 = ~a10244 & ~a10242;
assign a10248 = a5238 & a3466;
assign a10250 = a10248 & ~a10246;
assign a10252 = ~l1336 & ~l1252;
assign a10254 = l1336 & l1252;
assign a10256 = ~a10254 & ~a10252;
assign a10258 = a5238 & a4352;
assign a10260 = a10258 & ~a10256;
assign a10262 = ~a10260 & ~a10250;
assign a10264 = a10262 & ~a10240;
assign a10266 = a10264 & ~a10230;
assign a10268 = a10266 & ~a10220;
assign a10270 = a10268 & ~a10210;
assign a10272 = a10270 & ~a10170;
assign a10274 = ~a10272 & l1350;
assign a10276 = ~l734 & ~l732;
assign a10278 = a10276 & ~l730;
assign a10280 = l734 & ~l732;
assign a10282 = a10280 & ~l730;
assign a10284 = ~l734 & l732;
assign a10286 = a10284 & ~l730;
assign a10288 = l734 & l732;
assign a10290 = a10288 & ~l730;
assign a10292 = a10276 & l730;
assign a10294 = a10280 & l730;
assign a10296 = ~l738 & ~l736;
assign a10298 = l738 & ~l736;
assign a10300 = ~l738 & l736;
assign a10302 = l738 & l736;
assign a10304 = a10302 & ~l1312;
assign a10306 = a10304 & ~a10300;
assign a10308 = a10300 & ~l1298;
assign a10310 = ~a10308 & ~a10306;
assign a10312 = ~a10310 & ~a10298;
assign a10314 = a10298 & ~l1284;
assign a10316 = ~a10314 & ~a10312;
assign a10318 = ~a10316 & ~a10296;
assign a10320 = a10296 & ~l1270;
assign a10322 = ~a10320 & ~a10318;
assign a10324 = ~a10322 & a10294;
assign a10326 = a10324 & ~a10292;
assign a10328 = a10302 & ~l1228;
assign a10330 = a10328 & ~a10300;
assign a10332 = a10300 & ~l1214;
assign a10334 = ~a10332 & ~a10330;
assign a10336 = ~a10334 & ~a10298;
assign a10338 = a10298 & ~l1200;
assign a10340 = ~a10338 & ~a10336;
assign a10342 = ~a10340 & ~a10296;
assign a10344 = a10296 & ~l1186;
assign a10346 = ~a10344 & ~a10342;
assign a10348 = ~a10346 & a10292;
assign a10350 = ~a10348 & ~a10326;
assign a10352 = ~a10350 & ~a10290;
assign a10354 = a10302 & ~l1144;
assign a10356 = a10354 & ~a10300;
assign a10358 = a10300 & ~l1130;
assign a10360 = ~a10358 & ~a10356;
assign a10362 = ~a10360 & ~a10298;
assign a10364 = a10298 & ~l1116;
assign a10366 = ~a10364 & ~a10362;
assign a10368 = ~a10366 & ~a10296;
assign a10370 = a10296 & ~l1102;
assign a10372 = ~a10370 & ~a10368;
assign a10374 = ~a10372 & a10290;
assign a10376 = ~a10374 & ~a10352;
assign a10378 = ~a10376 & ~a10286;
assign a10380 = a10302 & ~l1060;
assign a10382 = a10380 & ~a10300;
assign a10384 = a10300 & ~l1046;
assign a10386 = ~a10384 & ~a10382;
assign a10388 = ~a10386 & ~a10298;
assign a10390 = a10298 & ~l1032;
assign a10392 = ~a10390 & ~a10388;
assign a10394 = ~a10392 & ~a10296;
assign a10396 = a10296 & ~l1018;
assign a10398 = ~a10396 & ~a10394;
assign a10400 = ~a10398 & a10286;
assign a10402 = ~a10400 & ~a10378;
assign a10404 = ~a10402 & ~a10282;
assign a10406 = a10302 & ~l976;
assign a10408 = a10406 & ~a10300;
assign a10410 = a10300 & ~l962;
assign a10412 = ~a10410 & ~a10408;
assign a10414 = ~a10412 & ~a10298;
assign a10416 = a10298 & ~l948;
assign a10418 = ~a10416 & ~a10414;
assign a10420 = ~a10418 & ~a10296;
assign a10422 = a10296 & ~l934;
assign a10424 = ~a10422 & ~a10420;
assign a10426 = ~a10424 & a10282;
assign a10428 = ~a10426 & ~a10404;
assign a10430 = a10428 & ~l930;
assign a10432 = ~a10428 & l930;
assign a10434 = ~a10432 & ~a10430;
assign a10436 = a10302 & l1314;
assign a10438 = a10436 & ~a10300;
assign a10440 = a10300 & l1300;
assign a10442 = ~a10440 & ~a10438;
assign a10444 = ~a10442 & ~a10298;
assign a10446 = a10298 & l1286;
assign a10448 = ~a10446 & ~a10444;
assign a10450 = ~a10448 & ~a10296;
assign a10452 = a10296 & l1272;
assign a10454 = ~a10452 & ~a10450;
assign a10456 = ~a10454 & a10294;
assign a10458 = a10456 & ~a10292;
assign a10460 = a10302 & l1230;
assign a10462 = a10460 & ~a10300;
assign a10464 = a10300 & l1216;
assign a10466 = ~a10464 & ~a10462;
assign a10468 = ~a10466 & ~a10298;
assign a10470 = a10298 & l1202;
assign a10472 = ~a10470 & ~a10468;
assign a10474 = ~a10472 & ~a10296;
assign a10476 = a10296 & l1188;
assign a10478 = ~a10476 & ~a10474;
assign a10480 = ~a10478 & a10292;
assign a10482 = ~a10480 & ~a10458;
assign a10484 = ~a10482 & ~a10290;
assign a10486 = a10302 & l1146;
assign a10488 = a10486 & ~a10300;
assign a10490 = a10300 & l1132;
assign a10492 = ~a10490 & ~a10488;
assign a10494 = ~a10492 & ~a10298;
assign a10496 = a10298 & l1118;
assign a10498 = ~a10496 & ~a10494;
assign a10500 = ~a10498 & ~a10296;
assign a10502 = a10296 & l1104;
assign a10504 = ~a10502 & ~a10500;
assign a10506 = ~a10504 & a10290;
assign a10508 = ~a10506 & ~a10484;
assign a10510 = ~a10508 & ~a10286;
assign a10512 = a10302 & l1062;
assign a10514 = a10512 & ~a10300;
assign a10516 = a10300 & l1048;
assign a10518 = ~a10516 & ~a10514;
assign a10520 = ~a10518 & ~a10298;
assign a10522 = a10298 & l1034;
assign a10524 = ~a10522 & ~a10520;
assign a10526 = ~a10524 & ~a10296;
assign a10528 = a10296 & l1020;
assign a10530 = ~a10528 & ~a10526;
assign a10532 = ~a10530 & a10286;
assign a10534 = ~a10532 & ~a10510;
assign a10536 = ~a10534 & ~a10282;
assign a10538 = a10302 & l978;
assign a10540 = a10538 & ~a10300;
assign a10542 = a10300 & l964;
assign a10544 = ~a10542 & ~a10540;
assign a10546 = ~a10544 & ~a10298;
assign a10548 = a10298 & l950;
assign a10550 = ~a10548 & ~a10546;
assign a10552 = ~a10550 & ~a10296;
assign a10554 = a10296 & l936;
assign a10556 = ~a10554 & ~a10552;
assign a10558 = ~a10556 & a10282;
assign a10560 = ~a10558 & ~a10536;
assign a10562 = a10560 & ~l932;
assign a10564 = ~a10560 & l932;
assign a10566 = ~a10564 & ~a10562;
assign a10568 = a10566 & a10434;
assign a10570 = ~a10568 & ~a10278;
assign a10572 = ~l744 & ~l742;
assign a10574 = a10572 & ~l740;
assign a10576 = l744 & ~l742;
assign a10578 = a10576 & ~l740;
assign a10580 = ~l744 & l742;
assign a10582 = a10580 & ~l740;
assign a10584 = l744 & l742;
assign a10586 = a10584 & ~l740;
assign a10588 = a10572 & l740;
assign a10590 = a10576 & l740;
assign a10592 = ~l748 & ~l746;
assign a10594 = l748 & ~l746;
assign a10596 = ~l748 & l746;
assign a10598 = l748 & l746;
assign a10600 = a10598 & ~l1312;
assign a10602 = a10600 & ~a10596;
assign a10604 = a10596 & ~l1298;
assign a10606 = ~a10604 & ~a10602;
assign a10608 = ~a10606 & ~a10594;
assign a10610 = a10594 & ~l1284;
assign a10612 = ~a10610 & ~a10608;
assign a10614 = ~a10612 & ~a10592;
assign a10616 = a10592 & ~l1270;
assign a10618 = ~a10616 & ~a10614;
assign a10620 = ~a10618 & a10590;
assign a10622 = a10620 & ~a10588;
assign a10624 = a10598 & ~l1228;
assign a10626 = a10624 & ~a10596;
assign a10628 = a10596 & ~l1214;
assign a10630 = ~a10628 & ~a10626;
assign a10632 = ~a10630 & ~a10594;
assign a10634 = a10594 & ~l1200;
assign a10636 = ~a10634 & ~a10632;
assign a10638 = ~a10636 & ~a10592;
assign a10640 = a10592 & ~l1186;
assign a10642 = ~a10640 & ~a10638;
assign a10644 = ~a10642 & a10588;
assign a10646 = ~a10644 & ~a10622;
assign a10648 = ~a10646 & ~a10586;
assign a10650 = a10598 & ~l1144;
assign a10652 = a10650 & ~a10596;
assign a10654 = a10596 & ~l1130;
assign a10656 = ~a10654 & ~a10652;
assign a10658 = ~a10656 & ~a10594;
assign a10660 = a10594 & ~l1116;
assign a10662 = ~a10660 & ~a10658;
assign a10664 = ~a10662 & ~a10592;
assign a10666 = a10592 & ~l1102;
assign a10668 = ~a10666 & ~a10664;
assign a10670 = ~a10668 & a10586;
assign a10672 = ~a10670 & ~a10648;
assign a10674 = ~a10672 & ~a10582;
assign a10676 = a10598 & ~l1060;
assign a10678 = a10676 & ~a10596;
assign a10680 = a10596 & ~l1046;
assign a10682 = ~a10680 & ~a10678;
assign a10684 = ~a10682 & ~a10594;
assign a10686 = a10594 & ~l1032;
assign a10688 = ~a10686 & ~a10684;
assign a10690 = ~a10688 & ~a10592;
assign a10692 = a10592 & ~l1018;
assign a10694 = ~a10692 & ~a10690;
assign a10696 = ~a10694 & a10582;
assign a10698 = ~a10696 & ~a10674;
assign a10700 = ~a10698 & ~a10578;
assign a10702 = a10598 & ~l976;
assign a10704 = a10702 & ~a10596;
assign a10706 = a10596 & ~l962;
assign a10708 = ~a10706 & ~a10704;
assign a10710 = ~a10708 & ~a10594;
assign a10712 = a10594 & ~l948;
assign a10714 = ~a10712 & ~a10710;
assign a10716 = ~a10714 & ~a10592;
assign a10718 = a10592 & ~l934;
assign a10720 = ~a10718 & ~a10716;
assign a10722 = ~a10720 & a10578;
assign a10724 = ~a10722 & ~a10700;
assign a10726 = a10724 & ~l944;
assign a10728 = ~a10724 & l944;
assign a10730 = ~a10728 & ~a10726;
assign a10732 = a10598 & l1314;
assign a10734 = a10732 & ~a10596;
assign a10736 = a10596 & l1300;
assign a10738 = ~a10736 & ~a10734;
assign a10740 = ~a10738 & ~a10594;
assign a10742 = a10594 & l1286;
assign a10744 = ~a10742 & ~a10740;
assign a10746 = ~a10744 & ~a10592;
assign a10748 = a10592 & l1272;
assign a10750 = ~a10748 & ~a10746;
assign a10752 = ~a10750 & a10590;
assign a10754 = a10752 & ~a10588;
assign a10756 = a10598 & l1230;
assign a10758 = a10756 & ~a10596;
assign a10760 = a10596 & l1216;
assign a10762 = ~a10760 & ~a10758;
assign a10764 = ~a10762 & ~a10594;
assign a10766 = a10594 & l1202;
assign a10768 = ~a10766 & ~a10764;
assign a10770 = ~a10768 & ~a10592;
assign a10772 = a10592 & l1188;
assign a10774 = ~a10772 & ~a10770;
assign a10776 = ~a10774 & a10588;
assign a10778 = ~a10776 & ~a10754;
assign a10780 = ~a10778 & ~a10586;
assign a10782 = a10598 & l1146;
assign a10784 = a10782 & ~a10596;
assign a10786 = a10596 & l1132;
assign a10788 = ~a10786 & ~a10784;
assign a10790 = ~a10788 & ~a10594;
assign a10792 = a10594 & l1118;
assign a10794 = ~a10792 & ~a10790;
assign a10796 = ~a10794 & ~a10592;
assign a10798 = a10592 & l1104;
assign a10800 = ~a10798 & ~a10796;
assign a10802 = ~a10800 & a10586;
assign a10804 = ~a10802 & ~a10780;
assign a10806 = ~a10804 & ~a10582;
assign a10808 = a10598 & l1062;
assign a10810 = a10808 & ~a10596;
assign a10812 = a10596 & l1048;
assign a10814 = ~a10812 & ~a10810;
assign a10816 = ~a10814 & ~a10594;
assign a10818 = a10594 & l1034;
assign a10820 = ~a10818 & ~a10816;
assign a10822 = ~a10820 & ~a10592;
assign a10824 = a10592 & l1020;
assign a10826 = ~a10824 & ~a10822;
assign a10828 = ~a10826 & a10582;
assign a10830 = ~a10828 & ~a10806;
assign a10832 = ~a10830 & ~a10578;
assign a10834 = a10598 & l978;
assign a10836 = a10834 & ~a10596;
assign a10838 = a10596 & l964;
assign a10840 = ~a10838 & ~a10836;
assign a10842 = ~a10840 & ~a10594;
assign a10844 = a10594 & l950;
assign a10846 = ~a10844 & ~a10842;
assign a10848 = ~a10846 & ~a10592;
assign a10850 = a10592 & l936;
assign a10852 = ~a10850 & ~a10848;
assign a10854 = ~a10852 & a10578;
assign a10856 = ~a10854 & ~a10832;
assign a10858 = a10856 & ~l946;
assign a10860 = ~a10856 & l946;
assign a10862 = ~a10860 & ~a10858;
assign a10864 = a10862 & a10730;
assign a10866 = ~a10864 & ~a10574;
assign a10868 = ~l754 & ~l752;
assign a10870 = a10868 & ~l750;
assign a10872 = l754 & ~l752;
assign a10874 = a10872 & ~l750;
assign a10876 = ~l754 & l752;
assign a10878 = a10876 & ~l750;
assign a10880 = l754 & l752;
assign a10882 = a10880 & ~l750;
assign a10884 = a10868 & l750;
assign a10886 = a10872 & l750;
assign a10888 = ~l758 & ~l756;
assign a10890 = l758 & ~l756;
assign a10892 = ~l758 & l756;
assign a10894 = l758 & l756;
assign a10896 = a10894 & ~l1312;
assign a10898 = a10896 & ~a10892;
assign a10900 = a10892 & ~l1298;
assign a10902 = ~a10900 & ~a10898;
assign a10904 = ~a10902 & ~a10890;
assign a10906 = a10890 & ~l1284;
assign a10908 = ~a10906 & ~a10904;
assign a10910 = ~a10908 & ~a10888;
assign a10912 = a10888 & ~l1270;
assign a10914 = ~a10912 & ~a10910;
assign a10916 = ~a10914 & a10886;
assign a10918 = a10916 & ~a10884;
assign a10920 = a10894 & ~l1228;
assign a10922 = a10920 & ~a10892;
assign a10924 = a10892 & ~l1214;
assign a10926 = ~a10924 & ~a10922;
assign a10928 = ~a10926 & ~a10890;
assign a10930 = a10890 & ~l1200;
assign a10932 = ~a10930 & ~a10928;
assign a10934 = ~a10932 & ~a10888;
assign a10936 = a10888 & ~l1186;
assign a10938 = ~a10936 & ~a10934;
assign a10940 = ~a10938 & a10884;
assign a10942 = ~a10940 & ~a10918;
assign a10944 = ~a10942 & ~a10882;
assign a10946 = a10894 & ~l1144;
assign a10948 = a10946 & ~a10892;
assign a10950 = a10892 & ~l1130;
assign a10952 = ~a10950 & ~a10948;
assign a10954 = ~a10952 & ~a10890;
assign a10956 = a10890 & ~l1116;
assign a10958 = ~a10956 & ~a10954;
assign a10960 = ~a10958 & ~a10888;
assign a10962 = a10888 & ~l1102;
assign a10964 = ~a10962 & ~a10960;
assign a10966 = ~a10964 & a10882;
assign a10968 = ~a10966 & ~a10944;
assign a10970 = ~a10968 & ~a10878;
assign a10972 = a10894 & ~l1060;
assign a10974 = a10972 & ~a10892;
assign a10976 = a10892 & ~l1046;
assign a10978 = ~a10976 & ~a10974;
assign a10980 = ~a10978 & ~a10890;
assign a10982 = a10890 & ~l1032;
assign a10984 = ~a10982 & ~a10980;
assign a10986 = ~a10984 & ~a10888;
assign a10988 = a10888 & ~l1018;
assign a10990 = ~a10988 & ~a10986;
assign a10992 = ~a10990 & a10878;
assign a10994 = ~a10992 & ~a10970;
assign a10996 = ~a10994 & ~a10874;
assign a10998 = a10894 & ~l976;
assign a11000 = a10998 & ~a10892;
assign a11002 = a10892 & ~l962;
assign a11004 = ~a11002 & ~a11000;
assign a11006 = ~a11004 & ~a10890;
assign a11008 = a10890 & ~l948;
assign a11010 = ~a11008 & ~a11006;
assign a11012 = ~a11010 & ~a10888;
assign a11014 = a10888 & ~l934;
assign a11016 = ~a11014 & ~a11012;
assign a11018 = ~a11016 & a10874;
assign a11020 = ~a11018 & ~a10996;
assign a11022 = a11020 & ~l958;
assign a11024 = ~a11020 & l958;
assign a11026 = ~a11024 & ~a11022;
assign a11028 = a10894 & l1314;
assign a11030 = a11028 & ~a10892;
assign a11032 = a10892 & l1300;
assign a11034 = ~a11032 & ~a11030;
assign a11036 = ~a11034 & ~a10890;
assign a11038 = a10890 & l1286;
assign a11040 = ~a11038 & ~a11036;
assign a11042 = ~a11040 & ~a10888;
assign a11044 = a10888 & l1272;
assign a11046 = ~a11044 & ~a11042;
assign a11048 = ~a11046 & a10886;
assign a11050 = a11048 & ~a10884;
assign a11052 = a10894 & l1230;
assign a11054 = a11052 & ~a10892;
assign a11056 = a10892 & l1216;
assign a11058 = ~a11056 & ~a11054;
assign a11060 = ~a11058 & ~a10890;
assign a11062 = a10890 & l1202;
assign a11064 = ~a11062 & ~a11060;
assign a11066 = ~a11064 & ~a10888;
assign a11068 = a10888 & l1188;
assign a11070 = ~a11068 & ~a11066;
assign a11072 = ~a11070 & a10884;
assign a11074 = ~a11072 & ~a11050;
assign a11076 = ~a11074 & ~a10882;
assign a11078 = a10894 & l1146;
assign a11080 = a11078 & ~a10892;
assign a11082 = a10892 & l1132;
assign a11084 = ~a11082 & ~a11080;
assign a11086 = ~a11084 & ~a10890;
assign a11088 = a10890 & l1118;
assign a11090 = ~a11088 & ~a11086;
assign a11092 = ~a11090 & ~a10888;
assign a11094 = a10888 & l1104;
assign a11096 = ~a11094 & ~a11092;
assign a11098 = ~a11096 & a10882;
assign a11100 = ~a11098 & ~a11076;
assign a11102 = ~a11100 & ~a10878;
assign a11104 = a10894 & l1062;
assign a11106 = a11104 & ~a10892;
assign a11108 = a10892 & l1048;
assign a11110 = ~a11108 & ~a11106;
assign a11112 = ~a11110 & ~a10890;
assign a11114 = a10890 & l1034;
assign a11116 = ~a11114 & ~a11112;
assign a11118 = ~a11116 & ~a10888;
assign a11120 = a10888 & l1020;
assign a11122 = ~a11120 & ~a11118;
assign a11124 = ~a11122 & a10878;
assign a11126 = ~a11124 & ~a11102;
assign a11128 = ~a11126 & ~a10874;
assign a11130 = a10894 & l978;
assign a11132 = a11130 & ~a10892;
assign a11134 = a10892 & l964;
assign a11136 = ~a11134 & ~a11132;
assign a11138 = ~a11136 & ~a10890;
assign a11140 = a10890 & l950;
assign a11142 = ~a11140 & ~a11138;
assign a11144 = ~a11142 & ~a10888;
assign a11146 = a10888 & l936;
assign a11148 = ~a11146 & ~a11144;
assign a11150 = ~a11148 & a10874;
assign a11152 = ~a11150 & ~a11128;
assign a11154 = a11152 & ~l960;
assign a11156 = ~a11152 & l960;
assign a11158 = ~a11156 & ~a11154;
assign a11160 = a11158 & a11026;
assign a11162 = ~a11160 & ~a10870;
assign a11164 = ~l764 & ~l762;
assign a11166 = a11164 & ~l760;
assign a11168 = l764 & ~l762;
assign a11170 = a11168 & ~l760;
assign a11172 = ~l764 & l762;
assign a11174 = a11172 & ~l760;
assign a11176 = l764 & l762;
assign a11178 = a11176 & ~l760;
assign a11180 = a11164 & l760;
assign a11182 = a11168 & l760;
assign a11184 = ~l768 & ~l766;
assign a11186 = l768 & ~l766;
assign a11188 = ~l768 & l766;
assign a11190 = l768 & l766;
assign a11192 = a11190 & ~l1312;
assign a11194 = a11192 & ~a11188;
assign a11196 = a11188 & ~l1298;
assign a11198 = ~a11196 & ~a11194;
assign a11200 = ~a11198 & ~a11186;
assign a11202 = a11186 & ~l1284;
assign a11204 = ~a11202 & ~a11200;
assign a11206 = ~a11204 & ~a11184;
assign a11208 = a11184 & ~l1270;
assign a11210 = ~a11208 & ~a11206;
assign a11212 = ~a11210 & a11182;
assign a11214 = a11212 & ~a11180;
assign a11216 = a11190 & ~l1228;
assign a11218 = a11216 & ~a11188;
assign a11220 = a11188 & ~l1214;
assign a11222 = ~a11220 & ~a11218;
assign a11224 = ~a11222 & ~a11186;
assign a11226 = a11186 & ~l1200;
assign a11228 = ~a11226 & ~a11224;
assign a11230 = ~a11228 & ~a11184;
assign a11232 = a11184 & ~l1186;
assign a11234 = ~a11232 & ~a11230;
assign a11236 = ~a11234 & a11180;
assign a11238 = ~a11236 & ~a11214;
assign a11240 = ~a11238 & ~a11178;
assign a11242 = a11190 & ~l1144;
assign a11244 = a11242 & ~a11188;
assign a11246 = a11188 & ~l1130;
assign a11248 = ~a11246 & ~a11244;
assign a11250 = ~a11248 & ~a11186;
assign a11252 = a11186 & ~l1116;
assign a11254 = ~a11252 & ~a11250;
assign a11256 = ~a11254 & ~a11184;
assign a11258 = a11184 & ~l1102;
assign a11260 = ~a11258 & ~a11256;
assign a11262 = ~a11260 & a11178;
assign a11264 = ~a11262 & ~a11240;
assign a11266 = ~a11264 & ~a11174;
assign a11268 = a11190 & ~l1060;
assign a11270 = a11268 & ~a11188;
assign a11272 = a11188 & ~l1046;
assign a11274 = ~a11272 & ~a11270;
assign a11276 = ~a11274 & ~a11186;
assign a11278 = a11186 & ~l1032;
assign a11280 = ~a11278 & ~a11276;
assign a11282 = ~a11280 & ~a11184;
assign a11284 = a11184 & ~l1018;
assign a11286 = ~a11284 & ~a11282;
assign a11288 = ~a11286 & a11174;
assign a11290 = ~a11288 & ~a11266;
assign a11292 = ~a11290 & ~a11170;
assign a11294 = a11190 & ~l976;
assign a11296 = a11294 & ~a11188;
assign a11298 = a11188 & ~l962;
assign a11300 = ~a11298 & ~a11296;
assign a11302 = ~a11300 & ~a11186;
assign a11304 = a11186 & ~l948;
assign a11306 = ~a11304 & ~a11302;
assign a11308 = ~a11306 & ~a11184;
assign a11310 = a11184 & ~l934;
assign a11312 = ~a11310 & ~a11308;
assign a11314 = ~a11312 & a11170;
assign a11316 = ~a11314 & ~a11292;
assign a11318 = a11316 & ~l972;
assign a11320 = ~a11316 & l972;
assign a11322 = ~a11320 & ~a11318;
assign a11324 = a11190 & l1314;
assign a11326 = a11324 & ~a11188;
assign a11328 = a11188 & l1300;
assign a11330 = ~a11328 & ~a11326;
assign a11332 = ~a11330 & ~a11186;
assign a11334 = a11186 & l1286;
assign a11336 = ~a11334 & ~a11332;
assign a11338 = ~a11336 & ~a11184;
assign a11340 = a11184 & l1272;
assign a11342 = ~a11340 & ~a11338;
assign a11344 = ~a11342 & a11182;
assign a11346 = a11344 & ~a11180;
assign a11348 = a11190 & l1230;
assign a11350 = a11348 & ~a11188;
assign a11352 = a11188 & l1216;
assign a11354 = ~a11352 & ~a11350;
assign a11356 = ~a11354 & ~a11186;
assign a11358 = a11186 & l1202;
assign a11360 = ~a11358 & ~a11356;
assign a11362 = ~a11360 & ~a11184;
assign a11364 = a11184 & l1188;
assign a11366 = ~a11364 & ~a11362;
assign a11368 = ~a11366 & a11180;
assign a11370 = ~a11368 & ~a11346;
assign a11372 = ~a11370 & ~a11178;
assign a11374 = a11190 & l1146;
assign a11376 = a11374 & ~a11188;
assign a11378 = a11188 & l1132;
assign a11380 = ~a11378 & ~a11376;
assign a11382 = ~a11380 & ~a11186;
assign a11384 = a11186 & l1118;
assign a11386 = ~a11384 & ~a11382;
assign a11388 = ~a11386 & ~a11184;
assign a11390 = a11184 & l1104;
assign a11392 = ~a11390 & ~a11388;
assign a11394 = ~a11392 & a11178;
assign a11396 = ~a11394 & ~a11372;
assign a11398 = ~a11396 & ~a11174;
assign a11400 = a11190 & l1062;
assign a11402 = a11400 & ~a11188;
assign a11404 = a11188 & l1048;
assign a11406 = ~a11404 & ~a11402;
assign a11408 = ~a11406 & ~a11186;
assign a11410 = a11186 & l1034;
assign a11412 = ~a11410 & ~a11408;
assign a11414 = ~a11412 & ~a11184;
assign a11416 = a11184 & l1020;
assign a11418 = ~a11416 & ~a11414;
assign a11420 = ~a11418 & a11174;
assign a11422 = ~a11420 & ~a11398;
assign a11424 = ~a11422 & ~a11170;
assign a11426 = a11190 & l978;
assign a11428 = a11426 & ~a11188;
assign a11430 = a11188 & l964;
assign a11432 = ~a11430 & ~a11428;
assign a11434 = ~a11432 & ~a11186;
assign a11436 = a11186 & l950;
assign a11438 = ~a11436 & ~a11434;
assign a11440 = ~a11438 & ~a11184;
assign a11442 = a11184 & l936;
assign a11444 = ~a11442 & ~a11440;
assign a11446 = ~a11444 & a11170;
assign a11448 = ~a11446 & ~a11424;
assign a11450 = a11448 & ~l974;
assign a11452 = ~a11448 & l974;
assign a11454 = ~a11452 & ~a11450;
assign a11456 = a11454 & a11322;
assign a11458 = ~a11456 & ~a11166;
assign a11460 = ~l774 & ~l772;
assign a11462 = a11460 & ~l770;
assign a11464 = l774 & ~l772;
assign a11466 = a11464 & ~l770;
assign a11468 = ~l774 & l772;
assign a11470 = a11468 & ~l770;
assign a11472 = l774 & l772;
assign a11474 = a11472 & ~l770;
assign a11476 = a11460 & l770;
assign a11478 = a11464 & l770;
assign a11480 = ~l778 & ~l776;
assign a11482 = l778 & ~l776;
assign a11484 = ~l778 & l776;
assign a11486 = l778 & l776;
assign a11488 = a11486 & ~l1312;
assign a11490 = a11488 & ~a11484;
assign a11492 = a11484 & ~l1298;
assign a11494 = ~a11492 & ~a11490;
assign a11496 = ~a11494 & ~a11482;
assign a11498 = a11482 & ~l1284;
assign a11500 = ~a11498 & ~a11496;
assign a11502 = ~a11500 & ~a11480;
assign a11504 = a11480 & ~l1270;
assign a11506 = ~a11504 & ~a11502;
assign a11508 = ~a11506 & a11478;
assign a11510 = a11508 & ~a11476;
assign a11512 = a11486 & ~l1228;
assign a11514 = a11512 & ~a11484;
assign a11516 = a11484 & ~l1214;
assign a11518 = ~a11516 & ~a11514;
assign a11520 = ~a11518 & ~a11482;
assign a11522 = a11482 & ~l1200;
assign a11524 = ~a11522 & ~a11520;
assign a11526 = ~a11524 & ~a11480;
assign a11528 = a11480 & ~l1186;
assign a11530 = ~a11528 & ~a11526;
assign a11532 = ~a11530 & a11476;
assign a11534 = ~a11532 & ~a11510;
assign a11536 = ~a11534 & ~a11474;
assign a11538 = a11486 & ~l1144;
assign a11540 = a11538 & ~a11484;
assign a11542 = a11484 & ~l1130;
assign a11544 = ~a11542 & ~a11540;
assign a11546 = ~a11544 & ~a11482;
assign a11548 = a11482 & ~l1116;
assign a11550 = ~a11548 & ~a11546;
assign a11552 = ~a11550 & ~a11480;
assign a11554 = a11480 & ~l1102;
assign a11556 = ~a11554 & ~a11552;
assign a11558 = ~a11556 & a11474;
assign a11560 = ~a11558 & ~a11536;
assign a11562 = ~a11560 & ~a11470;
assign a11564 = a11486 & ~l1060;
assign a11566 = a11564 & ~a11484;
assign a11568 = a11484 & ~l1046;
assign a11570 = ~a11568 & ~a11566;
assign a11572 = ~a11570 & ~a11482;
assign a11574 = a11482 & ~l1032;
assign a11576 = ~a11574 & ~a11572;
assign a11578 = ~a11576 & ~a11480;
assign a11580 = a11480 & ~l1018;
assign a11582 = ~a11580 & ~a11578;
assign a11584 = ~a11582 & a11470;
assign a11586 = ~a11584 & ~a11562;
assign a11588 = ~a11586 & ~a11466;
assign a11590 = a11486 & ~l976;
assign a11592 = a11590 & ~a11484;
assign a11594 = a11484 & ~l962;
assign a11596 = ~a11594 & ~a11592;
assign a11598 = ~a11596 & ~a11482;
assign a11600 = a11482 & ~l948;
assign a11602 = ~a11600 & ~a11598;
assign a11604 = ~a11602 & ~a11480;
assign a11606 = a11480 & ~l934;
assign a11608 = ~a11606 & ~a11604;
assign a11610 = ~a11608 & a11466;
assign a11612 = ~a11610 & ~a11588;
assign a11614 = a11612 & ~l1014;
assign a11616 = ~a11612 & l1014;
assign a11618 = ~a11616 & ~a11614;
assign a11620 = a11486 & l1314;
assign a11622 = a11620 & ~a11484;
assign a11624 = a11484 & l1300;
assign a11626 = ~a11624 & ~a11622;
assign a11628 = ~a11626 & ~a11482;
assign a11630 = a11482 & l1286;
assign a11632 = ~a11630 & ~a11628;
assign a11634 = ~a11632 & ~a11480;
assign a11636 = a11480 & l1272;
assign a11638 = ~a11636 & ~a11634;
assign a11640 = ~a11638 & a11478;
assign a11642 = a11640 & ~a11476;
assign a11644 = a11486 & l1230;
assign a11646 = a11644 & ~a11484;
assign a11648 = a11484 & l1216;
assign a11650 = ~a11648 & ~a11646;
assign a11652 = ~a11650 & ~a11482;
assign a11654 = a11482 & l1202;
assign a11656 = ~a11654 & ~a11652;
assign a11658 = ~a11656 & ~a11480;
assign a11660 = a11480 & l1188;
assign a11662 = ~a11660 & ~a11658;
assign a11664 = ~a11662 & a11476;
assign a11666 = ~a11664 & ~a11642;
assign a11668 = ~a11666 & ~a11474;
assign a11670 = a11486 & l1146;
assign a11672 = a11670 & ~a11484;
assign a11674 = a11484 & l1132;
assign a11676 = ~a11674 & ~a11672;
assign a11678 = ~a11676 & ~a11482;
assign a11680 = a11482 & l1118;
assign a11682 = ~a11680 & ~a11678;
assign a11684 = ~a11682 & ~a11480;
assign a11686 = a11480 & l1104;
assign a11688 = ~a11686 & ~a11684;
assign a11690 = ~a11688 & a11474;
assign a11692 = ~a11690 & ~a11668;
assign a11694 = ~a11692 & ~a11470;
assign a11696 = a11486 & l1062;
assign a11698 = a11696 & ~a11484;
assign a11700 = a11484 & l1048;
assign a11702 = ~a11700 & ~a11698;
assign a11704 = ~a11702 & ~a11482;
assign a11706 = a11482 & l1034;
assign a11708 = ~a11706 & ~a11704;
assign a11710 = ~a11708 & ~a11480;
assign a11712 = a11480 & l1020;
assign a11714 = ~a11712 & ~a11710;
assign a11716 = ~a11714 & a11470;
assign a11718 = ~a11716 & ~a11694;
assign a11720 = ~a11718 & ~a11466;
assign a11722 = a11486 & l978;
assign a11724 = a11722 & ~a11484;
assign a11726 = a11484 & l964;
assign a11728 = ~a11726 & ~a11724;
assign a11730 = ~a11728 & ~a11482;
assign a11732 = a11482 & l950;
assign a11734 = ~a11732 & ~a11730;
assign a11736 = ~a11734 & ~a11480;
assign a11738 = a11480 & l936;
assign a11740 = ~a11738 & ~a11736;
assign a11742 = ~a11740 & a11466;
assign a11744 = ~a11742 & ~a11720;
assign a11746 = a11744 & ~l1016;
assign a11748 = ~a11744 & l1016;
assign a11750 = ~a11748 & ~a11746;
assign a11752 = a11750 & a11618;
assign a11754 = ~a11752 & ~a11462;
assign a11756 = ~l784 & ~l782;
assign a11758 = a11756 & ~l780;
assign a11760 = l784 & ~l782;
assign a11762 = a11760 & ~l780;
assign a11764 = ~l784 & l782;
assign a11766 = a11764 & ~l780;
assign a11768 = l784 & l782;
assign a11770 = a11768 & ~l780;
assign a11772 = a11756 & l780;
assign a11774 = a11760 & l780;
assign a11776 = ~l788 & ~l786;
assign a11778 = l788 & ~l786;
assign a11780 = ~l788 & l786;
assign a11782 = l788 & l786;
assign a11784 = a11782 & ~l1312;
assign a11786 = a11784 & ~a11780;
assign a11788 = a11780 & ~l1298;
assign a11790 = ~a11788 & ~a11786;
assign a11792 = ~a11790 & ~a11778;
assign a11794 = a11778 & ~l1284;
assign a11796 = ~a11794 & ~a11792;
assign a11798 = ~a11796 & ~a11776;
assign a11800 = a11776 & ~l1270;
assign a11802 = ~a11800 & ~a11798;
assign a11804 = ~a11802 & a11774;
assign a11806 = a11804 & ~a11772;
assign a11808 = a11782 & ~l1228;
assign a11810 = a11808 & ~a11780;
assign a11812 = a11780 & ~l1214;
assign a11814 = ~a11812 & ~a11810;
assign a11816 = ~a11814 & ~a11778;
assign a11818 = a11778 & ~l1200;
assign a11820 = ~a11818 & ~a11816;
assign a11822 = ~a11820 & ~a11776;
assign a11824 = a11776 & ~l1186;
assign a11826 = ~a11824 & ~a11822;
assign a11828 = ~a11826 & a11772;
assign a11830 = ~a11828 & ~a11806;
assign a11832 = ~a11830 & ~a11770;
assign a11834 = a11782 & ~l1144;
assign a11836 = a11834 & ~a11780;
assign a11838 = a11780 & ~l1130;
assign a11840 = ~a11838 & ~a11836;
assign a11842 = ~a11840 & ~a11778;
assign a11844 = a11778 & ~l1116;
assign a11846 = ~a11844 & ~a11842;
assign a11848 = ~a11846 & ~a11776;
assign a11850 = a11776 & ~l1102;
assign a11852 = ~a11850 & ~a11848;
assign a11854 = ~a11852 & a11770;
assign a11856 = ~a11854 & ~a11832;
assign a11858 = ~a11856 & ~a11766;
assign a11860 = a11782 & ~l1060;
assign a11862 = a11860 & ~a11780;
assign a11864 = a11780 & ~l1046;
assign a11866 = ~a11864 & ~a11862;
assign a11868 = ~a11866 & ~a11778;
assign a11870 = a11778 & ~l1032;
assign a11872 = ~a11870 & ~a11868;
assign a11874 = ~a11872 & ~a11776;
assign a11876 = a11776 & ~l1018;
assign a11878 = ~a11876 & ~a11874;
assign a11880 = ~a11878 & a11766;
assign a11882 = ~a11880 & ~a11858;
assign a11884 = ~a11882 & ~a11762;
assign a11886 = a11782 & ~l976;
assign a11888 = a11886 & ~a11780;
assign a11890 = a11780 & ~l962;
assign a11892 = ~a11890 & ~a11888;
assign a11894 = ~a11892 & ~a11778;
assign a11896 = a11778 & ~l948;
assign a11898 = ~a11896 & ~a11894;
assign a11900 = ~a11898 & ~a11776;
assign a11902 = a11776 & ~l934;
assign a11904 = ~a11902 & ~a11900;
assign a11906 = ~a11904 & a11762;
assign a11908 = ~a11906 & ~a11884;
assign a11910 = a11908 & ~l1028;
assign a11912 = ~a11908 & l1028;
assign a11914 = ~a11912 & ~a11910;
assign a11916 = a11782 & l1314;
assign a11918 = a11916 & ~a11780;
assign a11920 = a11780 & l1300;
assign a11922 = ~a11920 & ~a11918;
assign a11924 = ~a11922 & ~a11778;
assign a11926 = a11778 & l1286;
assign a11928 = ~a11926 & ~a11924;
assign a11930 = ~a11928 & ~a11776;
assign a11932 = a11776 & l1272;
assign a11934 = ~a11932 & ~a11930;
assign a11936 = ~a11934 & a11774;
assign a11938 = a11936 & ~a11772;
assign a11940 = a11782 & l1230;
assign a11942 = a11940 & ~a11780;
assign a11944 = a11780 & l1216;
assign a11946 = ~a11944 & ~a11942;
assign a11948 = ~a11946 & ~a11778;
assign a11950 = a11778 & l1202;
assign a11952 = ~a11950 & ~a11948;
assign a11954 = ~a11952 & ~a11776;
assign a11956 = a11776 & l1188;
assign a11958 = ~a11956 & ~a11954;
assign a11960 = ~a11958 & a11772;
assign a11962 = ~a11960 & ~a11938;
assign a11964 = ~a11962 & ~a11770;
assign a11966 = a11782 & l1146;
assign a11968 = a11966 & ~a11780;
assign a11970 = a11780 & l1132;
assign a11972 = ~a11970 & ~a11968;
assign a11974 = ~a11972 & ~a11778;
assign a11976 = a11778 & l1118;
assign a11978 = ~a11976 & ~a11974;
assign a11980 = ~a11978 & ~a11776;
assign a11982 = a11776 & l1104;
assign a11984 = ~a11982 & ~a11980;
assign a11986 = ~a11984 & a11770;
assign a11988 = ~a11986 & ~a11964;
assign a11990 = ~a11988 & ~a11766;
assign a11992 = a11782 & l1062;
assign a11994 = a11992 & ~a11780;
assign a11996 = a11780 & l1048;
assign a11998 = ~a11996 & ~a11994;
assign a12000 = ~a11998 & ~a11778;
assign a12002 = a11778 & l1034;
assign a12004 = ~a12002 & ~a12000;
assign a12006 = ~a12004 & ~a11776;
assign a12008 = a11776 & l1020;
assign a12010 = ~a12008 & ~a12006;
assign a12012 = ~a12010 & a11766;
assign a12014 = ~a12012 & ~a11990;
assign a12016 = ~a12014 & ~a11762;
assign a12018 = a11782 & l978;
assign a12020 = a12018 & ~a11780;
assign a12022 = a11780 & l964;
assign a12024 = ~a12022 & ~a12020;
assign a12026 = ~a12024 & ~a11778;
assign a12028 = a11778 & l950;
assign a12030 = ~a12028 & ~a12026;
assign a12032 = ~a12030 & ~a11776;
assign a12034 = a11776 & l936;
assign a12036 = ~a12034 & ~a12032;
assign a12038 = ~a12036 & a11762;
assign a12040 = ~a12038 & ~a12016;
assign a12042 = a12040 & ~l1030;
assign a12044 = ~a12040 & l1030;
assign a12046 = ~a12044 & ~a12042;
assign a12048 = a12046 & a11914;
assign a12050 = ~a12048 & ~a11758;
assign a12052 = ~l794 & ~l792;
assign a12054 = a12052 & ~l790;
assign a12056 = l794 & ~l792;
assign a12058 = a12056 & ~l790;
assign a12060 = ~l794 & l792;
assign a12062 = a12060 & ~l790;
assign a12064 = l794 & l792;
assign a12066 = a12064 & ~l790;
assign a12068 = a12052 & l790;
assign a12070 = a12056 & l790;
assign a12072 = ~l798 & ~l796;
assign a12074 = l798 & ~l796;
assign a12076 = ~l798 & l796;
assign a12078 = l798 & l796;
assign a12080 = a12078 & ~l1312;
assign a12082 = a12080 & ~a12076;
assign a12084 = a12076 & ~l1298;
assign a12086 = ~a12084 & ~a12082;
assign a12088 = ~a12086 & ~a12074;
assign a12090 = a12074 & ~l1284;
assign a12092 = ~a12090 & ~a12088;
assign a12094 = ~a12092 & ~a12072;
assign a12096 = a12072 & ~l1270;
assign a12098 = ~a12096 & ~a12094;
assign a12100 = ~a12098 & a12070;
assign a12102 = a12100 & ~a12068;
assign a12104 = a12078 & ~l1228;
assign a12106 = a12104 & ~a12076;
assign a12108 = a12076 & ~l1214;
assign a12110 = ~a12108 & ~a12106;
assign a12112 = ~a12110 & ~a12074;
assign a12114 = a12074 & ~l1200;
assign a12116 = ~a12114 & ~a12112;
assign a12118 = ~a12116 & ~a12072;
assign a12120 = a12072 & ~l1186;
assign a12122 = ~a12120 & ~a12118;
assign a12124 = ~a12122 & a12068;
assign a12126 = ~a12124 & ~a12102;
assign a12128 = ~a12126 & ~a12066;
assign a12130 = a12078 & ~l1144;
assign a12132 = a12130 & ~a12076;
assign a12134 = a12076 & ~l1130;
assign a12136 = ~a12134 & ~a12132;
assign a12138 = ~a12136 & ~a12074;
assign a12140 = a12074 & ~l1116;
assign a12142 = ~a12140 & ~a12138;
assign a12144 = ~a12142 & ~a12072;
assign a12146 = a12072 & ~l1102;
assign a12148 = ~a12146 & ~a12144;
assign a12150 = ~a12148 & a12066;
assign a12152 = ~a12150 & ~a12128;
assign a12154 = ~a12152 & ~a12062;
assign a12156 = a12078 & ~l1060;
assign a12158 = a12156 & ~a12076;
assign a12160 = a12076 & ~l1046;
assign a12162 = ~a12160 & ~a12158;
assign a12164 = ~a12162 & ~a12074;
assign a12166 = a12074 & ~l1032;
assign a12168 = ~a12166 & ~a12164;
assign a12170 = ~a12168 & ~a12072;
assign a12172 = a12072 & ~l1018;
assign a12174 = ~a12172 & ~a12170;
assign a12176 = ~a12174 & a12062;
assign a12178 = ~a12176 & ~a12154;
assign a12180 = ~a12178 & ~a12058;
assign a12182 = a12078 & ~l976;
assign a12184 = a12182 & ~a12076;
assign a12186 = a12076 & ~l962;
assign a12188 = ~a12186 & ~a12184;
assign a12190 = ~a12188 & ~a12074;
assign a12192 = a12074 & ~l948;
assign a12194 = ~a12192 & ~a12190;
assign a12196 = ~a12194 & ~a12072;
assign a12198 = a12072 & ~l934;
assign a12200 = ~a12198 & ~a12196;
assign a12202 = ~a12200 & a12058;
assign a12204 = ~a12202 & ~a12180;
assign a12206 = a12204 & ~l1042;
assign a12208 = ~a12204 & l1042;
assign a12210 = ~a12208 & ~a12206;
assign a12212 = a12078 & l1314;
assign a12214 = a12212 & ~a12076;
assign a12216 = a12076 & l1300;
assign a12218 = ~a12216 & ~a12214;
assign a12220 = ~a12218 & ~a12074;
assign a12222 = a12074 & l1286;
assign a12224 = ~a12222 & ~a12220;
assign a12226 = ~a12224 & ~a12072;
assign a12228 = a12072 & l1272;
assign a12230 = ~a12228 & ~a12226;
assign a12232 = ~a12230 & a12070;
assign a12234 = a12232 & ~a12068;
assign a12236 = a12078 & l1230;
assign a12238 = a12236 & ~a12076;
assign a12240 = a12076 & l1216;
assign a12242 = ~a12240 & ~a12238;
assign a12244 = ~a12242 & ~a12074;
assign a12246 = a12074 & l1202;
assign a12248 = ~a12246 & ~a12244;
assign a12250 = ~a12248 & ~a12072;
assign a12252 = a12072 & l1188;
assign a12254 = ~a12252 & ~a12250;
assign a12256 = ~a12254 & a12068;
assign a12258 = ~a12256 & ~a12234;
assign a12260 = ~a12258 & ~a12066;
assign a12262 = a12078 & l1146;
assign a12264 = a12262 & ~a12076;
assign a12266 = a12076 & l1132;
assign a12268 = ~a12266 & ~a12264;
assign a12270 = ~a12268 & ~a12074;
assign a12272 = a12074 & l1118;
assign a12274 = ~a12272 & ~a12270;
assign a12276 = ~a12274 & ~a12072;
assign a12278 = a12072 & l1104;
assign a12280 = ~a12278 & ~a12276;
assign a12282 = ~a12280 & a12066;
assign a12284 = ~a12282 & ~a12260;
assign a12286 = ~a12284 & ~a12062;
assign a12288 = a12078 & l1062;
assign a12290 = a12288 & ~a12076;
assign a12292 = a12076 & l1048;
assign a12294 = ~a12292 & ~a12290;
assign a12296 = ~a12294 & ~a12074;
assign a12298 = a12074 & l1034;
assign a12300 = ~a12298 & ~a12296;
assign a12302 = ~a12300 & ~a12072;
assign a12304 = a12072 & l1020;
assign a12306 = ~a12304 & ~a12302;
assign a12308 = ~a12306 & a12062;
assign a12310 = ~a12308 & ~a12286;
assign a12312 = ~a12310 & ~a12058;
assign a12314 = a12078 & l978;
assign a12316 = a12314 & ~a12076;
assign a12318 = a12076 & l964;
assign a12320 = ~a12318 & ~a12316;
assign a12322 = ~a12320 & ~a12074;
assign a12324 = a12074 & l950;
assign a12326 = ~a12324 & ~a12322;
assign a12328 = ~a12326 & ~a12072;
assign a12330 = a12072 & l936;
assign a12332 = ~a12330 & ~a12328;
assign a12334 = ~a12332 & a12058;
assign a12336 = ~a12334 & ~a12312;
assign a12338 = a12336 & ~l1044;
assign a12340 = ~a12336 & l1044;
assign a12342 = ~a12340 & ~a12338;
assign a12344 = a12342 & a12210;
assign a12346 = ~a12344 & ~a12054;
assign a12348 = ~l804 & ~l802;
assign a12350 = a12348 & ~l800;
assign a12352 = l804 & ~l802;
assign a12354 = a12352 & ~l800;
assign a12356 = ~l804 & l802;
assign a12358 = a12356 & ~l800;
assign a12360 = l804 & l802;
assign a12362 = a12360 & ~l800;
assign a12364 = a12348 & l800;
assign a12366 = a12352 & l800;
assign a12368 = ~l808 & ~l806;
assign a12370 = l808 & ~l806;
assign a12372 = ~l808 & l806;
assign a12374 = l808 & l806;
assign a12376 = a12374 & ~l1312;
assign a12378 = a12376 & ~a12372;
assign a12380 = a12372 & ~l1298;
assign a12382 = ~a12380 & ~a12378;
assign a12384 = ~a12382 & ~a12370;
assign a12386 = a12370 & ~l1284;
assign a12388 = ~a12386 & ~a12384;
assign a12390 = ~a12388 & ~a12368;
assign a12392 = a12368 & ~l1270;
assign a12394 = ~a12392 & ~a12390;
assign a12396 = ~a12394 & a12366;
assign a12398 = a12396 & ~a12364;
assign a12400 = a12374 & ~l1228;
assign a12402 = a12400 & ~a12372;
assign a12404 = a12372 & ~l1214;
assign a12406 = ~a12404 & ~a12402;
assign a12408 = ~a12406 & ~a12370;
assign a12410 = a12370 & ~l1200;
assign a12412 = ~a12410 & ~a12408;
assign a12414 = ~a12412 & ~a12368;
assign a12416 = a12368 & ~l1186;
assign a12418 = ~a12416 & ~a12414;
assign a12420 = ~a12418 & a12364;
assign a12422 = ~a12420 & ~a12398;
assign a12424 = ~a12422 & ~a12362;
assign a12426 = a12374 & ~l1144;
assign a12428 = a12426 & ~a12372;
assign a12430 = a12372 & ~l1130;
assign a12432 = ~a12430 & ~a12428;
assign a12434 = ~a12432 & ~a12370;
assign a12436 = a12370 & ~l1116;
assign a12438 = ~a12436 & ~a12434;
assign a12440 = ~a12438 & ~a12368;
assign a12442 = a12368 & ~l1102;
assign a12444 = ~a12442 & ~a12440;
assign a12446 = ~a12444 & a12362;
assign a12448 = ~a12446 & ~a12424;
assign a12450 = ~a12448 & ~a12358;
assign a12452 = a12374 & ~l1060;
assign a12454 = a12452 & ~a12372;
assign a12456 = a12372 & ~l1046;
assign a12458 = ~a12456 & ~a12454;
assign a12460 = ~a12458 & ~a12370;
assign a12462 = a12370 & ~l1032;
assign a12464 = ~a12462 & ~a12460;
assign a12466 = ~a12464 & ~a12368;
assign a12468 = a12368 & ~l1018;
assign a12470 = ~a12468 & ~a12466;
assign a12472 = ~a12470 & a12358;
assign a12474 = ~a12472 & ~a12450;
assign a12476 = ~a12474 & ~a12354;
assign a12478 = a12374 & ~l976;
assign a12480 = a12478 & ~a12372;
assign a12482 = a12372 & ~l962;
assign a12484 = ~a12482 & ~a12480;
assign a12486 = ~a12484 & ~a12370;
assign a12488 = a12370 & ~l948;
assign a12490 = ~a12488 & ~a12486;
assign a12492 = ~a12490 & ~a12368;
assign a12494 = a12368 & ~l934;
assign a12496 = ~a12494 & ~a12492;
assign a12498 = ~a12496 & a12354;
assign a12500 = ~a12498 & ~a12476;
assign a12502 = a12500 & ~l1056;
assign a12504 = ~a12500 & l1056;
assign a12506 = ~a12504 & ~a12502;
assign a12508 = a12374 & l1314;
assign a12510 = a12508 & ~a12372;
assign a12512 = a12372 & l1300;
assign a12514 = ~a12512 & ~a12510;
assign a12516 = ~a12514 & ~a12370;
assign a12518 = a12370 & l1286;
assign a12520 = ~a12518 & ~a12516;
assign a12522 = ~a12520 & ~a12368;
assign a12524 = a12368 & l1272;
assign a12526 = ~a12524 & ~a12522;
assign a12528 = ~a12526 & a12366;
assign a12530 = a12528 & ~a12364;
assign a12532 = a12374 & l1230;
assign a12534 = a12532 & ~a12372;
assign a12536 = a12372 & l1216;
assign a12538 = ~a12536 & ~a12534;
assign a12540 = ~a12538 & ~a12370;
assign a12542 = a12370 & l1202;
assign a12544 = ~a12542 & ~a12540;
assign a12546 = ~a12544 & ~a12368;
assign a12548 = a12368 & l1188;
assign a12550 = ~a12548 & ~a12546;
assign a12552 = ~a12550 & a12364;
assign a12554 = ~a12552 & ~a12530;
assign a12556 = ~a12554 & ~a12362;
assign a12558 = a12374 & l1146;
assign a12560 = a12558 & ~a12372;
assign a12562 = a12372 & l1132;
assign a12564 = ~a12562 & ~a12560;
assign a12566 = ~a12564 & ~a12370;
assign a12568 = a12370 & l1118;
assign a12570 = ~a12568 & ~a12566;
assign a12572 = ~a12570 & ~a12368;
assign a12574 = a12368 & l1104;
assign a12576 = ~a12574 & ~a12572;
assign a12578 = ~a12576 & a12362;
assign a12580 = ~a12578 & ~a12556;
assign a12582 = ~a12580 & ~a12358;
assign a12584 = a12374 & l1062;
assign a12586 = a12584 & ~a12372;
assign a12588 = a12372 & l1048;
assign a12590 = ~a12588 & ~a12586;
assign a12592 = ~a12590 & ~a12370;
assign a12594 = a12370 & l1034;
assign a12596 = ~a12594 & ~a12592;
assign a12598 = ~a12596 & ~a12368;
assign a12600 = a12368 & l1020;
assign a12602 = ~a12600 & ~a12598;
assign a12604 = ~a12602 & a12358;
assign a12606 = ~a12604 & ~a12582;
assign a12608 = ~a12606 & ~a12354;
assign a12610 = a12374 & l978;
assign a12612 = a12610 & ~a12372;
assign a12614 = a12372 & l964;
assign a12616 = ~a12614 & ~a12612;
assign a12618 = ~a12616 & ~a12370;
assign a12620 = a12370 & l950;
assign a12622 = ~a12620 & ~a12618;
assign a12624 = ~a12622 & ~a12368;
assign a12626 = a12368 & l936;
assign a12628 = ~a12626 & ~a12624;
assign a12630 = ~a12628 & a12354;
assign a12632 = ~a12630 & ~a12608;
assign a12634 = a12632 & ~l1058;
assign a12636 = ~a12632 & l1058;
assign a12638 = ~a12636 & ~a12634;
assign a12640 = a12638 & a12506;
assign a12642 = ~a12640 & ~a12350;
assign a12644 = ~l814 & ~l812;
assign a12646 = a12644 & ~l810;
assign a12648 = l814 & ~l812;
assign a12650 = a12648 & ~l810;
assign a12652 = ~l814 & l812;
assign a12654 = a12652 & ~l810;
assign a12656 = l814 & l812;
assign a12658 = a12656 & ~l810;
assign a12660 = a12644 & l810;
assign a12662 = a12648 & l810;
assign a12664 = ~l818 & ~l816;
assign a12666 = l818 & ~l816;
assign a12668 = ~l818 & l816;
assign a12670 = l818 & l816;
assign a12672 = a12670 & ~l1312;
assign a12674 = a12672 & ~a12668;
assign a12676 = a12668 & ~l1298;
assign a12678 = ~a12676 & ~a12674;
assign a12680 = ~a12678 & ~a12666;
assign a12682 = a12666 & ~l1284;
assign a12684 = ~a12682 & ~a12680;
assign a12686 = ~a12684 & ~a12664;
assign a12688 = a12664 & ~l1270;
assign a12690 = ~a12688 & ~a12686;
assign a12692 = ~a12690 & a12662;
assign a12694 = a12692 & ~a12660;
assign a12696 = a12670 & ~l1228;
assign a12698 = a12696 & ~a12668;
assign a12700 = a12668 & ~l1214;
assign a12702 = ~a12700 & ~a12698;
assign a12704 = ~a12702 & ~a12666;
assign a12706 = a12666 & ~l1200;
assign a12708 = ~a12706 & ~a12704;
assign a12710 = ~a12708 & ~a12664;
assign a12712 = a12664 & ~l1186;
assign a12714 = ~a12712 & ~a12710;
assign a12716 = ~a12714 & a12660;
assign a12718 = ~a12716 & ~a12694;
assign a12720 = ~a12718 & ~a12658;
assign a12722 = a12670 & ~l1144;
assign a12724 = a12722 & ~a12668;
assign a12726 = a12668 & ~l1130;
assign a12728 = ~a12726 & ~a12724;
assign a12730 = ~a12728 & ~a12666;
assign a12732 = a12666 & ~l1116;
assign a12734 = ~a12732 & ~a12730;
assign a12736 = ~a12734 & ~a12664;
assign a12738 = a12664 & ~l1102;
assign a12740 = ~a12738 & ~a12736;
assign a12742 = ~a12740 & a12658;
assign a12744 = ~a12742 & ~a12720;
assign a12746 = ~a12744 & ~a12654;
assign a12748 = a12670 & ~l1060;
assign a12750 = a12748 & ~a12668;
assign a12752 = a12668 & ~l1046;
assign a12754 = ~a12752 & ~a12750;
assign a12756 = ~a12754 & ~a12666;
assign a12758 = a12666 & ~l1032;
assign a12760 = ~a12758 & ~a12756;
assign a12762 = ~a12760 & ~a12664;
assign a12764 = a12664 & ~l1018;
assign a12766 = ~a12764 & ~a12762;
assign a12768 = ~a12766 & a12654;
assign a12770 = ~a12768 & ~a12746;
assign a12772 = ~a12770 & ~a12650;
assign a12774 = a12670 & ~l976;
assign a12776 = a12774 & ~a12668;
assign a12778 = a12668 & ~l962;
assign a12780 = ~a12778 & ~a12776;
assign a12782 = ~a12780 & ~a12666;
assign a12784 = a12666 & ~l948;
assign a12786 = ~a12784 & ~a12782;
assign a12788 = ~a12786 & ~a12664;
assign a12790 = a12664 & ~l934;
assign a12792 = ~a12790 & ~a12788;
assign a12794 = ~a12792 & a12650;
assign a12796 = ~a12794 & ~a12772;
assign a12798 = a12796 & ~l1098;
assign a12800 = ~a12796 & l1098;
assign a12802 = ~a12800 & ~a12798;
assign a12804 = a12670 & l1314;
assign a12806 = a12804 & ~a12668;
assign a12808 = a12668 & l1300;
assign a12810 = ~a12808 & ~a12806;
assign a12812 = ~a12810 & ~a12666;
assign a12814 = a12666 & l1286;
assign a12816 = ~a12814 & ~a12812;
assign a12818 = ~a12816 & ~a12664;
assign a12820 = a12664 & l1272;
assign a12822 = ~a12820 & ~a12818;
assign a12824 = ~a12822 & a12662;
assign a12826 = a12824 & ~a12660;
assign a12828 = a12670 & l1230;
assign a12830 = a12828 & ~a12668;
assign a12832 = a12668 & l1216;
assign a12834 = ~a12832 & ~a12830;
assign a12836 = ~a12834 & ~a12666;
assign a12838 = a12666 & l1202;
assign a12840 = ~a12838 & ~a12836;
assign a12842 = ~a12840 & ~a12664;
assign a12844 = a12664 & l1188;
assign a12846 = ~a12844 & ~a12842;
assign a12848 = ~a12846 & a12660;
assign a12850 = ~a12848 & ~a12826;
assign a12852 = ~a12850 & ~a12658;
assign a12854 = a12670 & l1146;
assign a12856 = a12854 & ~a12668;
assign a12858 = a12668 & l1132;
assign a12860 = ~a12858 & ~a12856;
assign a12862 = ~a12860 & ~a12666;
assign a12864 = a12666 & l1118;
assign a12866 = ~a12864 & ~a12862;
assign a12868 = ~a12866 & ~a12664;
assign a12870 = a12664 & l1104;
assign a12872 = ~a12870 & ~a12868;
assign a12874 = ~a12872 & a12658;
assign a12876 = ~a12874 & ~a12852;
assign a12878 = ~a12876 & ~a12654;
assign a12880 = a12670 & l1062;
assign a12882 = a12880 & ~a12668;
assign a12884 = a12668 & l1048;
assign a12886 = ~a12884 & ~a12882;
assign a12888 = ~a12886 & ~a12666;
assign a12890 = a12666 & l1034;
assign a12892 = ~a12890 & ~a12888;
assign a12894 = ~a12892 & ~a12664;
assign a12896 = a12664 & l1020;
assign a12898 = ~a12896 & ~a12894;
assign a12900 = ~a12898 & a12654;
assign a12902 = ~a12900 & ~a12878;
assign a12904 = ~a12902 & ~a12650;
assign a12906 = a12670 & l978;
assign a12908 = a12906 & ~a12668;
assign a12910 = a12668 & l964;
assign a12912 = ~a12910 & ~a12908;
assign a12914 = ~a12912 & ~a12666;
assign a12916 = a12666 & l950;
assign a12918 = ~a12916 & ~a12914;
assign a12920 = ~a12918 & ~a12664;
assign a12922 = a12664 & l936;
assign a12924 = ~a12922 & ~a12920;
assign a12926 = ~a12924 & a12650;
assign a12928 = ~a12926 & ~a12904;
assign a12930 = a12928 & ~l1100;
assign a12932 = ~a12928 & l1100;
assign a12934 = ~a12932 & ~a12930;
assign a12936 = a12934 & a12802;
assign a12938 = ~a12936 & ~a12646;
assign a12940 = ~l824 & ~l822;
assign a12942 = a12940 & ~l820;
assign a12944 = l824 & ~l822;
assign a12946 = a12944 & ~l820;
assign a12948 = ~l824 & l822;
assign a12950 = a12948 & ~l820;
assign a12952 = l824 & l822;
assign a12954 = a12952 & ~l820;
assign a12956 = a12940 & l820;
assign a12958 = a12944 & l820;
assign a12960 = ~l828 & ~l826;
assign a12962 = l828 & ~l826;
assign a12964 = ~l828 & l826;
assign a12966 = l828 & l826;
assign a12968 = a12966 & ~l1312;
assign a12970 = a12968 & ~a12964;
assign a12972 = a12964 & ~l1298;
assign a12974 = ~a12972 & ~a12970;
assign a12976 = ~a12974 & ~a12962;
assign a12978 = a12962 & ~l1284;
assign a12980 = ~a12978 & ~a12976;
assign a12982 = ~a12980 & ~a12960;
assign a12984 = a12960 & ~l1270;
assign a12986 = ~a12984 & ~a12982;
assign a12988 = ~a12986 & a12958;
assign a12990 = a12988 & ~a12956;
assign a12992 = a12966 & ~l1228;
assign a12994 = a12992 & ~a12964;
assign a12996 = a12964 & ~l1214;
assign a12998 = ~a12996 & ~a12994;
assign a13000 = ~a12998 & ~a12962;
assign a13002 = a12962 & ~l1200;
assign a13004 = ~a13002 & ~a13000;
assign a13006 = ~a13004 & ~a12960;
assign a13008 = a12960 & ~l1186;
assign a13010 = ~a13008 & ~a13006;
assign a13012 = ~a13010 & a12956;
assign a13014 = ~a13012 & ~a12990;
assign a13016 = ~a13014 & ~a12954;
assign a13018 = a12966 & ~l1144;
assign a13020 = a13018 & ~a12964;
assign a13022 = a12964 & ~l1130;
assign a13024 = ~a13022 & ~a13020;
assign a13026 = ~a13024 & ~a12962;
assign a13028 = a12962 & ~l1116;
assign a13030 = ~a13028 & ~a13026;
assign a13032 = ~a13030 & ~a12960;
assign a13034 = a12960 & ~l1102;
assign a13036 = ~a13034 & ~a13032;
assign a13038 = ~a13036 & a12954;
assign a13040 = ~a13038 & ~a13016;
assign a13042 = ~a13040 & ~a12950;
assign a13044 = a12966 & ~l1060;
assign a13046 = a13044 & ~a12964;
assign a13048 = a12964 & ~l1046;
assign a13050 = ~a13048 & ~a13046;
assign a13052 = ~a13050 & ~a12962;
assign a13054 = a12962 & ~l1032;
assign a13056 = ~a13054 & ~a13052;
assign a13058 = ~a13056 & ~a12960;
assign a13060 = a12960 & ~l1018;
assign a13062 = ~a13060 & ~a13058;
assign a13064 = ~a13062 & a12950;
assign a13066 = ~a13064 & ~a13042;
assign a13068 = ~a13066 & ~a12946;
assign a13070 = a12966 & ~l976;
assign a13072 = a13070 & ~a12964;
assign a13074 = a12964 & ~l962;
assign a13076 = ~a13074 & ~a13072;
assign a13078 = ~a13076 & ~a12962;
assign a13080 = a12962 & ~l948;
assign a13082 = ~a13080 & ~a13078;
assign a13084 = ~a13082 & ~a12960;
assign a13086 = a12960 & ~l934;
assign a13088 = ~a13086 & ~a13084;
assign a13090 = ~a13088 & a12946;
assign a13092 = ~a13090 & ~a13068;
assign a13094 = a13092 & ~l1112;
assign a13096 = ~a13092 & l1112;
assign a13098 = ~a13096 & ~a13094;
assign a13100 = a12966 & l1314;
assign a13102 = a13100 & ~a12964;
assign a13104 = a12964 & l1300;
assign a13106 = ~a13104 & ~a13102;
assign a13108 = ~a13106 & ~a12962;
assign a13110 = a12962 & l1286;
assign a13112 = ~a13110 & ~a13108;
assign a13114 = ~a13112 & ~a12960;
assign a13116 = a12960 & l1272;
assign a13118 = ~a13116 & ~a13114;
assign a13120 = ~a13118 & a12958;
assign a13122 = a13120 & ~a12956;
assign a13124 = a12966 & l1230;
assign a13126 = a13124 & ~a12964;
assign a13128 = a12964 & l1216;
assign a13130 = ~a13128 & ~a13126;
assign a13132 = ~a13130 & ~a12962;
assign a13134 = a12962 & l1202;
assign a13136 = ~a13134 & ~a13132;
assign a13138 = ~a13136 & ~a12960;
assign a13140 = a12960 & l1188;
assign a13142 = ~a13140 & ~a13138;
assign a13144 = ~a13142 & a12956;
assign a13146 = ~a13144 & ~a13122;
assign a13148 = ~a13146 & ~a12954;
assign a13150 = a12966 & l1146;
assign a13152 = a13150 & ~a12964;
assign a13154 = a12964 & l1132;
assign a13156 = ~a13154 & ~a13152;
assign a13158 = ~a13156 & ~a12962;
assign a13160 = a12962 & l1118;
assign a13162 = ~a13160 & ~a13158;
assign a13164 = ~a13162 & ~a12960;
assign a13166 = a12960 & l1104;
assign a13168 = ~a13166 & ~a13164;
assign a13170 = ~a13168 & a12954;
assign a13172 = ~a13170 & ~a13148;
assign a13174 = ~a13172 & ~a12950;
assign a13176 = a12966 & l1062;
assign a13178 = a13176 & ~a12964;
assign a13180 = a12964 & l1048;
assign a13182 = ~a13180 & ~a13178;
assign a13184 = ~a13182 & ~a12962;
assign a13186 = a12962 & l1034;
assign a13188 = ~a13186 & ~a13184;
assign a13190 = ~a13188 & ~a12960;
assign a13192 = a12960 & l1020;
assign a13194 = ~a13192 & ~a13190;
assign a13196 = ~a13194 & a12950;
assign a13198 = ~a13196 & ~a13174;
assign a13200 = ~a13198 & ~a12946;
assign a13202 = a12966 & l978;
assign a13204 = a13202 & ~a12964;
assign a13206 = a12964 & l964;
assign a13208 = ~a13206 & ~a13204;
assign a13210 = ~a13208 & ~a12962;
assign a13212 = a12962 & l950;
assign a13214 = ~a13212 & ~a13210;
assign a13216 = ~a13214 & ~a12960;
assign a13218 = a12960 & l936;
assign a13220 = ~a13218 & ~a13216;
assign a13222 = ~a13220 & a12946;
assign a13224 = ~a13222 & ~a13200;
assign a13226 = a13224 & ~l1114;
assign a13228 = ~a13224 & l1114;
assign a13230 = ~a13228 & ~a13226;
assign a13232 = a13230 & a13098;
assign a13234 = ~a13232 & ~a12942;
assign a13236 = ~l834 & ~l832;
assign a13238 = a13236 & ~l830;
assign a13240 = l834 & ~l832;
assign a13242 = a13240 & ~l830;
assign a13244 = ~l834 & l832;
assign a13246 = a13244 & ~l830;
assign a13248 = l834 & l832;
assign a13250 = a13248 & ~l830;
assign a13252 = a13236 & l830;
assign a13254 = a13240 & l830;
assign a13256 = ~l838 & ~l836;
assign a13258 = l838 & ~l836;
assign a13260 = ~l838 & l836;
assign a13262 = l838 & l836;
assign a13264 = a13262 & ~l1312;
assign a13266 = a13264 & ~a13260;
assign a13268 = a13260 & ~l1298;
assign a13270 = ~a13268 & ~a13266;
assign a13272 = ~a13270 & ~a13258;
assign a13274 = a13258 & ~l1284;
assign a13276 = ~a13274 & ~a13272;
assign a13278 = ~a13276 & ~a13256;
assign a13280 = a13256 & ~l1270;
assign a13282 = ~a13280 & ~a13278;
assign a13284 = ~a13282 & a13254;
assign a13286 = a13284 & ~a13252;
assign a13288 = a13262 & ~l1228;
assign a13290 = a13288 & ~a13260;
assign a13292 = a13260 & ~l1214;
assign a13294 = ~a13292 & ~a13290;
assign a13296 = ~a13294 & ~a13258;
assign a13298 = a13258 & ~l1200;
assign a13300 = ~a13298 & ~a13296;
assign a13302 = ~a13300 & ~a13256;
assign a13304 = a13256 & ~l1186;
assign a13306 = ~a13304 & ~a13302;
assign a13308 = ~a13306 & a13252;
assign a13310 = ~a13308 & ~a13286;
assign a13312 = ~a13310 & ~a13250;
assign a13314 = a13262 & ~l1144;
assign a13316 = a13314 & ~a13260;
assign a13318 = a13260 & ~l1130;
assign a13320 = ~a13318 & ~a13316;
assign a13322 = ~a13320 & ~a13258;
assign a13324 = a13258 & ~l1116;
assign a13326 = ~a13324 & ~a13322;
assign a13328 = ~a13326 & ~a13256;
assign a13330 = a13256 & ~l1102;
assign a13332 = ~a13330 & ~a13328;
assign a13334 = ~a13332 & a13250;
assign a13336 = ~a13334 & ~a13312;
assign a13338 = ~a13336 & ~a13246;
assign a13340 = a13262 & ~l1060;
assign a13342 = a13340 & ~a13260;
assign a13344 = a13260 & ~l1046;
assign a13346 = ~a13344 & ~a13342;
assign a13348 = ~a13346 & ~a13258;
assign a13350 = a13258 & ~l1032;
assign a13352 = ~a13350 & ~a13348;
assign a13354 = ~a13352 & ~a13256;
assign a13356 = a13256 & ~l1018;
assign a13358 = ~a13356 & ~a13354;
assign a13360 = ~a13358 & a13246;
assign a13362 = ~a13360 & ~a13338;
assign a13364 = ~a13362 & ~a13242;
assign a13366 = a13262 & ~l976;
assign a13368 = a13366 & ~a13260;
assign a13370 = a13260 & ~l962;
assign a13372 = ~a13370 & ~a13368;
assign a13374 = ~a13372 & ~a13258;
assign a13376 = a13258 & ~l948;
assign a13378 = ~a13376 & ~a13374;
assign a13380 = ~a13378 & ~a13256;
assign a13382 = a13256 & ~l934;
assign a13384 = ~a13382 & ~a13380;
assign a13386 = ~a13384 & a13242;
assign a13388 = ~a13386 & ~a13364;
assign a13390 = a13388 & ~l1126;
assign a13392 = ~a13388 & l1126;
assign a13394 = ~a13392 & ~a13390;
assign a13396 = a13262 & l1314;
assign a13398 = a13396 & ~a13260;
assign a13400 = a13260 & l1300;
assign a13402 = ~a13400 & ~a13398;
assign a13404 = ~a13402 & ~a13258;
assign a13406 = a13258 & l1286;
assign a13408 = ~a13406 & ~a13404;
assign a13410 = ~a13408 & ~a13256;
assign a13412 = a13256 & l1272;
assign a13414 = ~a13412 & ~a13410;
assign a13416 = ~a13414 & a13254;
assign a13418 = a13416 & ~a13252;
assign a13420 = a13262 & l1230;
assign a13422 = a13420 & ~a13260;
assign a13424 = a13260 & l1216;
assign a13426 = ~a13424 & ~a13422;
assign a13428 = ~a13426 & ~a13258;
assign a13430 = a13258 & l1202;
assign a13432 = ~a13430 & ~a13428;
assign a13434 = ~a13432 & ~a13256;
assign a13436 = a13256 & l1188;
assign a13438 = ~a13436 & ~a13434;
assign a13440 = ~a13438 & a13252;
assign a13442 = ~a13440 & ~a13418;
assign a13444 = ~a13442 & ~a13250;
assign a13446 = a13262 & l1146;
assign a13448 = a13446 & ~a13260;
assign a13450 = a13260 & l1132;
assign a13452 = ~a13450 & ~a13448;
assign a13454 = ~a13452 & ~a13258;
assign a13456 = a13258 & l1118;
assign a13458 = ~a13456 & ~a13454;
assign a13460 = ~a13458 & ~a13256;
assign a13462 = a13256 & l1104;
assign a13464 = ~a13462 & ~a13460;
assign a13466 = ~a13464 & a13250;
assign a13468 = ~a13466 & ~a13444;
assign a13470 = ~a13468 & ~a13246;
assign a13472 = a13262 & l1062;
assign a13474 = a13472 & ~a13260;
assign a13476 = a13260 & l1048;
assign a13478 = ~a13476 & ~a13474;
assign a13480 = ~a13478 & ~a13258;
assign a13482 = a13258 & l1034;
assign a13484 = ~a13482 & ~a13480;
assign a13486 = ~a13484 & ~a13256;
assign a13488 = a13256 & l1020;
assign a13490 = ~a13488 & ~a13486;
assign a13492 = ~a13490 & a13246;
assign a13494 = ~a13492 & ~a13470;
assign a13496 = ~a13494 & ~a13242;
assign a13498 = a13262 & l978;
assign a13500 = a13498 & ~a13260;
assign a13502 = a13260 & l964;
assign a13504 = ~a13502 & ~a13500;
assign a13506 = ~a13504 & ~a13258;
assign a13508 = a13258 & l950;
assign a13510 = ~a13508 & ~a13506;
assign a13512 = ~a13510 & ~a13256;
assign a13514 = a13256 & l936;
assign a13516 = ~a13514 & ~a13512;
assign a13518 = ~a13516 & a13242;
assign a13520 = ~a13518 & ~a13496;
assign a13522 = a13520 & ~l1128;
assign a13524 = ~a13520 & l1128;
assign a13526 = ~a13524 & ~a13522;
assign a13528 = a13526 & a13394;
assign a13530 = ~a13528 & ~a13238;
assign a13532 = ~l844 & ~l842;
assign a13534 = a13532 & ~l840;
assign a13536 = l844 & ~l842;
assign a13538 = a13536 & ~l840;
assign a13540 = ~l844 & l842;
assign a13542 = a13540 & ~l840;
assign a13544 = l844 & l842;
assign a13546 = a13544 & ~l840;
assign a13548 = a13532 & l840;
assign a13550 = a13536 & l840;
assign a13552 = ~l848 & ~l846;
assign a13554 = l848 & ~l846;
assign a13556 = ~l848 & l846;
assign a13558 = l848 & l846;
assign a13560 = a13558 & ~l1312;
assign a13562 = a13560 & ~a13556;
assign a13564 = a13556 & ~l1298;
assign a13566 = ~a13564 & ~a13562;
assign a13568 = ~a13566 & ~a13554;
assign a13570 = a13554 & ~l1284;
assign a13572 = ~a13570 & ~a13568;
assign a13574 = ~a13572 & ~a13552;
assign a13576 = a13552 & ~l1270;
assign a13578 = ~a13576 & ~a13574;
assign a13580 = ~a13578 & a13550;
assign a13582 = a13580 & ~a13548;
assign a13584 = a13558 & ~l1228;
assign a13586 = a13584 & ~a13556;
assign a13588 = a13556 & ~l1214;
assign a13590 = ~a13588 & ~a13586;
assign a13592 = ~a13590 & ~a13554;
assign a13594 = a13554 & ~l1200;
assign a13596 = ~a13594 & ~a13592;
assign a13598 = ~a13596 & ~a13552;
assign a13600 = a13552 & ~l1186;
assign a13602 = ~a13600 & ~a13598;
assign a13604 = ~a13602 & a13548;
assign a13606 = ~a13604 & ~a13582;
assign a13608 = ~a13606 & ~a13546;
assign a13610 = a13558 & ~l1144;
assign a13612 = a13610 & ~a13556;
assign a13614 = a13556 & ~l1130;
assign a13616 = ~a13614 & ~a13612;
assign a13618 = ~a13616 & ~a13554;
assign a13620 = a13554 & ~l1116;
assign a13622 = ~a13620 & ~a13618;
assign a13624 = ~a13622 & ~a13552;
assign a13626 = a13552 & ~l1102;
assign a13628 = ~a13626 & ~a13624;
assign a13630 = ~a13628 & a13546;
assign a13632 = ~a13630 & ~a13608;
assign a13634 = ~a13632 & ~a13542;
assign a13636 = a13558 & ~l1060;
assign a13638 = a13636 & ~a13556;
assign a13640 = a13556 & ~l1046;
assign a13642 = ~a13640 & ~a13638;
assign a13644 = ~a13642 & ~a13554;
assign a13646 = a13554 & ~l1032;
assign a13648 = ~a13646 & ~a13644;
assign a13650 = ~a13648 & ~a13552;
assign a13652 = a13552 & ~l1018;
assign a13654 = ~a13652 & ~a13650;
assign a13656 = ~a13654 & a13542;
assign a13658 = ~a13656 & ~a13634;
assign a13660 = ~a13658 & ~a13538;
assign a13662 = a13558 & ~l976;
assign a13664 = a13662 & ~a13556;
assign a13666 = a13556 & ~l962;
assign a13668 = ~a13666 & ~a13664;
assign a13670 = ~a13668 & ~a13554;
assign a13672 = a13554 & ~l948;
assign a13674 = ~a13672 & ~a13670;
assign a13676 = ~a13674 & ~a13552;
assign a13678 = a13552 & ~l934;
assign a13680 = ~a13678 & ~a13676;
assign a13682 = ~a13680 & a13538;
assign a13684 = ~a13682 & ~a13660;
assign a13686 = a13684 & ~l1140;
assign a13688 = ~a13684 & l1140;
assign a13690 = ~a13688 & ~a13686;
assign a13692 = a13558 & l1314;
assign a13694 = a13692 & ~a13556;
assign a13696 = a13556 & l1300;
assign a13698 = ~a13696 & ~a13694;
assign a13700 = ~a13698 & ~a13554;
assign a13702 = a13554 & l1286;
assign a13704 = ~a13702 & ~a13700;
assign a13706 = ~a13704 & ~a13552;
assign a13708 = a13552 & l1272;
assign a13710 = ~a13708 & ~a13706;
assign a13712 = ~a13710 & a13550;
assign a13714 = a13712 & ~a13548;
assign a13716 = a13558 & l1230;
assign a13718 = a13716 & ~a13556;
assign a13720 = a13556 & l1216;
assign a13722 = ~a13720 & ~a13718;
assign a13724 = ~a13722 & ~a13554;
assign a13726 = a13554 & l1202;
assign a13728 = ~a13726 & ~a13724;
assign a13730 = ~a13728 & ~a13552;
assign a13732 = a13552 & l1188;
assign a13734 = ~a13732 & ~a13730;
assign a13736 = ~a13734 & a13548;
assign a13738 = ~a13736 & ~a13714;
assign a13740 = ~a13738 & ~a13546;
assign a13742 = a13558 & l1146;
assign a13744 = a13742 & ~a13556;
assign a13746 = a13556 & l1132;
assign a13748 = ~a13746 & ~a13744;
assign a13750 = ~a13748 & ~a13554;
assign a13752 = a13554 & l1118;
assign a13754 = ~a13752 & ~a13750;
assign a13756 = ~a13754 & ~a13552;
assign a13758 = a13552 & l1104;
assign a13760 = ~a13758 & ~a13756;
assign a13762 = ~a13760 & a13546;
assign a13764 = ~a13762 & ~a13740;
assign a13766 = ~a13764 & ~a13542;
assign a13768 = a13558 & l1062;
assign a13770 = a13768 & ~a13556;
assign a13772 = a13556 & l1048;
assign a13774 = ~a13772 & ~a13770;
assign a13776 = ~a13774 & ~a13554;
assign a13778 = a13554 & l1034;
assign a13780 = ~a13778 & ~a13776;
assign a13782 = ~a13780 & ~a13552;
assign a13784 = a13552 & l1020;
assign a13786 = ~a13784 & ~a13782;
assign a13788 = ~a13786 & a13542;
assign a13790 = ~a13788 & ~a13766;
assign a13792 = ~a13790 & ~a13538;
assign a13794 = a13558 & l978;
assign a13796 = a13794 & ~a13556;
assign a13798 = a13556 & l964;
assign a13800 = ~a13798 & ~a13796;
assign a13802 = ~a13800 & ~a13554;
assign a13804 = a13554 & l950;
assign a13806 = ~a13804 & ~a13802;
assign a13808 = ~a13806 & ~a13552;
assign a13810 = a13552 & l936;
assign a13812 = ~a13810 & ~a13808;
assign a13814 = ~a13812 & a13538;
assign a13816 = ~a13814 & ~a13792;
assign a13818 = a13816 & ~l1142;
assign a13820 = ~a13816 & l1142;
assign a13822 = ~a13820 & ~a13818;
assign a13824 = a13822 & a13690;
assign a13826 = ~a13824 & ~a13534;
assign a13828 = ~l854 & ~l852;
assign a13830 = a13828 & ~l850;
assign a13832 = l854 & ~l852;
assign a13834 = a13832 & ~l850;
assign a13836 = ~l854 & l852;
assign a13838 = a13836 & ~l850;
assign a13840 = l854 & l852;
assign a13842 = a13840 & ~l850;
assign a13844 = a13828 & l850;
assign a13846 = a13832 & l850;
assign a13848 = ~l858 & ~l856;
assign a13850 = l858 & ~l856;
assign a13852 = ~l858 & l856;
assign a13854 = l858 & l856;
assign a13856 = a13854 & ~l1312;
assign a13858 = a13856 & ~a13852;
assign a13860 = a13852 & ~l1298;
assign a13862 = ~a13860 & ~a13858;
assign a13864 = ~a13862 & ~a13850;
assign a13866 = a13850 & ~l1284;
assign a13868 = ~a13866 & ~a13864;
assign a13870 = ~a13868 & ~a13848;
assign a13872 = a13848 & ~l1270;
assign a13874 = ~a13872 & ~a13870;
assign a13876 = ~a13874 & a13846;
assign a13878 = a13876 & ~a13844;
assign a13880 = a13854 & ~l1228;
assign a13882 = a13880 & ~a13852;
assign a13884 = a13852 & ~l1214;
assign a13886 = ~a13884 & ~a13882;
assign a13888 = ~a13886 & ~a13850;
assign a13890 = a13850 & ~l1200;
assign a13892 = ~a13890 & ~a13888;
assign a13894 = ~a13892 & ~a13848;
assign a13896 = a13848 & ~l1186;
assign a13898 = ~a13896 & ~a13894;
assign a13900 = ~a13898 & a13844;
assign a13902 = ~a13900 & ~a13878;
assign a13904 = ~a13902 & ~a13842;
assign a13906 = a13854 & ~l1144;
assign a13908 = a13906 & ~a13852;
assign a13910 = a13852 & ~l1130;
assign a13912 = ~a13910 & ~a13908;
assign a13914 = ~a13912 & ~a13850;
assign a13916 = a13850 & ~l1116;
assign a13918 = ~a13916 & ~a13914;
assign a13920 = ~a13918 & ~a13848;
assign a13922 = a13848 & ~l1102;
assign a13924 = ~a13922 & ~a13920;
assign a13926 = ~a13924 & a13842;
assign a13928 = ~a13926 & ~a13904;
assign a13930 = ~a13928 & ~a13838;
assign a13932 = a13854 & ~l1060;
assign a13934 = a13932 & ~a13852;
assign a13936 = a13852 & ~l1046;
assign a13938 = ~a13936 & ~a13934;
assign a13940 = ~a13938 & ~a13850;
assign a13942 = a13850 & ~l1032;
assign a13944 = ~a13942 & ~a13940;
assign a13946 = ~a13944 & ~a13848;
assign a13948 = a13848 & ~l1018;
assign a13950 = ~a13948 & ~a13946;
assign a13952 = ~a13950 & a13838;
assign a13954 = ~a13952 & ~a13930;
assign a13956 = ~a13954 & ~a13834;
assign a13958 = a13854 & ~l976;
assign a13960 = a13958 & ~a13852;
assign a13962 = a13852 & ~l962;
assign a13964 = ~a13962 & ~a13960;
assign a13966 = ~a13964 & ~a13850;
assign a13968 = a13850 & ~l948;
assign a13970 = ~a13968 & ~a13966;
assign a13972 = ~a13970 & ~a13848;
assign a13974 = a13848 & ~l934;
assign a13976 = ~a13974 & ~a13972;
assign a13978 = ~a13976 & a13834;
assign a13980 = ~a13978 & ~a13956;
assign a13982 = a13980 & ~l1182;
assign a13984 = ~a13980 & l1182;
assign a13986 = ~a13984 & ~a13982;
assign a13988 = a13854 & l1314;
assign a13990 = a13988 & ~a13852;
assign a13992 = a13852 & l1300;
assign a13994 = ~a13992 & ~a13990;
assign a13996 = ~a13994 & ~a13850;
assign a13998 = a13850 & l1286;
assign a14000 = ~a13998 & ~a13996;
assign a14002 = ~a14000 & ~a13848;
assign a14004 = a13848 & l1272;
assign a14006 = ~a14004 & ~a14002;
assign a14008 = ~a14006 & a13846;
assign a14010 = a14008 & ~a13844;
assign a14012 = a13854 & l1230;
assign a14014 = a14012 & ~a13852;
assign a14016 = a13852 & l1216;
assign a14018 = ~a14016 & ~a14014;
assign a14020 = ~a14018 & ~a13850;
assign a14022 = a13850 & l1202;
assign a14024 = ~a14022 & ~a14020;
assign a14026 = ~a14024 & ~a13848;
assign a14028 = a13848 & l1188;
assign a14030 = ~a14028 & ~a14026;
assign a14032 = ~a14030 & a13844;
assign a14034 = ~a14032 & ~a14010;
assign a14036 = ~a14034 & ~a13842;
assign a14038 = a13854 & l1146;
assign a14040 = a14038 & ~a13852;
assign a14042 = a13852 & l1132;
assign a14044 = ~a14042 & ~a14040;
assign a14046 = ~a14044 & ~a13850;
assign a14048 = a13850 & l1118;
assign a14050 = ~a14048 & ~a14046;
assign a14052 = ~a14050 & ~a13848;
assign a14054 = a13848 & l1104;
assign a14056 = ~a14054 & ~a14052;
assign a14058 = ~a14056 & a13842;
assign a14060 = ~a14058 & ~a14036;
assign a14062 = ~a14060 & ~a13838;
assign a14064 = a13854 & l1062;
assign a14066 = a14064 & ~a13852;
assign a14068 = a13852 & l1048;
assign a14070 = ~a14068 & ~a14066;
assign a14072 = ~a14070 & ~a13850;
assign a14074 = a13850 & l1034;
assign a14076 = ~a14074 & ~a14072;
assign a14078 = ~a14076 & ~a13848;
assign a14080 = a13848 & l1020;
assign a14082 = ~a14080 & ~a14078;
assign a14084 = ~a14082 & a13838;
assign a14086 = ~a14084 & ~a14062;
assign a14088 = ~a14086 & ~a13834;
assign a14090 = a13854 & l978;
assign a14092 = a14090 & ~a13852;
assign a14094 = a13852 & l964;
assign a14096 = ~a14094 & ~a14092;
assign a14098 = ~a14096 & ~a13850;
assign a14100 = a13850 & l950;
assign a14102 = ~a14100 & ~a14098;
assign a14104 = ~a14102 & ~a13848;
assign a14106 = a13848 & l936;
assign a14108 = ~a14106 & ~a14104;
assign a14110 = ~a14108 & a13834;
assign a14112 = ~a14110 & ~a14088;
assign a14114 = a14112 & ~l1184;
assign a14116 = ~a14112 & l1184;
assign a14118 = ~a14116 & ~a14114;
assign a14120 = a14118 & a13986;
assign a14122 = ~a14120 & ~a13830;
assign a14124 = ~l864 & ~l862;
assign a14126 = a14124 & ~l860;
assign a14128 = l864 & ~l862;
assign a14130 = a14128 & ~l860;
assign a14132 = ~l864 & l862;
assign a14134 = a14132 & ~l860;
assign a14136 = l864 & l862;
assign a14138 = a14136 & ~l860;
assign a14140 = a14124 & l860;
assign a14142 = a14128 & l860;
assign a14144 = ~l868 & ~l866;
assign a14146 = l868 & ~l866;
assign a14148 = ~l868 & l866;
assign a14150 = l868 & l866;
assign a14152 = a14150 & ~l1312;
assign a14154 = a14152 & ~a14148;
assign a14156 = a14148 & ~l1298;
assign a14158 = ~a14156 & ~a14154;
assign a14160 = ~a14158 & ~a14146;
assign a14162 = a14146 & ~l1284;
assign a14164 = ~a14162 & ~a14160;
assign a14166 = ~a14164 & ~a14144;
assign a14168 = a14144 & ~l1270;
assign a14170 = ~a14168 & ~a14166;
assign a14172 = ~a14170 & a14142;
assign a14174 = a14172 & ~a14140;
assign a14176 = a14150 & ~l1228;
assign a14178 = a14176 & ~a14148;
assign a14180 = a14148 & ~l1214;
assign a14182 = ~a14180 & ~a14178;
assign a14184 = ~a14182 & ~a14146;
assign a14186 = a14146 & ~l1200;
assign a14188 = ~a14186 & ~a14184;
assign a14190 = ~a14188 & ~a14144;
assign a14192 = a14144 & ~l1186;
assign a14194 = ~a14192 & ~a14190;
assign a14196 = ~a14194 & a14140;
assign a14198 = ~a14196 & ~a14174;
assign a14200 = ~a14198 & ~a14138;
assign a14202 = a14150 & ~l1144;
assign a14204 = a14202 & ~a14148;
assign a14206 = a14148 & ~l1130;
assign a14208 = ~a14206 & ~a14204;
assign a14210 = ~a14208 & ~a14146;
assign a14212 = a14146 & ~l1116;
assign a14214 = ~a14212 & ~a14210;
assign a14216 = ~a14214 & ~a14144;
assign a14218 = a14144 & ~l1102;
assign a14220 = ~a14218 & ~a14216;
assign a14222 = ~a14220 & a14138;
assign a14224 = ~a14222 & ~a14200;
assign a14226 = ~a14224 & ~a14134;
assign a14228 = a14150 & ~l1060;
assign a14230 = a14228 & ~a14148;
assign a14232 = a14148 & ~l1046;
assign a14234 = ~a14232 & ~a14230;
assign a14236 = ~a14234 & ~a14146;
assign a14238 = a14146 & ~l1032;
assign a14240 = ~a14238 & ~a14236;
assign a14242 = ~a14240 & ~a14144;
assign a14244 = a14144 & ~l1018;
assign a14246 = ~a14244 & ~a14242;
assign a14248 = ~a14246 & a14134;
assign a14250 = ~a14248 & ~a14226;
assign a14252 = ~a14250 & ~a14130;
assign a14254 = a14150 & ~l976;
assign a14256 = a14254 & ~a14148;
assign a14258 = a14148 & ~l962;
assign a14260 = ~a14258 & ~a14256;
assign a14262 = ~a14260 & ~a14146;
assign a14264 = a14146 & ~l948;
assign a14266 = ~a14264 & ~a14262;
assign a14268 = ~a14266 & ~a14144;
assign a14270 = a14144 & ~l934;
assign a14272 = ~a14270 & ~a14268;
assign a14274 = ~a14272 & a14130;
assign a14276 = ~a14274 & ~a14252;
assign a14278 = a14276 & ~l1196;
assign a14280 = ~a14276 & l1196;
assign a14282 = ~a14280 & ~a14278;
assign a14284 = a14150 & l1314;
assign a14286 = a14284 & ~a14148;
assign a14288 = a14148 & l1300;
assign a14290 = ~a14288 & ~a14286;
assign a14292 = ~a14290 & ~a14146;
assign a14294 = a14146 & l1286;
assign a14296 = ~a14294 & ~a14292;
assign a14298 = ~a14296 & ~a14144;
assign a14300 = a14144 & l1272;
assign a14302 = ~a14300 & ~a14298;
assign a14304 = ~a14302 & a14142;
assign a14306 = a14304 & ~a14140;
assign a14308 = a14150 & l1230;
assign a14310 = a14308 & ~a14148;
assign a14312 = a14148 & l1216;
assign a14314 = ~a14312 & ~a14310;
assign a14316 = ~a14314 & ~a14146;
assign a14318 = a14146 & l1202;
assign a14320 = ~a14318 & ~a14316;
assign a14322 = ~a14320 & ~a14144;
assign a14324 = a14144 & l1188;
assign a14326 = ~a14324 & ~a14322;
assign a14328 = ~a14326 & a14140;
assign a14330 = ~a14328 & ~a14306;
assign a14332 = ~a14330 & ~a14138;
assign a14334 = a14150 & l1146;
assign a14336 = a14334 & ~a14148;
assign a14338 = a14148 & l1132;
assign a14340 = ~a14338 & ~a14336;
assign a14342 = ~a14340 & ~a14146;
assign a14344 = a14146 & l1118;
assign a14346 = ~a14344 & ~a14342;
assign a14348 = ~a14346 & ~a14144;
assign a14350 = a14144 & l1104;
assign a14352 = ~a14350 & ~a14348;
assign a14354 = ~a14352 & a14138;
assign a14356 = ~a14354 & ~a14332;
assign a14358 = ~a14356 & ~a14134;
assign a14360 = a14150 & l1062;
assign a14362 = a14360 & ~a14148;
assign a14364 = a14148 & l1048;
assign a14366 = ~a14364 & ~a14362;
assign a14368 = ~a14366 & ~a14146;
assign a14370 = a14146 & l1034;
assign a14372 = ~a14370 & ~a14368;
assign a14374 = ~a14372 & ~a14144;
assign a14376 = a14144 & l1020;
assign a14378 = ~a14376 & ~a14374;
assign a14380 = ~a14378 & a14134;
assign a14382 = ~a14380 & ~a14358;
assign a14384 = ~a14382 & ~a14130;
assign a14386 = a14150 & l978;
assign a14388 = a14386 & ~a14148;
assign a14390 = a14148 & l964;
assign a14392 = ~a14390 & ~a14388;
assign a14394 = ~a14392 & ~a14146;
assign a14396 = a14146 & l950;
assign a14398 = ~a14396 & ~a14394;
assign a14400 = ~a14398 & ~a14144;
assign a14402 = a14144 & l936;
assign a14404 = ~a14402 & ~a14400;
assign a14406 = ~a14404 & a14130;
assign a14408 = ~a14406 & ~a14384;
assign a14410 = a14408 & ~l1198;
assign a14412 = ~a14408 & l1198;
assign a14414 = ~a14412 & ~a14410;
assign a14416 = a14414 & a14282;
assign a14418 = ~a14416 & ~a14126;
assign a14420 = ~l874 & ~l872;
assign a14422 = a14420 & ~l870;
assign a14424 = l874 & ~l872;
assign a14426 = a14424 & ~l870;
assign a14428 = ~l874 & l872;
assign a14430 = a14428 & ~l870;
assign a14432 = l874 & l872;
assign a14434 = a14432 & ~l870;
assign a14436 = a14420 & l870;
assign a14438 = a14424 & l870;
assign a14440 = ~l878 & ~l876;
assign a14442 = l878 & ~l876;
assign a14444 = ~l878 & l876;
assign a14446 = l878 & l876;
assign a14448 = a14446 & ~l1312;
assign a14450 = a14448 & ~a14444;
assign a14452 = a14444 & ~l1298;
assign a14454 = ~a14452 & ~a14450;
assign a14456 = ~a14454 & ~a14442;
assign a14458 = a14442 & ~l1284;
assign a14460 = ~a14458 & ~a14456;
assign a14462 = ~a14460 & ~a14440;
assign a14464 = a14440 & ~l1270;
assign a14466 = ~a14464 & ~a14462;
assign a14468 = ~a14466 & a14438;
assign a14470 = a14468 & ~a14436;
assign a14472 = a14446 & ~l1228;
assign a14474 = a14472 & ~a14444;
assign a14476 = a14444 & ~l1214;
assign a14478 = ~a14476 & ~a14474;
assign a14480 = ~a14478 & ~a14442;
assign a14482 = a14442 & ~l1200;
assign a14484 = ~a14482 & ~a14480;
assign a14486 = ~a14484 & ~a14440;
assign a14488 = a14440 & ~l1186;
assign a14490 = ~a14488 & ~a14486;
assign a14492 = ~a14490 & a14436;
assign a14494 = ~a14492 & ~a14470;
assign a14496 = ~a14494 & ~a14434;
assign a14498 = a14446 & ~l1144;
assign a14500 = a14498 & ~a14444;
assign a14502 = a14444 & ~l1130;
assign a14504 = ~a14502 & ~a14500;
assign a14506 = ~a14504 & ~a14442;
assign a14508 = a14442 & ~l1116;
assign a14510 = ~a14508 & ~a14506;
assign a14512 = ~a14510 & ~a14440;
assign a14514 = a14440 & ~l1102;
assign a14516 = ~a14514 & ~a14512;
assign a14518 = ~a14516 & a14434;
assign a14520 = ~a14518 & ~a14496;
assign a14522 = ~a14520 & ~a14430;
assign a14524 = a14446 & ~l1060;
assign a14526 = a14524 & ~a14444;
assign a14528 = a14444 & ~l1046;
assign a14530 = ~a14528 & ~a14526;
assign a14532 = ~a14530 & ~a14442;
assign a14534 = a14442 & ~l1032;
assign a14536 = ~a14534 & ~a14532;
assign a14538 = ~a14536 & ~a14440;
assign a14540 = a14440 & ~l1018;
assign a14542 = ~a14540 & ~a14538;
assign a14544 = ~a14542 & a14430;
assign a14546 = ~a14544 & ~a14522;
assign a14548 = ~a14546 & ~a14426;
assign a14550 = a14446 & ~l976;
assign a14552 = a14550 & ~a14444;
assign a14554 = a14444 & ~l962;
assign a14556 = ~a14554 & ~a14552;
assign a14558 = ~a14556 & ~a14442;
assign a14560 = a14442 & ~l948;
assign a14562 = ~a14560 & ~a14558;
assign a14564 = ~a14562 & ~a14440;
assign a14566 = a14440 & ~l934;
assign a14568 = ~a14566 & ~a14564;
assign a14570 = ~a14568 & a14426;
assign a14572 = ~a14570 & ~a14548;
assign a14574 = a14572 & ~l1210;
assign a14576 = ~a14572 & l1210;
assign a14578 = ~a14576 & ~a14574;
assign a14580 = a14446 & l1314;
assign a14582 = a14580 & ~a14444;
assign a14584 = a14444 & l1300;
assign a14586 = ~a14584 & ~a14582;
assign a14588 = ~a14586 & ~a14442;
assign a14590 = a14442 & l1286;
assign a14592 = ~a14590 & ~a14588;
assign a14594 = ~a14592 & ~a14440;
assign a14596 = a14440 & l1272;
assign a14598 = ~a14596 & ~a14594;
assign a14600 = ~a14598 & a14438;
assign a14602 = a14600 & ~a14436;
assign a14604 = a14446 & l1230;
assign a14606 = a14604 & ~a14444;
assign a14608 = a14444 & l1216;
assign a14610 = ~a14608 & ~a14606;
assign a14612 = ~a14610 & ~a14442;
assign a14614 = a14442 & l1202;
assign a14616 = ~a14614 & ~a14612;
assign a14618 = ~a14616 & ~a14440;
assign a14620 = a14440 & l1188;
assign a14622 = ~a14620 & ~a14618;
assign a14624 = ~a14622 & a14436;
assign a14626 = ~a14624 & ~a14602;
assign a14628 = ~a14626 & ~a14434;
assign a14630 = a14446 & l1146;
assign a14632 = a14630 & ~a14444;
assign a14634 = a14444 & l1132;
assign a14636 = ~a14634 & ~a14632;
assign a14638 = ~a14636 & ~a14442;
assign a14640 = a14442 & l1118;
assign a14642 = ~a14640 & ~a14638;
assign a14644 = ~a14642 & ~a14440;
assign a14646 = a14440 & l1104;
assign a14648 = ~a14646 & ~a14644;
assign a14650 = ~a14648 & a14434;
assign a14652 = ~a14650 & ~a14628;
assign a14654 = ~a14652 & ~a14430;
assign a14656 = a14446 & l1062;
assign a14658 = a14656 & ~a14444;
assign a14660 = a14444 & l1048;
assign a14662 = ~a14660 & ~a14658;
assign a14664 = ~a14662 & ~a14442;
assign a14666 = a14442 & l1034;
assign a14668 = ~a14666 & ~a14664;
assign a14670 = ~a14668 & ~a14440;
assign a14672 = a14440 & l1020;
assign a14674 = ~a14672 & ~a14670;
assign a14676 = ~a14674 & a14430;
assign a14678 = ~a14676 & ~a14654;
assign a14680 = ~a14678 & ~a14426;
assign a14682 = a14446 & l978;
assign a14684 = a14682 & ~a14444;
assign a14686 = a14444 & l964;
assign a14688 = ~a14686 & ~a14684;
assign a14690 = ~a14688 & ~a14442;
assign a14692 = a14442 & l950;
assign a14694 = ~a14692 & ~a14690;
assign a14696 = ~a14694 & ~a14440;
assign a14698 = a14440 & l936;
assign a14700 = ~a14698 & ~a14696;
assign a14702 = ~a14700 & a14426;
assign a14704 = ~a14702 & ~a14680;
assign a14706 = a14704 & ~l1212;
assign a14708 = ~a14704 & l1212;
assign a14710 = ~a14708 & ~a14706;
assign a14712 = a14710 & a14578;
assign a14714 = ~a14712 & ~a14422;
assign a14716 = ~l884 & ~l882;
assign a14718 = a14716 & ~l880;
assign a14720 = l884 & ~l882;
assign a14722 = a14720 & ~l880;
assign a14724 = ~l884 & l882;
assign a14726 = a14724 & ~l880;
assign a14728 = l884 & l882;
assign a14730 = a14728 & ~l880;
assign a14732 = a14716 & l880;
assign a14734 = a14720 & l880;
assign a14736 = ~l888 & ~l886;
assign a14738 = l888 & ~l886;
assign a14740 = ~l888 & l886;
assign a14742 = l888 & l886;
assign a14744 = a14742 & ~l1312;
assign a14746 = a14744 & ~a14740;
assign a14748 = a14740 & ~l1298;
assign a14750 = ~a14748 & ~a14746;
assign a14752 = ~a14750 & ~a14738;
assign a14754 = a14738 & ~l1284;
assign a14756 = ~a14754 & ~a14752;
assign a14758 = ~a14756 & ~a14736;
assign a14760 = a14736 & ~l1270;
assign a14762 = ~a14760 & ~a14758;
assign a14764 = ~a14762 & a14734;
assign a14766 = a14764 & ~a14732;
assign a14768 = a14742 & ~l1228;
assign a14770 = a14768 & ~a14740;
assign a14772 = a14740 & ~l1214;
assign a14774 = ~a14772 & ~a14770;
assign a14776 = ~a14774 & ~a14738;
assign a14778 = a14738 & ~l1200;
assign a14780 = ~a14778 & ~a14776;
assign a14782 = ~a14780 & ~a14736;
assign a14784 = a14736 & ~l1186;
assign a14786 = ~a14784 & ~a14782;
assign a14788 = ~a14786 & a14732;
assign a14790 = ~a14788 & ~a14766;
assign a14792 = ~a14790 & ~a14730;
assign a14794 = a14742 & ~l1144;
assign a14796 = a14794 & ~a14740;
assign a14798 = a14740 & ~l1130;
assign a14800 = ~a14798 & ~a14796;
assign a14802 = ~a14800 & ~a14738;
assign a14804 = a14738 & ~l1116;
assign a14806 = ~a14804 & ~a14802;
assign a14808 = ~a14806 & ~a14736;
assign a14810 = a14736 & ~l1102;
assign a14812 = ~a14810 & ~a14808;
assign a14814 = ~a14812 & a14730;
assign a14816 = ~a14814 & ~a14792;
assign a14818 = ~a14816 & ~a14726;
assign a14820 = a14742 & ~l1060;
assign a14822 = a14820 & ~a14740;
assign a14824 = a14740 & ~l1046;
assign a14826 = ~a14824 & ~a14822;
assign a14828 = ~a14826 & ~a14738;
assign a14830 = a14738 & ~l1032;
assign a14832 = ~a14830 & ~a14828;
assign a14834 = ~a14832 & ~a14736;
assign a14836 = a14736 & ~l1018;
assign a14838 = ~a14836 & ~a14834;
assign a14840 = ~a14838 & a14726;
assign a14842 = ~a14840 & ~a14818;
assign a14844 = ~a14842 & ~a14722;
assign a14846 = a14742 & ~l976;
assign a14848 = a14846 & ~a14740;
assign a14850 = a14740 & ~l962;
assign a14852 = ~a14850 & ~a14848;
assign a14854 = ~a14852 & ~a14738;
assign a14856 = a14738 & ~l948;
assign a14858 = ~a14856 & ~a14854;
assign a14860 = ~a14858 & ~a14736;
assign a14862 = a14736 & ~l934;
assign a14864 = ~a14862 & ~a14860;
assign a14866 = ~a14864 & a14722;
assign a14868 = ~a14866 & ~a14844;
assign a14870 = a14868 & ~l1224;
assign a14872 = ~a14868 & l1224;
assign a14874 = ~a14872 & ~a14870;
assign a14876 = a14742 & l1314;
assign a14878 = a14876 & ~a14740;
assign a14880 = a14740 & l1300;
assign a14882 = ~a14880 & ~a14878;
assign a14884 = ~a14882 & ~a14738;
assign a14886 = a14738 & l1286;
assign a14888 = ~a14886 & ~a14884;
assign a14890 = ~a14888 & ~a14736;
assign a14892 = a14736 & l1272;
assign a14894 = ~a14892 & ~a14890;
assign a14896 = ~a14894 & a14734;
assign a14898 = a14896 & ~a14732;
assign a14900 = a14742 & l1230;
assign a14902 = a14900 & ~a14740;
assign a14904 = a14740 & l1216;
assign a14906 = ~a14904 & ~a14902;
assign a14908 = ~a14906 & ~a14738;
assign a14910 = a14738 & l1202;
assign a14912 = ~a14910 & ~a14908;
assign a14914 = ~a14912 & ~a14736;
assign a14916 = a14736 & l1188;
assign a14918 = ~a14916 & ~a14914;
assign a14920 = ~a14918 & a14732;
assign a14922 = ~a14920 & ~a14898;
assign a14924 = ~a14922 & ~a14730;
assign a14926 = a14742 & l1146;
assign a14928 = a14926 & ~a14740;
assign a14930 = a14740 & l1132;
assign a14932 = ~a14930 & ~a14928;
assign a14934 = ~a14932 & ~a14738;
assign a14936 = a14738 & l1118;
assign a14938 = ~a14936 & ~a14934;
assign a14940 = ~a14938 & ~a14736;
assign a14942 = a14736 & l1104;
assign a14944 = ~a14942 & ~a14940;
assign a14946 = ~a14944 & a14730;
assign a14948 = ~a14946 & ~a14924;
assign a14950 = ~a14948 & ~a14726;
assign a14952 = a14742 & l1062;
assign a14954 = a14952 & ~a14740;
assign a14956 = a14740 & l1048;
assign a14958 = ~a14956 & ~a14954;
assign a14960 = ~a14958 & ~a14738;
assign a14962 = a14738 & l1034;
assign a14964 = ~a14962 & ~a14960;
assign a14966 = ~a14964 & ~a14736;
assign a14968 = a14736 & l1020;
assign a14970 = ~a14968 & ~a14966;
assign a14972 = ~a14970 & a14726;
assign a14974 = ~a14972 & ~a14950;
assign a14976 = ~a14974 & ~a14722;
assign a14978 = a14742 & l978;
assign a14980 = a14978 & ~a14740;
assign a14982 = a14740 & l964;
assign a14984 = ~a14982 & ~a14980;
assign a14986 = ~a14984 & ~a14738;
assign a14988 = a14738 & l950;
assign a14990 = ~a14988 & ~a14986;
assign a14992 = ~a14990 & ~a14736;
assign a14994 = a14736 & l936;
assign a14996 = ~a14994 & ~a14992;
assign a14998 = ~a14996 & a14722;
assign a15000 = ~a14998 & ~a14976;
assign a15002 = a15000 & ~l1226;
assign a15004 = ~a15000 & l1226;
assign a15006 = ~a15004 & ~a15002;
assign a15008 = a15006 & a14874;
assign a15010 = ~a15008 & ~a14718;
assign a15012 = ~l894 & ~l892;
assign a15014 = a15012 & ~l890;
assign a15016 = l894 & ~l892;
assign a15018 = a15016 & ~l890;
assign a15020 = ~l894 & l892;
assign a15022 = a15020 & ~l890;
assign a15024 = l894 & l892;
assign a15026 = a15024 & ~l890;
assign a15028 = a15012 & l890;
assign a15030 = a15016 & l890;
assign a15032 = ~l898 & ~l896;
assign a15034 = l898 & ~l896;
assign a15036 = ~l898 & l896;
assign a15038 = l898 & l896;
assign a15040 = a15038 & ~l1312;
assign a15042 = a15040 & ~a15036;
assign a15044 = a15036 & ~l1298;
assign a15046 = ~a15044 & ~a15042;
assign a15048 = ~a15046 & ~a15034;
assign a15050 = a15034 & ~l1284;
assign a15052 = ~a15050 & ~a15048;
assign a15054 = ~a15052 & ~a15032;
assign a15056 = a15032 & ~l1270;
assign a15058 = ~a15056 & ~a15054;
assign a15060 = ~a15058 & a15030;
assign a15062 = a15060 & ~a15028;
assign a15064 = a15038 & ~l1228;
assign a15066 = a15064 & ~a15036;
assign a15068 = a15036 & ~l1214;
assign a15070 = ~a15068 & ~a15066;
assign a15072 = ~a15070 & ~a15034;
assign a15074 = a15034 & ~l1200;
assign a15076 = ~a15074 & ~a15072;
assign a15078 = ~a15076 & ~a15032;
assign a15080 = a15032 & ~l1186;
assign a15082 = ~a15080 & ~a15078;
assign a15084 = ~a15082 & a15028;
assign a15086 = ~a15084 & ~a15062;
assign a15088 = ~a15086 & ~a15026;
assign a15090 = a15038 & ~l1144;
assign a15092 = a15090 & ~a15036;
assign a15094 = a15036 & ~l1130;
assign a15096 = ~a15094 & ~a15092;
assign a15098 = ~a15096 & ~a15034;
assign a15100 = a15034 & ~l1116;
assign a15102 = ~a15100 & ~a15098;
assign a15104 = ~a15102 & ~a15032;
assign a15106 = a15032 & ~l1102;
assign a15108 = ~a15106 & ~a15104;
assign a15110 = ~a15108 & a15026;
assign a15112 = ~a15110 & ~a15088;
assign a15114 = ~a15112 & ~a15022;
assign a15116 = a15038 & ~l1060;
assign a15118 = a15116 & ~a15036;
assign a15120 = a15036 & ~l1046;
assign a15122 = ~a15120 & ~a15118;
assign a15124 = ~a15122 & ~a15034;
assign a15126 = a15034 & ~l1032;
assign a15128 = ~a15126 & ~a15124;
assign a15130 = ~a15128 & ~a15032;
assign a15132 = a15032 & ~l1018;
assign a15134 = ~a15132 & ~a15130;
assign a15136 = ~a15134 & a15022;
assign a15138 = ~a15136 & ~a15114;
assign a15140 = ~a15138 & ~a15018;
assign a15142 = a15038 & ~l976;
assign a15144 = a15142 & ~a15036;
assign a15146 = a15036 & ~l962;
assign a15148 = ~a15146 & ~a15144;
assign a15150 = ~a15148 & ~a15034;
assign a15152 = a15034 & ~l948;
assign a15154 = ~a15152 & ~a15150;
assign a15156 = ~a15154 & ~a15032;
assign a15158 = a15032 & ~l934;
assign a15160 = ~a15158 & ~a15156;
assign a15162 = ~a15160 & a15018;
assign a15164 = ~a15162 & ~a15140;
assign a15166 = a15164 & ~l1266;
assign a15168 = ~a15164 & l1266;
assign a15170 = ~a15168 & ~a15166;
assign a15172 = a15038 & l1314;
assign a15174 = a15172 & ~a15036;
assign a15176 = a15036 & l1300;
assign a15178 = ~a15176 & ~a15174;
assign a15180 = ~a15178 & ~a15034;
assign a15182 = a15034 & l1286;
assign a15184 = ~a15182 & ~a15180;
assign a15186 = ~a15184 & ~a15032;
assign a15188 = a15032 & l1272;
assign a15190 = ~a15188 & ~a15186;
assign a15192 = ~a15190 & a15030;
assign a15194 = a15192 & ~a15028;
assign a15196 = a15038 & l1230;
assign a15198 = a15196 & ~a15036;
assign a15200 = a15036 & l1216;
assign a15202 = ~a15200 & ~a15198;
assign a15204 = ~a15202 & ~a15034;
assign a15206 = a15034 & l1202;
assign a15208 = ~a15206 & ~a15204;
assign a15210 = ~a15208 & ~a15032;
assign a15212 = a15032 & l1188;
assign a15214 = ~a15212 & ~a15210;
assign a15216 = ~a15214 & a15028;
assign a15218 = ~a15216 & ~a15194;
assign a15220 = ~a15218 & ~a15026;
assign a15222 = a15038 & l1146;
assign a15224 = a15222 & ~a15036;
assign a15226 = a15036 & l1132;
assign a15228 = ~a15226 & ~a15224;
assign a15230 = ~a15228 & ~a15034;
assign a15232 = a15034 & l1118;
assign a15234 = ~a15232 & ~a15230;
assign a15236 = ~a15234 & ~a15032;
assign a15238 = a15032 & l1104;
assign a15240 = ~a15238 & ~a15236;
assign a15242 = ~a15240 & a15026;
assign a15244 = ~a15242 & ~a15220;
assign a15246 = ~a15244 & ~a15022;
assign a15248 = a15038 & l1062;
assign a15250 = a15248 & ~a15036;
assign a15252 = a15036 & l1048;
assign a15254 = ~a15252 & ~a15250;
assign a15256 = ~a15254 & ~a15034;
assign a15258 = a15034 & l1034;
assign a15260 = ~a15258 & ~a15256;
assign a15262 = ~a15260 & ~a15032;
assign a15264 = a15032 & l1020;
assign a15266 = ~a15264 & ~a15262;
assign a15268 = ~a15266 & a15022;
assign a15270 = ~a15268 & ~a15246;
assign a15272 = ~a15270 & ~a15018;
assign a15274 = a15038 & l978;
assign a15276 = a15274 & ~a15036;
assign a15278 = a15036 & l964;
assign a15280 = ~a15278 & ~a15276;
assign a15282 = ~a15280 & ~a15034;
assign a15284 = a15034 & l950;
assign a15286 = ~a15284 & ~a15282;
assign a15288 = ~a15286 & ~a15032;
assign a15290 = a15032 & l936;
assign a15292 = ~a15290 & ~a15288;
assign a15294 = ~a15292 & a15018;
assign a15296 = ~a15294 & ~a15272;
assign a15298 = a15296 & ~l1268;
assign a15300 = ~a15296 & l1268;
assign a15302 = ~a15300 & ~a15298;
assign a15304 = a15302 & a15170;
assign a15306 = ~a15304 & ~a15014;
assign a15308 = ~l904 & ~l902;
assign a15310 = a15308 & ~l900;
assign a15312 = l904 & ~l902;
assign a15314 = a15312 & ~l900;
assign a15316 = ~l904 & l902;
assign a15318 = a15316 & ~l900;
assign a15320 = l904 & l902;
assign a15322 = a15320 & ~l900;
assign a15324 = a15308 & l900;
assign a15326 = a15312 & l900;
assign a15328 = ~l908 & ~l906;
assign a15330 = l908 & ~l906;
assign a15332 = ~l908 & l906;
assign a15334 = l908 & l906;
assign a15336 = a15334 & ~l1312;
assign a15338 = a15336 & ~a15332;
assign a15340 = a15332 & ~l1298;
assign a15342 = ~a15340 & ~a15338;
assign a15344 = ~a15342 & ~a15330;
assign a15346 = a15330 & ~l1284;
assign a15348 = ~a15346 & ~a15344;
assign a15350 = ~a15348 & ~a15328;
assign a15352 = a15328 & ~l1270;
assign a15354 = ~a15352 & ~a15350;
assign a15356 = ~a15354 & a15326;
assign a15358 = a15356 & ~a15324;
assign a15360 = a15334 & ~l1228;
assign a15362 = a15360 & ~a15332;
assign a15364 = a15332 & ~l1214;
assign a15366 = ~a15364 & ~a15362;
assign a15368 = ~a15366 & ~a15330;
assign a15370 = a15330 & ~l1200;
assign a15372 = ~a15370 & ~a15368;
assign a15374 = ~a15372 & ~a15328;
assign a15376 = a15328 & ~l1186;
assign a15378 = ~a15376 & ~a15374;
assign a15380 = ~a15378 & a15324;
assign a15382 = ~a15380 & ~a15358;
assign a15384 = ~a15382 & ~a15322;
assign a15386 = a15334 & ~l1144;
assign a15388 = a15386 & ~a15332;
assign a15390 = a15332 & ~l1130;
assign a15392 = ~a15390 & ~a15388;
assign a15394 = ~a15392 & ~a15330;
assign a15396 = a15330 & ~l1116;
assign a15398 = ~a15396 & ~a15394;
assign a15400 = ~a15398 & ~a15328;
assign a15402 = a15328 & ~l1102;
assign a15404 = ~a15402 & ~a15400;
assign a15406 = ~a15404 & a15322;
assign a15408 = ~a15406 & ~a15384;
assign a15410 = ~a15408 & ~a15318;
assign a15412 = a15334 & ~l1060;
assign a15414 = a15412 & ~a15332;
assign a15416 = a15332 & ~l1046;
assign a15418 = ~a15416 & ~a15414;
assign a15420 = ~a15418 & ~a15330;
assign a15422 = a15330 & ~l1032;
assign a15424 = ~a15422 & ~a15420;
assign a15426 = ~a15424 & ~a15328;
assign a15428 = a15328 & ~l1018;
assign a15430 = ~a15428 & ~a15426;
assign a15432 = ~a15430 & a15318;
assign a15434 = ~a15432 & ~a15410;
assign a15436 = ~a15434 & ~a15314;
assign a15438 = a15334 & ~l976;
assign a15440 = a15438 & ~a15332;
assign a15442 = a15332 & ~l962;
assign a15444 = ~a15442 & ~a15440;
assign a15446 = ~a15444 & ~a15330;
assign a15448 = a15330 & ~l948;
assign a15450 = ~a15448 & ~a15446;
assign a15452 = ~a15450 & ~a15328;
assign a15454 = a15328 & ~l934;
assign a15456 = ~a15454 & ~a15452;
assign a15458 = ~a15456 & a15314;
assign a15460 = ~a15458 & ~a15436;
assign a15462 = a15460 & ~l1280;
assign a15464 = ~a15460 & l1280;
assign a15466 = ~a15464 & ~a15462;
assign a15468 = a15334 & l1314;
assign a15470 = a15468 & ~a15332;
assign a15472 = a15332 & l1300;
assign a15474 = ~a15472 & ~a15470;
assign a15476 = ~a15474 & ~a15330;
assign a15478 = a15330 & l1286;
assign a15480 = ~a15478 & ~a15476;
assign a15482 = ~a15480 & ~a15328;
assign a15484 = a15328 & l1272;
assign a15486 = ~a15484 & ~a15482;
assign a15488 = ~a15486 & a15326;
assign a15490 = a15488 & ~a15324;
assign a15492 = a15334 & l1230;
assign a15494 = a15492 & ~a15332;
assign a15496 = a15332 & l1216;
assign a15498 = ~a15496 & ~a15494;
assign a15500 = ~a15498 & ~a15330;
assign a15502 = a15330 & l1202;
assign a15504 = ~a15502 & ~a15500;
assign a15506 = ~a15504 & ~a15328;
assign a15508 = a15328 & l1188;
assign a15510 = ~a15508 & ~a15506;
assign a15512 = ~a15510 & a15324;
assign a15514 = ~a15512 & ~a15490;
assign a15516 = ~a15514 & ~a15322;
assign a15518 = a15334 & l1146;
assign a15520 = a15518 & ~a15332;
assign a15522 = a15332 & l1132;
assign a15524 = ~a15522 & ~a15520;
assign a15526 = ~a15524 & ~a15330;
assign a15528 = a15330 & l1118;
assign a15530 = ~a15528 & ~a15526;
assign a15532 = ~a15530 & ~a15328;
assign a15534 = a15328 & l1104;
assign a15536 = ~a15534 & ~a15532;
assign a15538 = ~a15536 & a15322;
assign a15540 = ~a15538 & ~a15516;
assign a15542 = ~a15540 & ~a15318;
assign a15544 = a15334 & l1062;
assign a15546 = a15544 & ~a15332;
assign a15548 = a15332 & l1048;
assign a15550 = ~a15548 & ~a15546;
assign a15552 = ~a15550 & ~a15330;
assign a15554 = a15330 & l1034;
assign a15556 = ~a15554 & ~a15552;
assign a15558 = ~a15556 & ~a15328;
assign a15560 = a15328 & l1020;
assign a15562 = ~a15560 & ~a15558;
assign a15564 = ~a15562 & a15318;
assign a15566 = ~a15564 & ~a15542;
assign a15568 = ~a15566 & ~a15314;
assign a15570 = a15334 & l978;
assign a15572 = a15570 & ~a15332;
assign a15574 = a15332 & l964;
assign a15576 = ~a15574 & ~a15572;
assign a15578 = ~a15576 & ~a15330;
assign a15580 = a15330 & l950;
assign a15582 = ~a15580 & ~a15578;
assign a15584 = ~a15582 & ~a15328;
assign a15586 = a15328 & l936;
assign a15588 = ~a15586 & ~a15584;
assign a15590 = ~a15588 & a15314;
assign a15592 = ~a15590 & ~a15568;
assign a15594 = a15592 & ~l1282;
assign a15596 = ~a15592 & l1282;
assign a15598 = ~a15596 & ~a15594;
assign a15600 = a15598 & a15466;
assign a15602 = ~a15600 & ~a15310;
assign a15604 = ~l914 & ~l912;
assign a15606 = a15604 & ~l910;
assign a15608 = l914 & ~l912;
assign a15610 = a15608 & ~l910;
assign a15612 = ~l914 & l912;
assign a15614 = a15612 & ~l910;
assign a15616 = l914 & l912;
assign a15618 = a15616 & ~l910;
assign a15620 = a15604 & l910;
assign a15622 = a15608 & l910;
assign a15624 = ~l918 & ~l916;
assign a15626 = l918 & ~l916;
assign a15628 = ~l918 & l916;
assign a15630 = l918 & l916;
assign a15632 = a15630 & ~l1312;
assign a15634 = a15632 & ~a15628;
assign a15636 = a15628 & ~l1298;
assign a15638 = ~a15636 & ~a15634;
assign a15640 = ~a15638 & ~a15626;
assign a15642 = a15626 & ~l1284;
assign a15644 = ~a15642 & ~a15640;
assign a15646 = ~a15644 & ~a15624;
assign a15648 = a15624 & ~l1270;
assign a15650 = ~a15648 & ~a15646;
assign a15652 = ~a15650 & a15622;
assign a15654 = a15652 & ~a15620;
assign a15656 = a15630 & ~l1228;
assign a15658 = a15656 & ~a15628;
assign a15660 = a15628 & ~l1214;
assign a15662 = ~a15660 & ~a15658;
assign a15664 = ~a15662 & ~a15626;
assign a15666 = a15626 & ~l1200;
assign a15668 = ~a15666 & ~a15664;
assign a15670 = ~a15668 & ~a15624;
assign a15672 = a15624 & ~l1186;
assign a15674 = ~a15672 & ~a15670;
assign a15676 = ~a15674 & a15620;
assign a15678 = ~a15676 & ~a15654;
assign a15680 = ~a15678 & ~a15618;
assign a15682 = a15630 & ~l1144;
assign a15684 = a15682 & ~a15628;
assign a15686 = a15628 & ~l1130;
assign a15688 = ~a15686 & ~a15684;
assign a15690 = ~a15688 & ~a15626;
assign a15692 = a15626 & ~l1116;
assign a15694 = ~a15692 & ~a15690;
assign a15696 = ~a15694 & ~a15624;
assign a15698 = a15624 & ~l1102;
assign a15700 = ~a15698 & ~a15696;
assign a15702 = ~a15700 & a15618;
assign a15704 = ~a15702 & ~a15680;
assign a15706 = ~a15704 & ~a15614;
assign a15708 = a15630 & ~l1060;
assign a15710 = a15708 & ~a15628;
assign a15712 = a15628 & ~l1046;
assign a15714 = ~a15712 & ~a15710;
assign a15716 = ~a15714 & ~a15626;
assign a15718 = a15626 & ~l1032;
assign a15720 = ~a15718 & ~a15716;
assign a15722 = ~a15720 & ~a15624;
assign a15724 = a15624 & ~l1018;
assign a15726 = ~a15724 & ~a15722;
assign a15728 = ~a15726 & a15614;
assign a15730 = ~a15728 & ~a15706;
assign a15732 = ~a15730 & ~a15610;
assign a15734 = a15630 & ~l976;
assign a15736 = a15734 & ~a15628;
assign a15738 = a15628 & ~l962;
assign a15740 = ~a15738 & ~a15736;
assign a15742 = ~a15740 & ~a15626;
assign a15744 = a15626 & ~l948;
assign a15746 = ~a15744 & ~a15742;
assign a15748 = ~a15746 & ~a15624;
assign a15750 = a15624 & ~l934;
assign a15752 = ~a15750 & ~a15748;
assign a15754 = ~a15752 & a15610;
assign a15756 = ~a15754 & ~a15732;
assign a15758 = a15756 & ~l1294;
assign a15760 = ~a15756 & l1294;
assign a15762 = ~a15760 & ~a15758;
assign a15764 = a15630 & l1314;
assign a15766 = a15764 & ~a15628;
assign a15768 = a15628 & l1300;
assign a15770 = ~a15768 & ~a15766;
assign a15772 = ~a15770 & ~a15626;
assign a15774 = a15626 & l1286;
assign a15776 = ~a15774 & ~a15772;
assign a15778 = ~a15776 & ~a15624;
assign a15780 = a15624 & l1272;
assign a15782 = ~a15780 & ~a15778;
assign a15784 = ~a15782 & a15622;
assign a15786 = a15784 & ~a15620;
assign a15788 = a15630 & l1230;
assign a15790 = a15788 & ~a15628;
assign a15792 = a15628 & l1216;
assign a15794 = ~a15792 & ~a15790;
assign a15796 = ~a15794 & ~a15626;
assign a15798 = a15626 & l1202;
assign a15800 = ~a15798 & ~a15796;
assign a15802 = ~a15800 & ~a15624;
assign a15804 = a15624 & l1188;
assign a15806 = ~a15804 & ~a15802;
assign a15808 = ~a15806 & a15620;
assign a15810 = ~a15808 & ~a15786;
assign a15812 = ~a15810 & ~a15618;
assign a15814 = a15630 & l1146;
assign a15816 = a15814 & ~a15628;
assign a15818 = a15628 & l1132;
assign a15820 = ~a15818 & ~a15816;
assign a15822 = ~a15820 & ~a15626;
assign a15824 = a15626 & l1118;
assign a15826 = ~a15824 & ~a15822;
assign a15828 = ~a15826 & ~a15624;
assign a15830 = a15624 & l1104;
assign a15832 = ~a15830 & ~a15828;
assign a15834 = ~a15832 & a15618;
assign a15836 = ~a15834 & ~a15812;
assign a15838 = ~a15836 & ~a15614;
assign a15840 = a15630 & l1062;
assign a15842 = a15840 & ~a15628;
assign a15844 = a15628 & l1048;
assign a15846 = ~a15844 & ~a15842;
assign a15848 = ~a15846 & ~a15626;
assign a15850 = a15626 & l1034;
assign a15852 = ~a15850 & ~a15848;
assign a15854 = ~a15852 & ~a15624;
assign a15856 = a15624 & l1020;
assign a15858 = ~a15856 & ~a15854;
assign a15860 = ~a15858 & a15614;
assign a15862 = ~a15860 & ~a15838;
assign a15864 = ~a15862 & ~a15610;
assign a15866 = a15630 & l978;
assign a15868 = a15866 & ~a15628;
assign a15870 = a15628 & l964;
assign a15872 = ~a15870 & ~a15868;
assign a15874 = ~a15872 & ~a15626;
assign a15876 = a15626 & l950;
assign a15878 = ~a15876 & ~a15874;
assign a15880 = ~a15878 & ~a15624;
assign a15882 = a15624 & l936;
assign a15884 = ~a15882 & ~a15880;
assign a15886 = ~a15884 & a15610;
assign a15888 = ~a15886 & ~a15864;
assign a15890 = a15888 & ~l1296;
assign a15892 = ~a15888 & l1296;
assign a15894 = ~a15892 & ~a15890;
assign a15896 = a15894 & a15762;
assign a15898 = ~a15896 & ~a15606;
assign a15900 = ~l924 & ~l922;
assign a15902 = a15900 & ~l920;
assign a15904 = l924 & ~l922;
assign a15906 = a15904 & ~l920;
assign a15908 = ~l924 & l922;
assign a15910 = a15908 & ~l920;
assign a15912 = l924 & l922;
assign a15914 = a15912 & ~l920;
assign a15916 = a15900 & l920;
assign a15918 = a15904 & l920;
assign a15920 = ~l928 & ~l926;
assign a15922 = l928 & ~l926;
assign a15924 = ~l928 & l926;
assign a15926 = l928 & l926;
assign a15928 = a15926 & ~l1312;
assign a15930 = a15928 & ~a15924;
assign a15932 = a15924 & ~l1298;
assign a15934 = ~a15932 & ~a15930;
assign a15936 = ~a15934 & ~a15922;
assign a15938 = a15922 & ~l1284;
assign a15940 = ~a15938 & ~a15936;
assign a15942 = ~a15940 & ~a15920;
assign a15944 = a15920 & ~l1270;
assign a15946 = ~a15944 & ~a15942;
assign a15948 = ~a15946 & a15918;
assign a15950 = a15948 & ~a15916;
assign a15952 = a15926 & ~l1228;
assign a15954 = a15952 & ~a15924;
assign a15956 = a15924 & ~l1214;
assign a15958 = ~a15956 & ~a15954;
assign a15960 = ~a15958 & ~a15922;
assign a15962 = a15922 & ~l1200;
assign a15964 = ~a15962 & ~a15960;
assign a15966 = ~a15964 & ~a15920;
assign a15968 = a15920 & ~l1186;
assign a15970 = ~a15968 & ~a15966;
assign a15972 = ~a15970 & a15916;
assign a15974 = ~a15972 & ~a15950;
assign a15976 = ~a15974 & ~a15914;
assign a15978 = a15926 & ~l1144;
assign a15980 = a15978 & ~a15924;
assign a15982 = a15924 & ~l1130;
assign a15984 = ~a15982 & ~a15980;
assign a15986 = ~a15984 & ~a15922;
assign a15988 = a15922 & ~l1116;
assign a15990 = ~a15988 & ~a15986;
assign a15992 = ~a15990 & ~a15920;
assign a15994 = a15920 & ~l1102;
assign a15996 = ~a15994 & ~a15992;
assign a15998 = ~a15996 & a15914;
assign a16000 = ~a15998 & ~a15976;
assign a16002 = ~a16000 & ~a15910;
assign a16004 = a15926 & ~l1060;
assign a16006 = a16004 & ~a15924;
assign a16008 = a15924 & ~l1046;
assign a16010 = ~a16008 & ~a16006;
assign a16012 = ~a16010 & ~a15922;
assign a16014 = a15922 & ~l1032;
assign a16016 = ~a16014 & ~a16012;
assign a16018 = ~a16016 & ~a15920;
assign a16020 = a15920 & ~l1018;
assign a16022 = ~a16020 & ~a16018;
assign a16024 = ~a16022 & a15910;
assign a16026 = ~a16024 & ~a16002;
assign a16028 = ~a16026 & ~a15906;
assign a16030 = a15926 & ~l976;
assign a16032 = a16030 & ~a15924;
assign a16034 = a15924 & ~l962;
assign a16036 = ~a16034 & ~a16032;
assign a16038 = ~a16036 & ~a15922;
assign a16040 = a15922 & ~l948;
assign a16042 = ~a16040 & ~a16038;
assign a16044 = ~a16042 & ~a15920;
assign a16046 = a15920 & ~l934;
assign a16048 = ~a16046 & ~a16044;
assign a16050 = ~a16048 & a15906;
assign a16052 = ~a16050 & ~a16028;
assign a16054 = a16052 & ~l1308;
assign a16056 = ~a16052 & l1308;
assign a16058 = ~a16056 & ~a16054;
assign a16060 = a15926 & l1314;
assign a16062 = a16060 & ~a15924;
assign a16064 = a15924 & l1300;
assign a16066 = ~a16064 & ~a16062;
assign a16068 = ~a16066 & ~a15922;
assign a16070 = a15922 & l1286;
assign a16072 = ~a16070 & ~a16068;
assign a16074 = ~a16072 & ~a15920;
assign a16076 = a15920 & l1272;
assign a16078 = ~a16076 & ~a16074;
assign a16080 = ~a16078 & a15918;
assign a16082 = a16080 & ~a15916;
assign a16084 = a15926 & l1230;
assign a16086 = a16084 & ~a15924;
assign a16088 = a15924 & l1216;
assign a16090 = ~a16088 & ~a16086;
assign a16092 = ~a16090 & ~a15922;
assign a16094 = a15922 & l1202;
assign a16096 = ~a16094 & ~a16092;
assign a16098 = ~a16096 & ~a15920;
assign a16100 = a15920 & l1188;
assign a16102 = ~a16100 & ~a16098;
assign a16104 = ~a16102 & a15916;
assign a16106 = ~a16104 & ~a16082;
assign a16108 = ~a16106 & ~a15914;
assign a16110 = a15926 & l1146;
assign a16112 = a16110 & ~a15924;
assign a16114 = a15924 & l1132;
assign a16116 = ~a16114 & ~a16112;
assign a16118 = ~a16116 & ~a15922;
assign a16120 = a15922 & l1118;
assign a16122 = ~a16120 & ~a16118;
assign a16124 = ~a16122 & ~a15920;
assign a16126 = a15920 & l1104;
assign a16128 = ~a16126 & ~a16124;
assign a16130 = ~a16128 & a15914;
assign a16132 = ~a16130 & ~a16108;
assign a16134 = ~a16132 & ~a15910;
assign a16136 = a15926 & l1062;
assign a16138 = a16136 & ~a15924;
assign a16140 = a15924 & l1048;
assign a16142 = ~a16140 & ~a16138;
assign a16144 = ~a16142 & ~a15922;
assign a16146 = a15922 & l1034;
assign a16148 = ~a16146 & ~a16144;
assign a16150 = ~a16148 & ~a15920;
assign a16152 = a15920 & l1020;
assign a16154 = ~a16152 & ~a16150;
assign a16156 = ~a16154 & a15910;
assign a16158 = ~a16156 & ~a16134;
assign a16160 = ~a16158 & ~a15906;
assign a16162 = a15926 & l978;
assign a16164 = a16162 & ~a15924;
assign a16166 = a15924 & l964;
assign a16168 = ~a16166 & ~a16164;
assign a16170 = ~a16168 & ~a15922;
assign a16172 = a15922 & l950;
assign a16174 = ~a16172 & ~a16170;
assign a16176 = ~a16174 & ~a15920;
assign a16178 = a15920 & l936;
assign a16180 = ~a16178 & ~a16176;
assign a16182 = ~a16180 & a15906;
assign a16184 = ~a16182 & ~a16160;
assign a16186 = a16184 & ~l1310;
assign a16188 = ~a16184 & l1310;
assign a16190 = ~a16188 & ~a16186;
assign a16192 = a16190 & a16058;
assign a16194 = ~a16192 & ~a15902;
assign a16196 = a15920 & a15906;
assign a16198 = ~a16196 & a10302;
assign a16200 = a16198 & ~a10300;
assign a16202 = a15624 & a15610;
assign a16204 = ~a16202 & a10300;
assign a16206 = ~a16204 & ~a16200;
assign a16208 = ~a16206 & ~a10298;
assign a16210 = a15328 & a15314;
assign a16212 = ~a16210 & a10298;
assign a16214 = ~a16212 & ~a16208;
assign a16216 = ~a16214 & ~a10296;
assign a16218 = a15032 & a15018;
assign a16220 = ~a16218 & a10296;
assign a16222 = ~a16220 & ~a16216;
assign a16224 = ~a16222 & a10294;
assign a16226 = a16224 & ~a10292;
assign a16228 = a14736 & a14722;
assign a16230 = ~a16228 & a10302;
assign a16232 = a16230 & ~a10300;
assign a16234 = a14440 & a14426;
assign a16236 = ~a16234 & a10300;
assign a16238 = ~a16236 & ~a16232;
assign a16240 = ~a16238 & ~a10298;
assign a16242 = a14144 & a14130;
assign a16244 = ~a16242 & a10298;
assign a16246 = ~a16244 & ~a16240;
assign a16248 = ~a16246 & ~a10296;
assign a16250 = a13848 & a13834;
assign a16252 = ~a16250 & a10296;
assign a16254 = ~a16252 & ~a16248;
assign a16256 = ~a16254 & a10292;
assign a16258 = ~a16256 & ~a16226;
assign a16260 = ~a16258 & ~a10290;
assign a16262 = a13552 & a13538;
assign a16264 = ~a16262 & a10302;
assign a16266 = a16264 & ~a10300;
assign a16268 = a13256 & a13242;
assign a16270 = ~a16268 & a10300;
assign a16272 = ~a16270 & ~a16266;
assign a16274 = ~a16272 & ~a10298;
assign a16276 = a12960 & a12946;
assign a16278 = ~a16276 & a10298;
assign a16280 = ~a16278 & ~a16274;
assign a16282 = ~a16280 & ~a10296;
assign a16284 = a12664 & a12650;
assign a16286 = ~a16284 & a10296;
assign a16288 = ~a16286 & ~a16282;
assign a16290 = ~a16288 & a10290;
assign a16292 = ~a16290 & ~a16260;
assign a16294 = ~a16292 & ~a10286;
assign a16296 = a12368 & a12354;
assign a16298 = ~a16296 & a10302;
assign a16300 = a16298 & ~a10300;
assign a16302 = a12072 & a12058;
assign a16304 = ~a16302 & a10300;
assign a16306 = ~a16304 & ~a16300;
assign a16308 = ~a16306 & ~a10298;
assign a16310 = a11776 & a11762;
assign a16312 = ~a16310 & a10298;
assign a16314 = ~a16312 & ~a16308;
assign a16316 = ~a16314 & ~a10296;
assign a16318 = a11480 & a11466;
assign a16320 = ~a16318 & a10296;
assign a16322 = ~a16320 & ~a16316;
assign a16324 = ~a16322 & a10286;
assign a16326 = ~a16324 & ~a16294;
assign a16328 = ~a16326 & ~a10282;
assign a16330 = a11184 & a11170;
assign a16332 = ~a16330 & a10302;
assign a16334 = a16332 & ~a10300;
assign a16336 = a10888 & a10874;
assign a16338 = ~a16336 & a10300;
assign a16340 = ~a16338 & ~a16334;
assign a16342 = ~a16340 & ~a10298;
assign a16344 = a10592 & a10578;
assign a16346 = ~a16344 & a10298;
assign a16348 = ~a16346 & ~a16342;
assign a16350 = ~a16348 & ~a10296;
assign a16352 = a10296 & ~a10282;
assign a16354 = ~a16352 & ~a16350;
assign a16356 = ~a16354 & a10282;
assign a16358 = ~a16356 & ~a16328;
assign a16360 = a15922 & a15906;
assign a16362 = ~a16360 & a10598;
assign a16364 = a16362 & ~a10596;
assign a16366 = a15626 & a15610;
assign a16368 = ~a16366 & a10596;
assign a16370 = ~a16368 & ~a16364;
assign a16372 = ~a16370 & ~a10594;
assign a16374 = a15330 & a15314;
assign a16376 = ~a16374 & a10594;
assign a16378 = ~a16376 & ~a16372;
assign a16380 = ~a16378 & ~a10592;
assign a16382 = a15034 & a15018;
assign a16384 = ~a16382 & a10592;
assign a16386 = ~a16384 & ~a16380;
assign a16388 = ~a16386 & a10590;
assign a16390 = a16388 & ~a10588;
assign a16392 = a14738 & a14722;
assign a16394 = ~a16392 & a10598;
assign a16396 = a16394 & ~a10596;
assign a16398 = a14442 & a14426;
assign a16400 = ~a16398 & a10596;
assign a16402 = ~a16400 & ~a16396;
assign a16404 = ~a16402 & ~a10594;
assign a16406 = a14146 & a14130;
assign a16408 = ~a16406 & a10594;
assign a16410 = ~a16408 & ~a16404;
assign a16412 = ~a16410 & ~a10592;
assign a16414 = a13850 & a13834;
assign a16416 = ~a16414 & a10592;
assign a16418 = ~a16416 & ~a16412;
assign a16420 = ~a16418 & a10588;
assign a16422 = ~a16420 & ~a16390;
assign a16424 = ~a16422 & ~a10586;
assign a16426 = a13554 & a13538;
assign a16428 = ~a16426 & a10598;
assign a16430 = a16428 & ~a10596;
assign a16432 = a13258 & a13242;
assign a16434 = ~a16432 & a10596;
assign a16436 = ~a16434 & ~a16430;
assign a16438 = ~a16436 & ~a10594;
assign a16440 = a12962 & a12946;
assign a16442 = ~a16440 & a10594;
assign a16444 = ~a16442 & ~a16438;
assign a16446 = ~a16444 & ~a10592;
assign a16448 = a12666 & a12650;
assign a16450 = ~a16448 & a10592;
assign a16452 = ~a16450 & ~a16446;
assign a16454 = ~a16452 & a10586;
assign a16456 = ~a16454 & ~a16424;
assign a16458 = ~a16456 & ~a10582;
assign a16460 = a12370 & a12354;
assign a16462 = ~a16460 & a10598;
assign a16464 = a16462 & ~a10596;
assign a16466 = a12074 & a12058;
assign a16468 = ~a16466 & a10596;
assign a16470 = ~a16468 & ~a16464;
assign a16472 = ~a16470 & ~a10594;
assign a16474 = a11778 & a11762;
assign a16476 = ~a16474 & a10594;
assign a16478 = ~a16476 & ~a16472;
assign a16480 = ~a16478 & ~a10592;
assign a16482 = a11482 & a11466;
assign a16484 = ~a16482 & a10592;
assign a16486 = ~a16484 & ~a16480;
assign a16488 = ~a16486 & a10582;
assign a16490 = ~a16488 & ~a16458;
assign a16492 = ~a16490 & ~a10578;
assign a16494 = a11186 & a11170;
assign a16496 = ~a16494 & a10598;
assign a16498 = a16496 & ~a10596;
assign a16500 = a10890 & a10874;
assign a16502 = ~a16500 & a10596;
assign a16504 = ~a16502 & ~a16498;
assign a16506 = ~a16504 & ~a10594;
assign a16508 = a10594 & ~a10578;
assign a16510 = ~a16508 & ~a16506;
assign a16512 = ~a16510 & ~a10592;
assign a16514 = a10298 & a10282;
assign a16516 = ~a16514 & a10592;
assign a16518 = ~a16516 & ~a16512;
assign a16520 = ~a16518 & a10578;
assign a16522 = ~a16520 & ~a16492;
assign a16524 = a15924 & a15906;
assign a16526 = ~a16524 & a10894;
assign a16528 = a16526 & ~a10892;
assign a16530 = a15628 & a15610;
assign a16532 = ~a16530 & a10892;
assign a16534 = ~a16532 & ~a16528;
assign a16536 = ~a16534 & ~a10890;
assign a16538 = a15332 & a15314;
assign a16540 = ~a16538 & a10890;
assign a16542 = ~a16540 & ~a16536;
assign a16544 = ~a16542 & ~a10888;
assign a16546 = a15036 & a15018;
assign a16548 = ~a16546 & a10888;
assign a16550 = ~a16548 & ~a16544;
assign a16552 = ~a16550 & a10886;
assign a16554 = a16552 & ~a10884;
assign a16556 = a14740 & a14722;
assign a16558 = ~a16556 & a10894;
assign a16560 = a16558 & ~a10892;
assign a16562 = a14444 & a14426;
assign a16564 = ~a16562 & a10892;
assign a16566 = ~a16564 & ~a16560;
assign a16568 = ~a16566 & ~a10890;
assign a16570 = a14148 & a14130;
assign a16572 = ~a16570 & a10890;
assign a16574 = ~a16572 & ~a16568;
assign a16576 = ~a16574 & ~a10888;
assign a16578 = a13852 & a13834;
assign a16580 = ~a16578 & a10888;
assign a16582 = ~a16580 & ~a16576;
assign a16584 = ~a16582 & a10884;
assign a16586 = ~a16584 & ~a16554;
assign a16588 = ~a16586 & ~a10882;
assign a16590 = a13556 & a13538;
assign a16592 = ~a16590 & a10894;
assign a16594 = a16592 & ~a10892;
assign a16596 = a13260 & a13242;
assign a16598 = ~a16596 & a10892;
assign a16600 = ~a16598 & ~a16594;
assign a16602 = ~a16600 & ~a10890;
assign a16604 = a12964 & a12946;
assign a16606 = ~a16604 & a10890;
assign a16608 = ~a16606 & ~a16602;
assign a16610 = ~a16608 & ~a10888;
assign a16612 = a12668 & a12650;
assign a16614 = ~a16612 & a10888;
assign a16616 = ~a16614 & ~a16610;
assign a16618 = ~a16616 & a10882;
assign a16620 = ~a16618 & ~a16588;
assign a16622 = ~a16620 & ~a10878;
assign a16624 = a12372 & a12354;
assign a16626 = ~a16624 & a10894;
assign a16628 = a16626 & ~a10892;
assign a16630 = a12076 & a12058;
assign a16632 = ~a16630 & a10892;
assign a16634 = ~a16632 & ~a16628;
assign a16636 = ~a16634 & ~a10890;
assign a16638 = a11780 & a11762;
assign a16640 = ~a16638 & a10890;
assign a16642 = ~a16640 & ~a16636;
assign a16644 = ~a16642 & ~a10888;
assign a16646 = a11484 & a11466;
assign a16648 = ~a16646 & a10888;
assign a16650 = ~a16648 & ~a16644;
assign a16652 = ~a16650 & a10878;
assign a16654 = ~a16652 & ~a16622;
assign a16656 = ~a16654 & ~a10874;
assign a16658 = a11188 & a11170;
assign a16660 = ~a16658 & a10894;
assign a16662 = a16660 & ~a10892;
assign a16664 = a10892 & ~a10874;
assign a16666 = ~a16664 & ~a16662;
assign a16668 = ~a16666 & ~a10890;
assign a16670 = a10596 & a10578;
assign a16672 = ~a16670 & a10890;
assign a16674 = ~a16672 & ~a16668;
assign a16676 = ~a16674 & ~a10888;
assign a16678 = a10300 & a10282;
assign a16680 = ~a16678 & a10888;
assign a16682 = ~a16680 & ~a16676;
assign a16684 = ~a16682 & a10874;
assign a16686 = ~a16684 & ~a16656;
assign a16688 = a15926 & a15906;
assign a16690 = ~a16688 & a11190;
assign a16692 = a16690 & ~a11188;
assign a16694 = a15630 & a15610;
assign a16696 = ~a16694 & a11188;
assign a16698 = ~a16696 & ~a16692;
assign a16700 = ~a16698 & ~a11186;
assign a16702 = a15334 & a15314;
assign a16704 = ~a16702 & a11186;
assign a16706 = ~a16704 & ~a16700;
assign a16708 = ~a16706 & ~a11184;
assign a16710 = a15038 & a15018;
assign a16712 = ~a16710 & a11184;
assign a16714 = ~a16712 & ~a16708;
assign a16716 = ~a16714 & a11182;
assign a16718 = a16716 & ~a11180;
assign a16720 = a14742 & a14722;
assign a16722 = ~a16720 & a11190;
assign a16724 = a16722 & ~a11188;
assign a16726 = a14446 & a14426;
assign a16728 = ~a16726 & a11188;
assign a16730 = ~a16728 & ~a16724;
assign a16732 = ~a16730 & ~a11186;
assign a16734 = a14150 & a14130;
assign a16736 = ~a16734 & a11186;
assign a16738 = ~a16736 & ~a16732;
assign a16740 = ~a16738 & ~a11184;
assign a16742 = a13854 & a13834;
assign a16744 = ~a16742 & a11184;
assign a16746 = ~a16744 & ~a16740;
assign a16748 = ~a16746 & a11180;
assign a16750 = ~a16748 & ~a16718;
assign a16752 = ~a16750 & ~a11178;
assign a16754 = a13558 & a13538;
assign a16756 = ~a16754 & a11190;
assign a16758 = a16756 & ~a11188;
assign a16760 = a13262 & a13242;
assign a16762 = ~a16760 & a11188;
assign a16764 = ~a16762 & ~a16758;
assign a16766 = ~a16764 & ~a11186;
assign a16768 = a12966 & a12946;
assign a16770 = ~a16768 & a11186;
assign a16772 = ~a16770 & ~a16766;
assign a16774 = ~a16772 & ~a11184;
assign a16776 = a12670 & a12650;
assign a16778 = ~a16776 & a11184;
assign a16780 = ~a16778 & ~a16774;
assign a16782 = ~a16780 & a11178;
assign a16784 = ~a16782 & ~a16752;
assign a16786 = ~a16784 & ~a11174;
assign a16788 = a12374 & a12354;
assign a16790 = ~a16788 & a11190;
assign a16792 = a16790 & ~a11188;
assign a16794 = a12078 & a12058;
assign a16796 = ~a16794 & a11188;
assign a16798 = ~a16796 & ~a16792;
assign a16800 = ~a16798 & ~a11186;
assign a16802 = a11782 & a11762;
assign a16804 = ~a16802 & a11186;
assign a16806 = ~a16804 & ~a16800;
assign a16808 = ~a16806 & ~a11184;
assign a16810 = a11486 & a11466;
assign a16812 = ~a16810 & a11184;
assign a16814 = ~a16812 & ~a16808;
assign a16816 = ~a16814 & a11174;
assign a16818 = ~a16816 & ~a16786;
assign a16820 = ~a16818 & ~a11170;
assign a16822 = a11190 & ~a11170;
assign a16824 = a16822 & ~a11188;
assign a16826 = a10894 & a10874;
assign a16828 = ~a16826 & a11188;
assign a16830 = ~a16828 & ~a16824;
assign a16832 = ~a16830 & ~a11186;
assign a16834 = a10598 & a10578;
assign a16836 = ~a16834 & a11186;
assign a16838 = ~a16836 & ~a16832;
assign a16840 = ~a16838 & ~a11184;
assign a16842 = a10302 & a10282;
assign a16844 = ~a16842 & a11184;
assign a16846 = ~a16844 & ~a16840;
assign a16848 = ~a16846 & a11170;
assign a16850 = ~a16848 & ~a16820;
assign a16852 = a15920 & a15910;
assign a16854 = ~a16852 & a11486;
assign a16856 = a16854 & ~a11484;
assign a16858 = a15624 & a15614;
assign a16860 = ~a16858 & a11484;
assign a16862 = ~a16860 & ~a16856;
assign a16864 = ~a16862 & ~a11482;
assign a16866 = a15328 & a15318;
assign a16868 = ~a16866 & a11482;
assign a16870 = ~a16868 & ~a16864;
assign a16872 = ~a16870 & ~a11480;
assign a16874 = a15032 & a15022;
assign a16876 = ~a16874 & a11480;
assign a16878 = ~a16876 & ~a16872;
assign a16880 = ~a16878 & a11478;
assign a16882 = a16880 & ~a11476;
assign a16884 = a14736 & a14726;
assign a16886 = ~a16884 & a11486;
assign a16888 = a16886 & ~a11484;
assign a16890 = a14440 & a14430;
assign a16892 = ~a16890 & a11484;
assign a16894 = ~a16892 & ~a16888;
assign a16896 = ~a16894 & ~a11482;
assign a16898 = a14144 & a14134;
assign a16900 = ~a16898 & a11482;
assign a16902 = ~a16900 & ~a16896;
assign a16904 = ~a16902 & ~a11480;
assign a16906 = a13848 & a13838;
assign a16908 = ~a16906 & a11480;
assign a16910 = ~a16908 & ~a16904;
assign a16912 = ~a16910 & a11476;
assign a16914 = ~a16912 & ~a16882;
assign a16916 = ~a16914 & ~a11474;
assign a16918 = a13552 & a13542;
assign a16920 = ~a16918 & a11486;
assign a16922 = a16920 & ~a11484;
assign a16924 = a13256 & a13246;
assign a16926 = ~a16924 & a11484;
assign a16928 = ~a16926 & ~a16922;
assign a16930 = ~a16928 & ~a11482;
assign a16932 = a12960 & a12950;
assign a16934 = ~a16932 & a11482;
assign a16936 = ~a16934 & ~a16930;
assign a16938 = ~a16936 & ~a11480;
assign a16940 = a12664 & a12654;
assign a16942 = ~a16940 & a11480;
assign a16944 = ~a16942 & ~a16938;
assign a16946 = ~a16944 & a11474;
assign a16948 = ~a16946 & ~a16916;
assign a16950 = ~a16948 & ~a11470;
assign a16952 = a12368 & a12358;
assign a16954 = ~a16952 & a11486;
assign a16956 = a16954 & ~a11484;
assign a16958 = a12072 & a12062;
assign a16960 = ~a16958 & a11484;
assign a16962 = ~a16960 & ~a16956;
assign a16964 = ~a16962 & ~a11482;
assign a16966 = a11776 & a11766;
assign a16968 = ~a16966 & a11482;
assign a16970 = ~a16968 & ~a16964;
assign a16972 = ~a16970 & ~a11480;
assign a16974 = a11480 & ~a11470;
assign a16976 = ~a16974 & ~a16972;
assign a16978 = ~a16976 & a11470;
assign a16980 = ~a16978 & ~a16950;
assign a16982 = ~a16980 & ~a11466;
assign a16984 = a11184 & a11174;
assign a16986 = ~a16984 & a11486;
assign a16988 = a16986 & ~a11484;
assign a16990 = a10888 & a10878;
assign a16992 = ~a16990 & a11484;
assign a16994 = ~a16992 & ~a16988;
assign a16996 = ~a16994 & ~a11482;
assign a16998 = a10592 & a10582;
assign a17000 = ~a16998 & a11482;
assign a17002 = ~a17000 & ~a16996;
assign a17004 = ~a17002 & ~a11480;
assign a17006 = a10296 & a10286;
assign a17008 = ~a17006 & a11480;
assign a17010 = ~a17008 & ~a17004;
assign a17012 = ~a17010 & a11466;
assign a17014 = ~a17012 & ~a16982;
assign a17016 = a15922 & a15910;
assign a17018 = ~a17016 & a11782;
assign a17020 = a17018 & ~a11780;
assign a17022 = a15626 & a15614;
assign a17024 = ~a17022 & a11780;
assign a17026 = ~a17024 & ~a17020;
assign a17028 = ~a17026 & ~a11778;
assign a17030 = a15330 & a15318;
assign a17032 = ~a17030 & a11778;
assign a17034 = ~a17032 & ~a17028;
assign a17036 = ~a17034 & ~a11776;
assign a17038 = a15034 & a15022;
assign a17040 = ~a17038 & a11776;
assign a17042 = ~a17040 & ~a17036;
assign a17044 = ~a17042 & a11774;
assign a17046 = a17044 & ~a11772;
assign a17048 = a14738 & a14726;
assign a17050 = ~a17048 & a11782;
assign a17052 = a17050 & ~a11780;
assign a17054 = a14442 & a14430;
assign a17056 = ~a17054 & a11780;
assign a17058 = ~a17056 & ~a17052;
assign a17060 = ~a17058 & ~a11778;
assign a17062 = a14146 & a14134;
assign a17064 = ~a17062 & a11778;
assign a17066 = ~a17064 & ~a17060;
assign a17068 = ~a17066 & ~a11776;
assign a17070 = a13850 & a13838;
assign a17072 = ~a17070 & a11776;
assign a17074 = ~a17072 & ~a17068;
assign a17076 = ~a17074 & a11772;
assign a17078 = ~a17076 & ~a17046;
assign a17080 = ~a17078 & ~a11770;
assign a17082 = a13554 & a13542;
assign a17084 = ~a17082 & a11782;
assign a17086 = a17084 & ~a11780;
assign a17088 = a13258 & a13246;
assign a17090 = ~a17088 & a11780;
assign a17092 = ~a17090 & ~a17086;
assign a17094 = ~a17092 & ~a11778;
assign a17096 = a12962 & a12950;
assign a17098 = ~a17096 & a11778;
assign a17100 = ~a17098 & ~a17094;
assign a17102 = ~a17100 & ~a11776;
assign a17104 = a12666 & a12654;
assign a17106 = ~a17104 & a11776;
assign a17108 = ~a17106 & ~a17102;
assign a17110 = ~a17108 & a11770;
assign a17112 = ~a17110 & ~a17080;
assign a17114 = ~a17112 & ~a11766;
assign a17116 = a12370 & a12358;
assign a17118 = ~a17116 & a11782;
assign a17120 = a17118 & ~a11780;
assign a17122 = a12074 & a12062;
assign a17124 = ~a17122 & a11780;
assign a17126 = ~a17124 & ~a17120;
assign a17128 = ~a17126 & ~a11778;
assign a17130 = a11778 & ~a11766;
assign a17132 = ~a17130 & ~a17128;
assign a17134 = ~a17132 & ~a11776;
assign a17136 = a11482 & a11470;
assign a17138 = ~a17136 & a11776;
assign a17140 = ~a17138 & ~a17134;
assign a17142 = ~a17140 & a11766;
assign a17144 = ~a17142 & ~a17114;
assign a17146 = ~a17144 & ~a11762;
assign a17148 = a11186 & a11174;
assign a17150 = ~a17148 & a11782;
assign a17152 = a17150 & ~a11780;
assign a17154 = a10890 & a10878;
assign a17156 = ~a17154 & a11780;
assign a17158 = ~a17156 & ~a17152;
assign a17160 = ~a17158 & ~a11778;
assign a17162 = a10594 & a10582;
assign a17164 = ~a17162 & a11778;
assign a17166 = ~a17164 & ~a17160;
assign a17168 = ~a17166 & ~a11776;
assign a17170 = a10298 & a10286;
assign a17172 = ~a17170 & a11776;
assign a17174 = ~a17172 & ~a17168;
assign a17176 = ~a17174 & a11762;
assign a17178 = ~a17176 & ~a17146;
assign a17180 = a15924 & a15910;
assign a17182 = ~a17180 & a12078;
assign a17184 = a17182 & ~a12076;
assign a17186 = a15628 & a15614;
assign a17188 = ~a17186 & a12076;
assign a17190 = ~a17188 & ~a17184;
assign a17192 = ~a17190 & ~a12074;
assign a17194 = a15332 & a15318;
assign a17196 = ~a17194 & a12074;
assign a17198 = ~a17196 & ~a17192;
assign a17200 = ~a17198 & ~a12072;
assign a17202 = a15036 & a15022;
assign a17204 = ~a17202 & a12072;
assign a17206 = ~a17204 & ~a17200;
assign a17208 = ~a17206 & a12070;
assign a17210 = a17208 & ~a12068;
assign a17212 = a14740 & a14726;
assign a17214 = ~a17212 & a12078;
assign a17216 = a17214 & ~a12076;
assign a17218 = a14444 & a14430;
assign a17220 = ~a17218 & a12076;
assign a17222 = ~a17220 & ~a17216;
assign a17224 = ~a17222 & ~a12074;
assign a17226 = a14148 & a14134;
assign a17228 = ~a17226 & a12074;
assign a17230 = ~a17228 & ~a17224;
assign a17232 = ~a17230 & ~a12072;
assign a17234 = a13852 & a13838;
assign a17236 = ~a17234 & a12072;
assign a17238 = ~a17236 & ~a17232;
assign a17240 = ~a17238 & a12068;
assign a17242 = ~a17240 & ~a17210;
assign a17244 = ~a17242 & ~a12066;
assign a17246 = a13556 & a13542;
assign a17248 = ~a17246 & a12078;
assign a17250 = a17248 & ~a12076;
assign a17252 = a13260 & a13246;
assign a17254 = ~a17252 & a12076;
assign a17256 = ~a17254 & ~a17250;
assign a17258 = ~a17256 & ~a12074;
assign a17260 = a12964 & a12950;
assign a17262 = ~a17260 & a12074;
assign a17264 = ~a17262 & ~a17258;
assign a17266 = ~a17264 & ~a12072;
assign a17268 = a12668 & a12654;
assign a17270 = ~a17268 & a12072;
assign a17272 = ~a17270 & ~a17266;
assign a17274 = ~a17272 & a12066;
assign a17276 = ~a17274 & ~a17244;
assign a17278 = ~a17276 & ~a12062;
assign a17280 = a12372 & a12358;
assign a17282 = ~a17280 & a12078;
assign a17284 = a17282 & ~a12076;
assign a17286 = a12076 & ~a12062;
assign a17288 = ~a17286 & ~a17284;
assign a17290 = ~a17288 & ~a12074;
assign a17292 = a11780 & a11766;
assign a17294 = ~a17292 & a12074;
assign a17296 = ~a17294 & ~a17290;
assign a17298 = ~a17296 & ~a12072;
assign a17300 = a11484 & a11470;
assign a17302 = ~a17300 & a12072;
assign a17304 = ~a17302 & ~a17298;
assign a17306 = ~a17304 & a12062;
assign a17308 = ~a17306 & ~a17278;
assign a17310 = ~a17308 & ~a12058;
assign a17312 = a11188 & a11174;
assign a17314 = ~a17312 & a12078;
assign a17316 = a17314 & ~a12076;
assign a17318 = a10892 & a10878;
assign a17320 = ~a17318 & a12076;
assign a17322 = ~a17320 & ~a17316;
assign a17324 = ~a17322 & ~a12074;
assign a17326 = a10596 & a10582;
assign a17328 = ~a17326 & a12074;
assign a17330 = ~a17328 & ~a17324;
assign a17332 = ~a17330 & ~a12072;
assign a17334 = a10300 & a10286;
assign a17336 = ~a17334 & a12072;
assign a17338 = ~a17336 & ~a17332;
assign a17340 = ~a17338 & a12058;
assign a17342 = ~a17340 & ~a17310;
assign a17344 = a15926 & a15910;
assign a17346 = ~a17344 & a12374;
assign a17348 = a17346 & ~a12372;
assign a17350 = a15630 & a15614;
assign a17352 = ~a17350 & a12372;
assign a17354 = ~a17352 & ~a17348;
assign a17356 = ~a17354 & ~a12370;
assign a17358 = a15334 & a15318;
assign a17360 = ~a17358 & a12370;
assign a17362 = ~a17360 & ~a17356;
assign a17364 = ~a17362 & ~a12368;
assign a17366 = a15038 & a15022;
assign a17368 = ~a17366 & a12368;
assign a17370 = ~a17368 & ~a17364;
assign a17372 = ~a17370 & a12366;
assign a17374 = a17372 & ~a12364;
assign a17376 = a14742 & a14726;
assign a17378 = ~a17376 & a12374;
assign a17380 = a17378 & ~a12372;
assign a17382 = a14446 & a14430;
assign a17384 = ~a17382 & a12372;
assign a17386 = ~a17384 & ~a17380;
assign a17388 = ~a17386 & ~a12370;
assign a17390 = a14150 & a14134;
assign a17392 = ~a17390 & a12370;
assign a17394 = ~a17392 & ~a17388;
assign a17396 = ~a17394 & ~a12368;
assign a17398 = a13854 & a13838;
assign a17400 = ~a17398 & a12368;
assign a17402 = ~a17400 & ~a17396;
assign a17404 = ~a17402 & a12364;
assign a17406 = ~a17404 & ~a17374;
assign a17408 = ~a17406 & ~a12362;
assign a17410 = a13558 & a13542;
assign a17412 = ~a17410 & a12374;
assign a17414 = a17412 & ~a12372;
assign a17416 = a13262 & a13246;
assign a17418 = ~a17416 & a12372;
assign a17420 = ~a17418 & ~a17414;
assign a17422 = ~a17420 & ~a12370;
assign a17424 = a12966 & a12950;
assign a17426 = ~a17424 & a12370;
assign a17428 = ~a17426 & ~a17422;
assign a17430 = ~a17428 & ~a12368;
assign a17432 = a12670 & a12654;
assign a17434 = ~a17432 & a12368;
assign a17436 = ~a17434 & ~a17430;
assign a17438 = ~a17436 & a12362;
assign a17440 = ~a17438 & ~a17408;
assign a17442 = ~a17440 & ~a12358;
assign a17444 = a12374 & ~a12358;
assign a17446 = a17444 & ~a12372;
assign a17448 = a12078 & a12062;
assign a17450 = ~a17448 & a12372;
assign a17452 = ~a17450 & ~a17446;
assign a17454 = ~a17452 & ~a12370;
assign a17456 = a11782 & a11766;
assign a17458 = ~a17456 & a12370;
assign a17460 = ~a17458 & ~a17454;
assign a17462 = ~a17460 & ~a12368;
assign a17464 = a11486 & a11470;
assign a17466 = ~a17464 & a12368;
assign a17468 = ~a17466 & ~a17462;
assign a17470 = ~a17468 & a12358;
assign a17472 = ~a17470 & ~a17442;
assign a17474 = ~a17472 & ~a12354;
assign a17476 = a11190 & a11174;
assign a17478 = ~a17476 & a12374;
assign a17480 = a17478 & ~a12372;
assign a17482 = a10894 & a10878;
assign a17484 = ~a17482 & a12372;
assign a17486 = ~a17484 & ~a17480;
assign a17488 = ~a17486 & ~a12370;
assign a17490 = a10598 & a10582;
assign a17492 = ~a17490 & a12370;
assign a17494 = ~a17492 & ~a17488;
assign a17496 = ~a17494 & ~a12368;
assign a17498 = a10302 & a10286;
assign a17500 = ~a17498 & a12368;
assign a17502 = ~a17500 & ~a17496;
assign a17504 = ~a17502 & a12354;
assign a17506 = ~a17504 & ~a17474;
assign a17508 = a15920 & a15914;
assign a17510 = ~a17508 & a12670;
assign a17512 = a17510 & ~a12668;
assign a17514 = a15624 & a15618;
assign a17516 = ~a17514 & a12668;
assign a17518 = ~a17516 & ~a17512;
assign a17520 = ~a17518 & ~a12666;
assign a17522 = a15328 & a15322;
assign a17524 = ~a17522 & a12666;
assign a17526 = ~a17524 & ~a17520;
assign a17528 = ~a17526 & ~a12664;
assign a17530 = a15032 & a15026;
assign a17532 = ~a17530 & a12664;
assign a17534 = ~a17532 & ~a17528;
assign a17536 = ~a17534 & a12662;
assign a17538 = a17536 & ~a12660;
assign a17540 = a14736 & a14730;
assign a17542 = ~a17540 & a12670;
assign a17544 = a17542 & ~a12668;
assign a17546 = a14440 & a14434;
assign a17548 = ~a17546 & a12668;
assign a17550 = ~a17548 & ~a17544;
assign a17552 = ~a17550 & ~a12666;
assign a17554 = a14144 & a14138;
assign a17556 = ~a17554 & a12666;
assign a17558 = ~a17556 & ~a17552;
assign a17560 = ~a17558 & ~a12664;
assign a17562 = a13848 & a13842;
assign a17564 = ~a17562 & a12664;
assign a17566 = ~a17564 & ~a17560;
assign a17568 = ~a17566 & a12660;
assign a17570 = ~a17568 & ~a17538;
assign a17572 = ~a17570 & ~a12658;
assign a17574 = a13552 & a13546;
assign a17576 = ~a17574 & a12670;
assign a17578 = a17576 & ~a12668;
assign a17580 = a13256 & a13250;
assign a17582 = ~a17580 & a12668;
assign a17584 = ~a17582 & ~a17578;
assign a17586 = ~a17584 & ~a12666;
assign a17588 = a12960 & a12954;
assign a17590 = ~a17588 & a12666;
assign a17592 = ~a17590 & ~a17586;
assign a17594 = ~a17592 & ~a12664;
assign a17596 = a12664 & ~a12658;
assign a17598 = ~a17596 & ~a17594;
assign a17600 = ~a17598 & a12658;
assign a17602 = ~a17600 & ~a17572;
assign a17604 = ~a17602 & ~a12654;
assign a17606 = a12368 & a12362;
assign a17608 = ~a17606 & a12670;
assign a17610 = a17608 & ~a12668;
assign a17612 = a12072 & a12066;
assign a17614 = ~a17612 & a12668;
assign a17616 = ~a17614 & ~a17610;
assign a17618 = ~a17616 & ~a12666;
assign a17620 = a11776 & a11770;
assign a17622 = ~a17620 & a12666;
assign a17624 = ~a17622 & ~a17618;
assign a17626 = ~a17624 & ~a12664;
assign a17628 = a11480 & a11474;
assign a17630 = ~a17628 & a12664;
assign a17632 = ~a17630 & ~a17626;
assign a17634 = ~a17632 & a12654;
assign a17636 = ~a17634 & ~a17604;
assign a17638 = ~a17636 & ~a12650;
assign a17640 = a11184 & a11178;
assign a17642 = ~a17640 & a12670;
assign a17644 = a17642 & ~a12668;
assign a17646 = a10888 & a10882;
assign a17648 = ~a17646 & a12668;
assign a17650 = ~a17648 & ~a17644;
assign a17652 = ~a17650 & ~a12666;
assign a17654 = a10592 & a10586;
assign a17656 = ~a17654 & a12666;
assign a17658 = ~a17656 & ~a17652;
assign a17660 = ~a17658 & ~a12664;
assign a17662 = a10296 & a10290;
assign a17664 = ~a17662 & a12664;
assign a17666 = ~a17664 & ~a17660;
assign a17668 = ~a17666 & a12650;
assign a17670 = ~a17668 & ~a17638;
assign a17672 = a15922 & a15914;
assign a17674 = ~a17672 & a12966;
assign a17676 = a17674 & ~a12964;
assign a17678 = a15626 & a15618;
assign a17680 = ~a17678 & a12964;
assign a17682 = ~a17680 & ~a17676;
assign a17684 = ~a17682 & ~a12962;
assign a17686 = a15330 & a15322;
assign a17688 = ~a17686 & a12962;
assign a17690 = ~a17688 & ~a17684;
assign a17692 = ~a17690 & ~a12960;
assign a17694 = a15034 & a15026;
assign a17696 = ~a17694 & a12960;
assign a17698 = ~a17696 & ~a17692;
assign a17700 = ~a17698 & a12958;
assign a17702 = a17700 & ~a12956;
assign a17704 = a14738 & a14730;
assign a17706 = ~a17704 & a12966;
assign a17708 = a17706 & ~a12964;
assign a17710 = a14442 & a14434;
assign a17712 = ~a17710 & a12964;
assign a17714 = ~a17712 & ~a17708;
assign a17716 = ~a17714 & ~a12962;
assign a17718 = a14146 & a14138;
assign a17720 = ~a17718 & a12962;
assign a17722 = ~a17720 & ~a17716;
assign a17724 = ~a17722 & ~a12960;
assign a17726 = a13850 & a13842;
assign a17728 = ~a17726 & a12960;
assign a17730 = ~a17728 & ~a17724;
assign a17732 = ~a17730 & a12956;
assign a17734 = ~a17732 & ~a17702;
assign a17736 = ~a17734 & ~a12954;
assign a17738 = a13554 & a13546;
assign a17740 = ~a17738 & a12966;
assign a17742 = a17740 & ~a12964;
assign a17744 = a13258 & a13250;
assign a17746 = ~a17744 & a12964;
assign a17748 = ~a17746 & ~a17742;
assign a17750 = ~a17748 & ~a12962;
assign a17752 = a12962 & ~a12954;
assign a17754 = ~a17752 & ~a17750;
assign a17756 = ~a17754 & ~a12960;
assign a17758 = a12666 & a12658;
assign a17760 = ~a17758 & a12960;
assign a17762 = ~a17760 & ~a17756;
assign a17764 = ~a17762 & a12954;
assign a17766 = ~a17764 & ~a17736;
assign a17768 = ~a17766 & ~a12950;
assign a17770 = a12370 & a12362;
assign a17772 = ~a17770 & a12966;
assign a17774 = a17772 & ~a12964;
assign a17776 = a12074 & a12066;
assign a17778 = ~a17776 & a12964;
assign a17780 = ~a17778 & ~a17774;
assign a17782 = ~a17780 & ~a12962;
assign a17784 = a11778 & a11770;
assign a17786 = ~a17784 & a12962;
assign a17788 = ~a17786 & ~a17782;
assign a17790 = ~a17788 & ~a12960;
assign a17792 = a11482 & a11474;
assign a17794 = ~a17792 & a12960;
assign a17796 = ~a17794 & ~a17790;
assign a17798 = ~a17796 & a12950;
assign a17800 = ~a17798 & ~a17768;
assign a17802 = ~a17800 & ~a12946;
assign a17804 = a11186 & a11178;
assign a17806 = ~a17804 & a12966;
assign a17808 = a17806 & ~a12964;
assign a17810 = a10890 & a10882;
assign a17812 = ~a17810 & a12964;
assign a17814 = ~a17812 & ~a17808;
assign a17816 = ~a17814 & ~a12962;
assign a17818 = a10594 & a10586;
assign a17820 = ~a17818 & a12962;
assign a17822 = ~a17820 & ~a17816;
assign a17824 = ~a17822 & ~a12960;
assign a17826 = a10298 & a10290;
assign a17828 = ~a17826 & a12960;
assign a17830 = ~a17828 & ~a17824;
assign a17832 = ~a17830 & a12946;
assign a17834 = ~a17832 & ~a17802;
assign a17836 = a15924 & a15914;
assign a17838 = ~a17836 & a13262;
assign a17840 = a17838 & ~a13260;
assign a17842 = a15628 & a15618;
assign a17844 = ~a17842 & a13260;
assign a17846 = ~a17844 & ~a17840;
assign a17848 = ~a17846 & ~a13258;
assign a17850 = a15332 & a15322;
assign a17852 = ~a17850 & a13258;
assign a17854 = ~a17852 & ~a17848;
assign a17856 = ~a17854 & ~a13256;
assign a17858 = a15036 & a15026;
assign a17860 = ~a17858 & a13256;
assign a17862 = ~a17860 & ~a17856;
assign a17864 = ~a17862 & a13254;
assign a17866 = a17864 & ~a13252;
assign a17868 = a14740 & a14730;
assign a17870 = ~a17868 & a13262;
assign a17872 = a17870 & ~a13260;
assign a17874 = a14444 & a14434;
assign a17876 = ~a17874 & a13260;
assign a17878 = ~a17876 & ~a17872;
assign a17880 = ~a17878 & ~a13258;
assign a17882 = a14148 & a14138;
assign a17884 = ~a17882 & a13258;
assign a17886 = ~a17884 & ~a17880;
assign a17888 = ~a17886 & ~a13256;
assign a17890 = a13852 & a13842;
assign a17892 = ~a17890 & a13256;
assign a17894 = ~a17892 & ~a17888;
assign a17896 = ~a17894 & a13252;
assign a17898 = ~a17896 & ~a17866;
assign a17900 = ~a17898 & ~a13250;
assign a17902 = a13556 & a13546;
assign a17904 = ~a17902 & a13262;
assign a17906 = a17904 & ~a13260;
assign a17908 = a13260 & ~a13250;
assign a17910 = ~a17908 & ~a17906;
assign a17912 = ~a17910 & ~a13258;
assign a17914 = a12964 & a12954;
assign a17916 = ~a17914 & a13258;
assign a17918 = ~a17916 & ~a17912;
assign a17920 = ~a17918 & ~a13256;
assign a17922 = a12668 & a12658;
assign a17924 = ~a17922 & a13256;
assign a17926 = ~a17924 & ~a17920;
assign a17928 = ~a17926 & a13250;
assign a17930 = ~a17928 & ~a17900;
assign a17932 = ~a17930 & ~a13246;
assign a17934 = a12372 & a12362;
assign a17936 = ~a17934 & a13262;
assign a17938 = a17936 & ~a13260;
assign a17940 = a12076 & a12066;
assign a17942 = ~a17940 & a13260;
assign a17944 = ~a17942 & ~a17938;
assign a17946 = ~a17944 & ~a13258;
assign a17948 = a11780 & a11770;
assign a17950 = ~a17948 & a13258;
assign a17952 = ~a17950 & ~a17946;
assign a17954 = ~a17952 & ~a13256;
assign a17956 = a11484 & a11474;
assign a17958 = ~a17956 & a13256;
assign a17960 = ~a17958 & ~a17954;
assign a17962 = ~a17960 & a13246;
assign a17964 = ~a17962 & ~a17932;
assign a17966 = ~a17964 & ~a13242;
assign a17968 = a11188 & a11178;
assign a17970 = ~a17968 & a13262;
assign a17972 = a17970 & ~a13260;
assign a17974 = a10892 & a10882;
assign a17976 = ~a17974 & a13260;
assign a17978 = ~a17976 & ~a17972;
assign a17980 = ~a17978 & ~a13258;
assign a17982 = a10596 & a10586;
assign a17984 = ~a17982 & a13258;
assign a17986 = ~a17984 & ~a17980;
assign a17988 = ~a17986 & ~a13256;
assign a17990 = a10300 & a10290;
assign a17992 = ~a17990 & a13256;
assign a17994 = ~a17992 & ~a17988;
assign a17996 = ~a17994 & a13242;
assign a17998 = ~a17996 & ~a17966;
assign a18000 = a15926 & a15914;
assign a18002 = ~a18000 & a13558;
assign a18004 = a18002 & ~a13556;
assign a18006 = a15630 & a15618;
assign a18008 = ~a18006 & a13556;
assign a18010 = ~a18008 & ~a18004;
assign a18012 = ~a18010 & ~a13554;
assign a18014 = a15334 & a15322;
assign a18016 = ~a18014 & a13554;
assign a18018 = ~a18016 & ~a18012;
assign a18020 = ~a18018 & ~a13552;
assign a18022 = a15038 & a15026;
assign a18024 = ~a18022 & a13552;
assign a18026 = ~a18024 & ~a18020;
assign a18028 = ~a18026 & a13550;
assign a18030 = a18028 & ~a13548;
assign a18032 = a14742 & a14730;
assign a18034 = ~a18032 & a13558;
assign a18036 = a18034 & ~a13556;
assign a18038 = a14446 & a14434;
assign a18040 = ~a18038 & a13556;
assign a18042 = ~a18040 & ~a18036;
assign a18044 = ~a18042 & ~a13554;
assign a18046 = a14150 & a14138;
assign a18048 = ~a18046 & a13554;
assign a18050 = ~a18048 & ~a18044;
assign a18052 = ~a18050 & ~a13552;
assign a18054 = a13854 & a13842;
assign a18056 = ~a18054 & a13552;
assign a18058 = ~a18056 & ~a18052;
assign a18060 = ~a18058 & a13548;
assign a18062 = ~a18060 & ~a18030;
assign a18064 = ~a18062 & ~a13546;
assign a18066 = a13558 & ~a13546;
assign a18068 = a18066 & ~a13556;
assign a18070 = a13262 & a13250;
assign a18072 = ~a18070 & a13556;
assign a18074 = ~a18072 & ~a18068;
assign a18076 = ~a18074 & ~a13554;
assign a18078 = a12966 & a12954;
assign a18080 = ~a18078 & a13554;
assign a18082 = ~a18080 & ~a18076;
assign a18084 = ~a18082 & ~a13552;
assign a18086 = a12670 & a12658;
assign a18088 = ~a18086 & a13552;
assign a18090 = ~a18088 & ~a18084;
assign a18092 = ~a18090 & a13546;
assign a18094 = ~a18092 & ~a18064;
assign a18096 = ~a18094 & ~a13542;
assign a18098 = a12374 & a12362;
assign a18100 = ~a18098 & a13558;
assign a18102 = a18100 & ~a13556;
assign a18104 = a12078 & a12066;
assign a18106 = ~a18104 & a13556;
assign a18108 = ~a18106 & ~a18102;
assign a18110 = ~a18108 & ~a13554;
assign a18112 = a11782 & a11770;
assign a18114 = ~a18112 & a13554;
assign a18116 = ~a18114 & ~a18110;
assign a18118 = ~a18116 & ~a13552;
assign a18120 = a11486 & a11474;
assign a18122 = ~a18120 & a13552;
assign a18124 = ~a18122 & ~a18118;
assign a18126 = ~a18124 & a13542;
assign a18128 = ~a18126 & ~a18096;
assign a18130 = ~a18128 & ~a13538;
assign a18132 = a11190 & a11178;
assign a18134 = ~a18132 & a13558;
assign a18136 = a18134 & ~a13556;
assign a18138 = a10894 & a10882;
assign a18140 = ~a18138 & a13556;
assign a18142 = ~a18140 & ~a18136;
assign a18144 = ~a18142 & ~a13554;
assign a18146 = a10598 & a10586;
assign a18148 = ~a18146 & a13554;
assign a18150 = ~a18148 & ~a18144;
assign a18152 = ~a18150 & ~a13552;
assign a18154 = a10302 & a10290;
assign a18156 = ~a18154 & a13552;
assign a18158 = ~a18156 & ~a18152;
assign a18160 = ~a18158 & a13538;
assign a18162 = ~a18160 & ~a18130;
assign a18164 = a15920 & a15916;
assign a18166 = ~a18164 & a13854;
assign a18168 = a18166 & ~a13852;
assign a18170 = a15624 & a15620;
assign a18172 = ~a18170 & a13852;
assign a18174 = ~a18172 & ~a18168;
assign a18176 = ~a18174 & ~a13850;
assign a18178 = a15328 & a15324;
assign a18180 = ~a18178 & a13850;
assign a18182 = ~a18180 & ~a18176;
assign a18184 = ~a18182 & ~a13848;
assign a18186 = a15032 & a15028;
assign a18188 = ~a18186 & a13848;
assign a18190 = ~a18188 & ~a18184;
assign a18192 = ~a18190 & a13846;
assign a18194 = a18192 & ~a13844;
assign a18196 = a14736 & a14732;
assign a18198 = ~a18196 & a13854;
assign a18200 = a18198 & ~a13852;
assign a18202 = a14440 & a14436;
assign a18204 = ~a18202 & a13852;
assign a18206 = ~a18204 & ~a18200;
assign a18208 = ~a18206 & ~a13850;
assign a18210 = a14144 & a14140;
assign a18212 = ~a18210 & a13850;
assign a18214 = ~a18212 & ~a18208;
assign a18216 = ~a18214 & ~a13848;
assign a18218 = a13848 & ~a13844;
assign a18220 = ~a18218 & ~a18216;
assign a18222 = ~a18220 & a13844;
assign a18224 = ~a18222 & ~a18194;
assign a18226 = ~a18224 & ~a13842;
assign a18228 = a13552 & a13548;
assign a18230 = ~a18228 & a13854;
assign a18232 = a18230 & ~a13852;
assign a18234 = a13256 & a13252;
assign a18236 = ~a18234 & a13852;
assign a18238 = ~a18236 & ~a18232;
assign a18240 = ~a18238 & ~a13850;
assign a18242 = a12960 & a12956;
assign a18244 = ~a18242 & a13850;
assign a18246 = ~a18244 & ~a18240;
assign a18248 = ~a18246 & ~a13848;
assign a18250 = a12664 & a12660;
assign a18252 = ~a18250 & a13848;
assign a18254 = ~a18252 & ~a18248;
assign a18256 = ~a18254 & a13842;
assign a18258 = ~a18256 & ~a18226;
assign a18260 = ~a18258 & ~a13838;
assign a18262 = a12368 & a12364;
assign a18264 = ~a18262 & a13854;
assign a18266 = a18264 & ~a13852;
assign a18268 = a12072 & a12068;
assign a18270 = ~a18268 & a13852;
assign a18272 = ~a18270 & ~a18266;
assign a18274 = ~a18272 & ~a13850;
assign a18276 = a11776 & a11772;
assign a18278 = ~a18276 & a13850;
assign a18280 = ~a18278 & ~a18274;
assign a18282 = ~a18280 & ~a13848;
assign a18284 = a11480 & a11476;
assign a18286 = ~a18284 & a13848;
assign a18288 = ~a18286 & ~a18282;
assign a18290 = ~a18288 & a13838;
assign a18292 = ~a18290 & ~a18260;
assign a18294 = ~a18292 & ~a13834;
assign a18296 = a11184 & a11180;
assign a18298 = ~a18296 & a13854;
assign a18300 = a18298 & ~a13852;
assign a18302 = a10888 & a10884;
assign a18304 = ~a18302 & a13852;
assign a18306 = ~a18304 & ~a18300;
assign a18308 = ~a18306 & ~a13850;
assign a18310 = a10592 & a10588;
assign a18312 = ~a18310 & a13850;
assign a18314 = ~a18312 & ~a18308;
assign a18316 = ~a18314 & ~a13848;
assign a18318 = a10296 & a10292;
assign a18320 = ~a18318 & a13848;
assign a18322 = ~a18320 & ~a18316;
assign a18324 = ~a18322 & a13834;
assign a18326 = ~a18324 & ~a18294;
assign a18328 = a15922 & a15916;
assign a18330 = ~a18328 & a14150;
assign a18332 = a18330 & ~a14148;
assign a18334 = a15626 & a15620;
assign a18336 = ~a18334 & a14148;
assign a18338 = ~a18336 & ~a18332;
assign a18340 = ~a18338 & ~a14146;
assign a18342 = a15330 & a15324;
assign a18344 = ~a18342 & a14146;
assign a18346 = ~a18344 & ~a18340;
assign a18348 = ~a18346 & ~a14144;
assign a18350 = a15034 & a15028;
assign a18352 = ~a18350 & a14144;
assign a18354 = ~a18352 & ~a18348;
assign a18356 = ~a18354 & a14142;
assign a18358 = a18356 & ~a14140;
assign a18360 = a14738 & a14732;
assign a18362 = ~a18360 & a14150;
assign a18364 = a18362 & ~a14148;
assign a18366 = a14442 & a14436;
assign a18368 = ~a18366 & a14148;
assign a18370 = ~a18368 & ~a18364;
assign a18372 = ~a18370 & ~a14146;
assign a18374 = a14146 & ~a14140;
assign a18376 = ~a18374 & ~a18372;
assign a18378 = ~a18376 & ~a14144;
assign a18380 = a13850 & a13844;
assign a18382 = ~a18380 & a14144;
assign a18384 = ~a18382 & ~a18378;
assign a18386 = ~a18384 & a14140;
assign a18388 = ~a18386 & ~a18358;
assign a18390 = ~a18388 & ~a14138;
assign a18392 = a13554 & a13548;
assign a18394 = ~a18392 & a14150;
assign a18396 = a18394 & ~a14148;
assign a18398 = a13258 & a13252;
assign a18400 = ~a18398 & a14148;
assign a18402 = ~a18400 & ~a18396;
assign a18404 = ~a18402 & ~a14146;
assign a18406 = a12962 & a12956;
assign a18408 = ~a18406 & a14146;
assign a18410 = ~a18408 & ~a18404;
assign a18412 = ~a18410 & ~a14144;
assign a18414 = a12666 & a12660;
assign a18416 = ~a18414 & a14144;
assign a18418 = ~a18416 & ~a18412;
assign a18420 = ~a18418 & a14138;
assign a18422 = ~a18420 & ~a18390;
assign a18424 = ~a18422 & ~a14134;
assign a18426 = a12370 & a12364;
assign a18428 = ~a18426 & a14150;
assign a18430 = a18428 & ~a14148;
assign a18432 = a12074 & a12068;
assign a18434 = ~a18432 & a14148;
assign a18436 = ~a18434 & ~a18430;
assign a18438 = ~a18436 & ~a14146;
assign a18440 = a11778 & a11772;
assign a18442 = ~a18440 & a14146;
assign a18444 = ~a18442 & ~a18438;
assign a18446 = ~a18444 & ~a14144;
assign a18448 = a11482 & a11476;
assign a18450 = ~a18448 & a14144;
assign a18452 = ~a18450 & ~a18446;
assign a18454 = ~a18452 & a14134;
assign a18456 = ~a18454 & ~a18424;
assign a18458 = ~a18456 & ~a14130;
assign a18460 = a11186 & a11180;
assign a18462 = ~a18460 & a14150;
assign a18464 = a18462 & ~a14148;
assign a18466 = a10890 & a10884;
assign a18468 = ~a18466 & a14148;
assign a18470 = ~a18468 & ~a18464;
assign a18472 = ~a18470 & ~a14146;
assign a18474 = a10594 & a10588;
assign a18476 = ~a18474 & a14146;
assign a18478 = ~a18476 & ~a18472;
assign a18480 = ~a18478 & ~a14144;
assign a18482 = a10298 & a10292;
assign a18484 = ~a18482 & a14144;
assign a18486 = ~a18484 & ~a18480;
assign a18488 = ~a18486 & a14130;
assign a18490 = ~a18488 & ~a18458;
assign a18492 = a15924 & a15916;
assign a18494 = ~a18492 & a14446;
assign a18496 = a18494 & ~a14444;
assign a18498 = a15628 & a15620;
assign a18500 = ~a18498 & a14444;
assign a18502 = ~a18500 & ~a18496;
assign a18504 = ~a18502 & ~a14442;
assign a18506 = a15332 & a15324;
assign a18508 = ~a18506 & a14442;
assign a18510 = ~a18508 & ~a18504;
assign a18512 = ~a18510 & ~a14440;
assign a18514 = a15036 & a15028;
assign a18516 = ~a18514 & a14440;
assign a18518 = ~a18516 & ~a18512;
assign a18520 = ~a18518 & a14438;
assign a18522 = a18520 & ~a14436;
assign a18524 = a14740 & a14732;
assign a18526 = ~a18524 & a14446;
assign a18528 = a18526 & ~a14444;
assign a18530 = a14444 & ~a14436;
assign a18532 = ~a18530 & ~a18528;
assign a18534 = ~a18532 & ~a14442;
assign a18536 = a14148 & a14140;
assign a18538 = ~a18536 & a14442;
assign a18540 = ~a18538 & ~a18534;
assign a18542 = ~a18540 & ~a14440;
assign a18544 = a13852 & a13844;
assign a18546 = ~a18544 & a14440;
assign a18548 = ~a18546 & ~a18542;
assign a18550 = ~a18548 & a14436;
assign a18552 = ~a18550 & ~a18522;
assign a18554 = ~a18552 & ~a14434;
assign a18556 = a13556 & a13548;
assign a18558 = ~a18556 & a14446;
assign a18560 = a18558 & ~a14444;
assign a18562 = a13260 & a13252;
assign a18564 = ~a18562 & a14444;
assign a18566 = ~a18564 & ~a18560;
assign a18568 = ~a18566 & ~a14442;
assign a18570 = a12964 & a12956;
assign a18572 = ~a18570 & a14442;
assign a18574 = ~a18572 & ~a18568;
assign a18576 = ~a18574 & ~a14440;
assign a18578 = a12668 & a12660;
assign a18580 = ~a18578 & a14440;
assign a18582 = ~a18580 & ~a18576;
assign a18584 = ~a18582 & a14434;
assign a18586 = ~a18584 & ~a18554;
assign a18588 = ~a18586 & ~a14430;
assign a18590 = a12372 & a12364;
assign a18592 = ~a18590 & a14446;
assign a18594 = a18592 & ~a14444;
assign a18596 = a12076 & a12068;
assign a18598 = ~a18596 & a14444;
assign a18600 = ~a18598 & ~a18594;
assign a18602 = ~a18600 & ~a14442;
assign a18604 = a11780 & a11772;
assign a18606 = ~a18604 & a14442;
assign a18608 = ~a18606 & ~a18602;
assign a18610 = ~a18608 & ~a14440;
assign a18612 = a11484 & a11476;
assign a18614 = ~a18612 & a14440;
assign a18616 = ~a18614 & ~a18610;
assign a18618 = ~a18616 & a14430;
assign a18620 = ~a18618 & ~a18588;
assign a18622 = ~a18620 & ~a14426;
assign a18624 = a11188 & a11180;
assign a18626 = ~a18624 & a14446;
assign a18628 = a18626 & ~a14444;
assign a18630 = a10892 & a10884;
assign a18632 = ~a18630 & a14444;
assign a18634 = ~a18632 & ~a18628;
assign a18636 = ~a18634 & ~a14442;
assign a18638 = a10596 & a10588;
assign a18640 = ~a18638 & a14442;
assign a18642 = ~a18640 & ~a18636;
assign a18644 = ~a18642 & ~a14440;
assign a18646 = a10300 & a10292;
assign a18648 = ~a18646 & a14440;
assign a18650 = ~a18648 & ~a18644;
assign a18652 = ~a18650 & a14426;
assign a18654 = ~a18652 & ~a18622;
assign a18656 = a15926 & a15916;
assign a18658 = ~a18656 & a14742;
assign a18660 = a18658 & ~a14740;
assign a18662 = a15630 & a15620;
assign a18664 = ~a18662 & a14740;
assign a18666 = ~a18664 & ~a18660;
assign a18668 = ~a18666 & ~a14738;
assign a18670 = a15334 & a15324;
assign a18672 = ~a18670 & a14738;
assign a18674 = ~a18672 & ~a18668;
assign a18676 = ~a18674 & ~a14736;
assign a18678 = a15038 & a15028;
assign a18680 = ~a18678 & a14736;
assign a18682 = ~a18680 & ~a18676;
assign a18684 = ~a18682 & a14734;
assign a18686 = a18684 & ~a14732;
assign a18688 = a14742 & ~a14732;
assign a18690 = a18688 & ~a14740;
assign a18692 = a14446 & a14436;
assign a18694 = ~a18692 & a14740;
assign a18696 = ~a18694 & ~a18690;
assign a18698 = ~a18696 & ~a14738;
assign a18700 = a14150 & a14140;
assign a18702 = ~a18700 & a14738;
assign a18704 = ~a18702 & ~a18698;
assign a18706 = ~a18704 & ~a14736;
assign a18708 = a13854 & a13844;
assign a18710 = ~a18708 & a14736;
assign a18712 = ~a18710 & ~a18706;
assign a18714 = ~a18712 & a14732;
assign a18716 = ~a18714 & ~a18686;
assign a18718 = ~a18716 & ~a14730;
assign a18720 = a13558 & a13548;
assign a18722 = ~a18720 & a14742;
assign a18724 = a18722 & ~a14740;
assign a18726 = a13262 & a13252;
assign a18728 = ~a18726 & a14740;
assign a18730 = ~a18728 & ~a18724;
assign a18732 = ~a18730 & ~a14738;
assign a18734 = a12966 & a12956;
assign a18736 = ~a18734 & a14738;
assign a18738 = ~a18736 & ~a18732;
assign a18740 = ~a18738 & ~a14736;
assign a18742 = a12670 & a12660;
assign a18744 = ~a18742 & a14736;
assign a18746 = ~a18744 & ~a18740;
assign a18748 = ~a18746 & a14730;
assign a18750 = ~a18748 & ~a18718;
assign a18752 = ~a18750 & ~a14726;
assign a18754 = a12374 & a12364;
assign a18756 = ~a18754 & a14742;
assign a18758 = a18756 & ~a14740;
assign a18760 = a12078 & a12068;
assign a18762 = ~a18760 & a14740;
assign a18764 = ~a18762 & ~a18758;
assign a18766 = ~a18764 & ~a14738;
assign a18768 = a11782 & a11772;
assign a18770 = ~a18768 & a14738;
assign a18772 = ~a18770 & ~a18766;
assign a18774 = ~a18772 & ~a14736;
assign a18776 = a11486 & a11476;
assign a18778 = ~a18776 & a14736;
assign a18780 = ~a18778 & ~a18774;
assign a18782 = ~a18780 & a14726;
assign a18784 = ~a18782 & ~a18752;
assign a18786 = ~a18784 & ~a14722;
assign a18788 = a11190 & a11180;
assign a18790 = ~a18788 & a14742;
assign a18792 = a18790 & ~a14740;
assign a18794 = a10894 & a10884;
assign a18796 = ~a18794 & a14740;
assign a18798 = ~a18796 & ~a18792;
assign a18800 = ~a18798 & ~a14738;
assign a18802 = a10598 & a10588;
assign a18804 = ~a18802 & a14738;
assign a18806 = ~a18804 & ~a18800;
assign a18808 = ~a18806 & ~a14736;
assign a18810 = a10302 & a10292;
assign a18812 = ~a18810 & a14736;
assign a18814 = ~a18812 & ~a18808;
assign a18816 = ~a18814 & a14722;
assign a18818 = ~a18816 & ~a18786;
assign a18820 = a15920 & a15918;
assign a18822 = ~a18820 & a15038;
assign a18824 = a18822 & ~a15036;
assign a18826 = a15624 & a15622;
assign a18828 = ~a18826 & a15036;
assign a18830 = ~a18828 & ~a18824;
assign a18832 = ~a18830 & ~a15034;
assign a18834 = a15328 & a15326;
assign a18836 = ~a18834 & a15034;
assign a18838 = ~a18836 & ~a18832;
assign a18840 = ~a18838 & ~a15032;
assign a18842 = a15032 & ~a15030;
assign a18844 = ~a18842 & ~a18840;
assign a18846 = ~a18844 & a15030;
assign a18848 = a18846 & ~a15028;
assign a18850 = a14736 & a14734;
assign a18852 = ~a18850 & a15038;
assign a18854 = a18852 & ~a15036;
assign a18856 = a14440 & a14438;
assign a18858 = ~a18856 & a15036;
assign a18860 = ~a18858 & ~a18854;
assign a18862 = ~a18860 & ~a15034;
assign a18864 = a14144 & a14142;
assign a18866 = ~a18864 & a15034;
assign a18868 = ~a18866 & ~a18862;
assign a18870 = ~a18868 & ~a15032;
assign a18872 = a13848 & a13846;
assign a18874 = ~a18872 & a15032;
assign a18876 = ~a18874 & ~a18870;
assign a18878 = ~a18876 & a15028;
assign a18880 = ~a18878 & ~a18848;
assign a18882 = ~a18880 & ~a15026;
assign a18884 = a13552 & a13550;
assign a18886 = ~a18884 & a15038;
assign a18888 = a18886 & ~a15036;
assign a18890 = a13256 & a13254;
assign a18892 = ~a18890 & a15036;
assign a18894 = ~a18892 & ~a18888;
assign a18896 = ~a18894 & ~a15034;
assign a18898 = a12960 & a12958;
assign a18900 = ~a18898 & a15034;
assign a18902 = ~a18900 & ~a18896;
assign a18904 = ~a18902 & ~a15032;
assign a18906 = a12664 & a12662;
assign a18908 = ~a18906 & a15032;
assign a18910 = ~a18908 & ~a18904;
assign a18912 = ~a18910 & a15026;
assign a18914 = ~a18912 & ~a18882;
assign a18916 = ~a18914 & ~a15022;
assign a18918 = a12368 & a12366;
assign a18920 = ~a18918 & a15038;
assign a18922 = a18920 & ~a15036;
assign a18924 = a12072 & a12070;
assign a18926 = ~a18924 & a15036;
assign a18928 = ~a18926 & ~a18922;
assign a18930 = ~a18928 & ~a15034;
assign a18932 = a11776 & a11774;
assign a18934 = ~a18932 & a15034;
assign a18936 = ~a18934 & ~a18930;
assign a18938 = ~a18936 & ~a15032;
assign a18940 = a11480 & a11478;
assign a18942 = ~a18940 & a15032;
assign a18944 = ~a18942 & ~a18938;
assign a18946 = ~a18944 & a15022;
assign a18948 = ~a18946 & ~a18916;
assign a18950 = ~a18948 & ~a15018;
assign a18952 = a11184 & a11182;
assign a18954 = ~a18952 & a15038;
assign a18956 = a18954 & ~a15036;
assign a18958 = a10888 & a10886;
assign a18960 = ~a18958 & a15036;
assign a18962 = ~a18960 & ~a18956;
assign a18964 = ~a18962 & ~a15034;
assign a18966 = a10592 & a10590;
assign a18968 = ~a18966 & a15034;
assign a18970 = ~a18968 & ~a18964;
assign a18972 = ~a18970 & ~a15032;
assign a18974 = a10296 & a10294;
assign a18976 = ~a18974 & a15032;
assign a18978 = ~a18976 & ~a18972;
assign a18980 = ~a18978 & a15018;
assign a18982 = ~a18980 & ~a18950;
assign a18984 = a15922 & a15918;
assign a18986 = ~a18984 & a15334;
assign a18988 = a18986 & ~a15332;
assign a18990 = a15626 & a15622;
assign a18992 = ~a18990 & a15332;
assign a18994 = ~a18992 & ~a18988;
assign a18996 = ~a18994 & ~a15330;
assign a18998 = a15330 & ~a15326;
assign a19000 = ~a18998 & ~a18996;
assign a19002 = ~a19000 & ~a15328;
assign a19004 = a15034 & a15030;
assign a19006 = ~a19004 & a15328;
assign a19008 = ~a19006 & ~a19002;
assign a19010 = ~a19008 & a15326;
assign a19012 = a19010 & ~a15324;
assign a19014 = a14738 & a14734;
assign a19016 = ~a19014 & a15334;
assign a19018 = a19016 & ~a15332;
assign a19020 = a14442 & a14438;
assign a19022 = ~a19020 & a15332;
assign a19024 = ~a19022 & ~a19018;
assign a19026 = ~a19024 & ~a15330;
assign a19028 = a14146 & a14142;
assign a19030 = ~a19028 & a15330;
assign a19032 = ~a19030 & ~a19026;
assign a19034 = ~a19032 & ~a15328;
assign a19036 = a13850 & a13846;
assign a19038 = ~a19036 & a15328;
assign a19040 = ~a19038 & ~a19034;
assign a19042 = ~a19040 & a15324;
assign a19044 = ~a19042 & ~a19012;
assign a19046 = ~a19044 & ~a15322;
assign a19048 = a13554 & a13550;
assign a19050 = ~a19048 & a15334;
assign a19052 = a19050 & ~a15332;
assign a19054 = a13258 & a13254;
assign a19056 = ~a19054 & a15332;
assign a19058 = ~a19056 & ~a19052;
assign a19060 = ~a19058 & ~a15330;
assign a19062 = a12962 & a12958;
assign a19064 = ~a19062 & a15330;
assign a19066 = ~a19064 & ~a19060;
assign a19068 = ~a19066 & ~a15328;
assign a19070 = a12666 & a12662;
assign a19072 = ~a19070 & a15328;
assign a19074 = ~a19072 & ~a19068;
assign a19076 = ~a19074 & a15322;
assign a19078 = ~a19076 & ~a19046;
assign a19080 = ~a19078 & ~a15318;
assign a19082 = a12370 & a12366;
assign a19084 = ~a19082 & a15334;
assign a19086 = a19084 & ~a15332;
assign a19088 = a12074 & a12070;
assign a19090 = ~a19088 & a15332;
assign a19092 = ~a19090 & ~a19086;
assign a19094 = ~a19092 & ~a15330;
assign a19096 = a11778 & a11774;
assign a19098 = ~a19096 & a15330;
assign a19100 = ~a19098 & ~a19094;
assign a19102 = ~a19100 & ~a15328;
assign a19104 = a11482 & a11478;
assign a19106 = ~a19104 & a15328;
assign a19108 = ~a19106 & ~a19102;
assign a19110 = ~a19108 & a15318;
assign a19112 = ~a19110 & ~a19080;
assign a19114 = ~a19112 & ~a15314;
assign a19116 = a11186 & a11182;
assign a19118 = ~a19116 & a15334;
assign a19120 = a19118 & ~a15332;
assign a19122 = a10890 & a10886;
assign a19124 = ~a19122 & a15332;
assign a19126 = ~a19124 & ~a19120;
assign a19128 = ~a19126 & ~a15330;
assign a19130 = a10594 & a10590;
assign a19132 = ~a19130 & a15330;
assign a19134 = ~a19132 & ~a19128;
assign a19136 = ~a19134 & ~a15328;
assign a19138 = a10298 & a10294;
assign a19140 = ~a19138 & a15328;
assign a19142 = ~a19140 & ~a19136;
assign a19144 = ~a19142 & a15314;
assign a19146 = ~a19144 & ~a19114;
assign a19148 = a15924 & a15918;
assign a19150 = ~a19148 & a15630;
assign a19152 = a19150 & ~a15628;
assign a19154 = a15628 & ~a15622;
assign a19156 = ~a19154 & ~a19152;
assign a19158 = ~a19156 & ~a15626;
assign a19160 = a15332 & a15326;
assign a19162 = ~a19160 & a15626;
assign a19164 = ~a19162 & ~a19158;
assign a19166 = ~a19164 & ~a15624;
assign a19168 = a15036 & a15030;
assign a19170 = ~a19168 & a15624;
assign a19172 = ~a19170 & ~a19166;
assign a19174 = ~a19172 & a15622;
assign a19176 = a19174 & ~a15620;
assign a19178 = a14740 & a14734;
assign a19180 = ~a19178 & a15630;
assign a19182 = a19180 & ~a15628;
assign a19184 = a14444 & a14438;
assign a19186 = ~a19184 & a15628;
assign a19188 = ~a19186 & ~a19182;
assign a19190 = ~a19188 & ~a15626;
assign a19192 = a14148 & a14142;
assign a19194 = ~a19192 & a15626;
assign a19196 = ~a19194 & ~a19190;
assign a19198 = ~a19196 & ~a15624;
assign a19200 = a13852 & a13846;
assign a19202 = ~a19200 & a15624;
assign a19204 = ~a19202 & ~a19198;
assign a19206 = ~a19204 & a15620;
assign a19208 = ~a19206 & ~a19176;
assign a19210 = ~a19208 & ~a15618;
assign a19212 = a13556 & a13550;
assign a19214 = ~a19212 & a15630;
assign a19216 = a19214 & ~a15628;
assign a19218 = a13260 & a13254;
assign a19220 = ~a19218 & a15628;
assign a19222 = ~a19220 & ~a19216;
assign a19224 = ~a19222 & ~a15626;
assign a19226 = a12964 & a12958;
assign a19228 = ~a19226 & a15626;
assign a19230 = ~a19228 & ~a19224;
assign a19232 = ~a19230 & ~a15624;
assign a19234 = a12668 & a12662;
assign a19236 = ~a19234 & a15624;
assign a19238 = ~a19236 & ~a19232;
assign a19240 = ~a19238 & a15618;
assign a19242 = ~a19240 & ~a19210;
assign a19244 = ~a19242 & ~a15614;
assign a19246 = a12372 & a12366;
assign a19248 = ~a19246 & a15630;
assign a19250 = a19248 & ~a15628;
assign a19252 = a12076 & a12070;
assign a19254 = ~a19252 & a15628;
assign a19256 = ~a19254 & ~a19250;
assign a19258 = ~a19256 & ~a15626;
assign a19260 = a11780 & a11774;
assign a19262 = ~a19260 & a15626;
assign a19264 = ~a19262 & ~a19258;
assign a19266 = ~a19264 & ~a15624;
assign a19268 = a11484 & a11478;
assign a19270 = ~a19268 & a15624;
assign a19272 = ~a19270 & ~a19266;
assign a19274 = ~a19272 & a15614;
assign a19276 = ~a19274 & ~a19244;
assign a19278 = ~a19276 & ~a15610;
assign a19280 = a11188 & a11182;
assign a19282 = ~a19280 & a15630;
assign a19284 = a19282 & ~a15628;
assign a19286 = a10892 & a10886;
assign a19288 = ~a19286 & a15628;
assign a19290 = ~a19288 & ~a19284;
assign a19292 = ~a19290 & ~a15626;
assign a19294 = a10596 & a10590;
assign a19296 = ~a19294 & a15626;
assign a19298 = ~a19296 & ~a19292;
assign a19300 = ~a19298 & ~a15624;
assign a19302 = a10300 & a10294;
assign a19304 = ~a19302 & a15624;
assign a19306 = ~a19304 & ~a19300;
assign a19308 = ~a19306 & a15610;
assign a19310 = ~a19308 & ~a19278;
assign a19312 = a15926 & ~a15918;
assign a19314 = a19312 & ~a15924;
assign a19316 = a15630 & a15622;
assign a19318 = ~a19316 & a15924;
assign a19320 = ~a19318 & ~a19314;
assign a19322 = ~a19320 & ~a15922;
assign a19324 = a15334 & a15326;
assign a19326 = ~a19324 & a15922;
assign a19328 = ~a19326 & ~a19322;
assign a19330 = ~a19328 & ~a15920;
assign a19332 = a15038 & a15030;
assign a19334 = ~a19332 & a15920;
assign a19336 = ~a19334 & ~a19330;
assign a19338 = ~a19336 & a15918;
assign a19340 = a19338 & ~a15916;
assign a19342 = a14742 & a14734;
assign a19344 = ~a19342 & a15926;
assign a19346 = a19344 & ~a15924;
assign a19348 = a14446 & a14438;
assign a19350 = ~a19348 & a15924;
assign a19352 = ~a19350 & ~a19346;
assign a19354 = ~a19352 & ~a15922;
assign a19356 = a14150 & a14142;
assign a19358 = ~a19356 & a15922;
assign a19360 = ~a19358 & ~a19354;
assign a19362 = ~a19360 & ~a15920;
assign a19364 = a13854 & a13846;
assign a19366 = ~a19364 & a15920;
assign a19368 = ~a19366 & ~a19362;
assign a19370 = ~a19368 & a15916;
assign a19372 = ~a19370 & ~a19340;
assign a19374 = ~a19372 & ~a15914;
assign a19376 = a13558 & a13550;
assign a19378 = ~a19376 & a15926;
assign a19380 = a19378 & ~a15924;
assign a19382 = a13262 & a13254;
assign a19384 = ~a19382 & a15924;
assign a19386 = ~a19384 & ~a19380;
assign a19388 = ~a19386 & ~a15922;
assign a19390 = a12966 & a12958;
assign a19392 = ~a19390 & a15922;
assign a19394 = ~a19392 & ~a19388;
assign a19396 = ~a19394 & ~a15920;
assign a19398 = a12670 & a12662;
assign a19400 = ~a19398 & a15920;
assign a19402 = ~a19400 & ~a19396;
assign a19404 = ~a19402 & a15914;
assign a19406 = ~a19404 & ~a19374;
assign a19408 = ~a19406 & ~a15910;
assign a19410 = a12374 & a12366;
assign a19412 = ~a19410 & a15926;
assign a19414 = a19412 & ~a15924;
assign a19416 = a12078 & a12070;
assign a19418 = ~a19416 & a15924;
assign a19420 = ~a19418 & ~a19414;
assign a19422 = ~a19420 & ~a15922;
assign a19424 = a11782 & a11774;
assign a19426 = ~a19424 & a15922;
assign a19428 = ~a19426 & ~a19422;
assign a19430 = ~a19428 & ~a15920;
assign a19432 = a11486 & a11478;
assign a19434 = ~a19432 & a15920;
assign a19436 = ~a19434 & ~a19430;
assign a19438 = ~a19436 & a15910;
assign a19440 = ~a19438 & ~a19408;
assign a19442 = ~a19440 & ~a15906;
assign a19444 = a11190 & a11182;
assign a19446 = ~a19444 & a15926;
assign a19448 = a19446 & ~a15924;
assign a19450 = a10894 & a10886;
assign a19452 = ~a19450 & a15924;
assign a19454 = ~a19452 & ~a19448;
assign a19456 = ~a19454 & ~a15922;
assign a19458 = a10598 & a10590;
assign a19460 = ~a19458 & a15922;
assign a19462 = ~a19460 & ~a19456;
assign a19464 = ~a19462 & ~a15920;
assign a19466 = a10302 & a10294;
assign a19468 = ~a19466 & a15920;
assign a19470 = ~a19468 & ~a19464;
assign a19472 = ~a19470 & a15906;
assign a19474 = ~a19472 & ~a19442;
assign a19476 = ~a11480 & a11466;
assign a19478 = ~a11776 & a11762;
assign a19480 = ~a19478 & ~a19476;
assign a19482 = ~a12072 & a12058;
assign a19484 = ~a19482 & a19480;
assign a19486 = ~a12368 & a12354;
assign a19488 = ~a19486 & a19484;
assign a19490 = ~a12664 & a12650;
assign a19492 = ~a11770 & ~a11474;
assign a19494 = a19492 & ~a12066;
assign a19496 = a19494 & ~a12362;
assign a19498 = ~a11772 & ~a11476;
assign a19500 = a19498 & ~a12068;
assign a19502 = a19500 & ~a12364;
assign a19504 = ~a14138 & ~a13842;
assign a19506 = a19504 & ~a14434;
assign a19508 = a19506 & ~a14730;
assign a19510 = ~a19508 & ~a19502;
assign a19512 = ~a11774 & ~a11478;
assign a19514 = a19512 & ~a12070;
assign a19516 = a19514 & ~a12366;
assign a19518 = ~a15322 & ~a15026;
assign a19520 = a19518 & ~a15618;
assign a19522 = a19520 & ~a15914;
assign a19524 = ~a19522 & ~a19516;
assign a19526 = ~a19524 & ~a19510;
assign a19528 = a19526 & a19496;
assign a19530 = ~a14142 & ~a13846;
assign a19532 = a19530 & ~a14438;
assign a19534 = a19532 & ~a14734;
assign a19536 = ~a19534 & ~a19522;
assign a19538 = a19536 & ~a19502;
assign a19540 = ~a15324 & ~a15028;
assign a19542 = a19540 & ~a15620;
assign a19544 = a19542 & ~a15916;
assign a19546 = ~a19544 & ~a19508;
assign a19548 = a19546 & ~a19516;
assign a19550 = ~a19548 & ~a19538;
assign a19552 = a19550 & a19528;
assign a19554 = ~a19552 & a19490;
assign a19556 = ~a12960 & a12946;
assign a19558 = a19556 & ~a19552;
assign a19560 = ~a13256 & a13242;
assign a19562 = a19560 & ~a19552;
assign a19564 = ~a13552 & a13538;
assign a19566 = a19564 & ~a19552;
assign a19568 = ~a13848 & a13834;
assign a19570 = ~a12956 & ~a12660;
assign a19572 = a19570 & ~a13252;
assign a19574 = a19572 & ~a13548;
assign a19576 = ~a19574 & ~a19496;
assign a19578 = ~a19544 & ~a19516;
assign a19580 = ~a19578 & ~a19576;
assign a19582 = a19580 & a19502;
assign a19584 = ~a12958 & ~a12662;
assign a19586 = a19584 & ~a13254;
assign a19588 = a19586 & ~a13550;
assign a19590 = ~a19588 & ~a19544;
assign a19592 = a19590 & ~a19496;
assign a19594 = ~a19574 & ~a19522;
assign a19596 = a19594 & ~a19516;
assign a19598 = ~a19596 & ~a19592;
assign a19600 = a19598 & a19582;
assign a19602 = ~a19600 & a19568;
assign a19604 = ~a14144 & a14130;
assign a19606 = a19604 & ~a19600;
assign a19608 = ~a14440 & a14426;
assign a19610 = a19608 & ~a19600;
assign a19612 = ~a14736 & a14722;
assign a19614 = a19612 & ~a19600;
assign a19616 = ~a15032 & a15018;
assign a19618 = ~a19588 & ~a19496;
assign a19620 = ~a19534 & ~a19502;
assign a19622 = ~a19620 & ~a19618;
assign a19624 = a19622 & a19516;
assign a19626 = ~a19574 & ~a19534;
assign a19628 = a19626 & ~a19496;
assign a19630 = ~a19588 & ~a19508;
assign a19632 = a19630 & ~a19502;
assign a19634 = ~a19632 & ~a19628;
assign a19636 = a19634 & a19624;
assign a19638 = ~a19636 & a19616;
assign a19640 = ~a15328 & a15314;
assign a19642 = a19640 & ~a19636;
assign a19644 = ~a15624 & a15610;
assign a19646 = a19644 & ~a19636;
assign a19648 = ~a15920 & a15906;
assign a19650 = a19648 & ~a19636;
assign a19652 = ~a19650 & ~a19646;
assign a19654 = a19652 & ~a19642;
assign a19656 = a19654 & ~a19638;
assign a19658 = a19656 & ~a19614;
assign a19660 = a19658 & ~a19610;
assign a19662 = a19660 & ~a19606;
assign a19664 = a19662 & ~a19602;
assign a19666 = a19664 & ~a19566;
assign a19668 = a19666 & ~a19562;
assign a19670 = a19668 & ~a19558;
assign a19672 = a19670 & ~a19554;
assign a19674 = a19672 & a19488;
assign a19676 = ~a19674 & a10286;
assign a19678 = ~a11482 & a11466;
assign a19680 = ~a11778 & a11762;
assign a19682 = ~a19680 & ~a19678;
assign a19684 = ~a12074 & a12058;
assign a19686 = ~a19684 & a19682;
assign a19688 = ~a12370 & a12354;
assign a19690 = ~a19688 & a19686;
assign a19692 = ~a12666 & a12650;
assign a19694 = a19692 & ~a19552;
assign a19696 = ~a12962 & a12946;
assign a19698 = a19696 & ~a19552;
assign a19700 = ~a13258 & a13242;
assign a19702 = a19700 & ~a19552;
assign a19704 = ~a13554 & a13538;
assign a19706 = a19704 & ~a19552;
assign a19708 = ~a13850 & a13834;
assign a19710 = a19708 & ~a19600;
assign a19712 = ~a14146 & a14130;
assign a19714 = a19712 & ~a19600;
assign a19716 = ~a14442 & a14426;
assign a19718 = a19716 & ~a19600;
assign a19720 = ~a14738 & a14722;
assign a19722 = a19720 & ~a19600;
assign a19724 = ~a15034 & a15018;
assign a19726 = a19724 & ~a19636;
assign a19728 = ~a15330 & a15314;
assign a19730 = a19728 & ~a19636;
assign a19732 = ~a15626 & a15610;
assign a19734 = a19732 & ~a19636;
assign a19736 = ~a15922 & a15906;
assign a19738 = a19736 & ~a19636;
assign a19740 = ~a19738 & ~a19734;
assign a19742 = a19740 & ~a19730;
assign a19744 = a19742 & ~a19726;
assign a19746 = a19744 & ~a19722;
assign a19748 = a19746 & ~a19718;
assign a19750 = a19748 & ~a19714;
assign a19752 = a19750 & ~a19710;
assign a19754 = a19752 & ~a19706;
assign a19756 = a19754 & ~a19702;
assign a19758 = a19756 & ~a19698;
assign a19760 = a19758 & ~a19694;
assign a19762 = a19760 & a19690;
assign a19764 = ~a19762 & a10582;
assign a19766 = ~a11484 & a11466;
assign a19768 = ~a11780 & a11762;
assign a19770 = ~a19768 & ~a19766;
assign a19772 = ~a12076 & a12058;
assign a19774 = ~a19772 & a19770;
assign a19776 = ~a12372 & a12354;
assign a19778 = ~a19776 & a19774;
assign a19780 = ~a12668 & a12650;
assign a19782 = a19780 & ~a19552;
assign a19784 = ~a12964 & a12946;
assign a19786 = a19784 & ~a19552;
assign a19788 = ~a13260 & a13242;
assign a19790 = a19788 & ~a19552;
assign a19792 = ~a13556 & a13538;
assign a19794 = a19792 & ~a19552;
assign a19796 = ~a13852 & a13834;
assign a19798 = a19796 & ~a19600;
assign a19800 = ~a14148 & a14130;
assign a19802 = a19800 & ~a19600;
assign a19804 = ~a14444 & a14426;
assign a19806 = a19804 & ~a19600;
assign a19808 = ~a14740 & a14722;
assign a19810 = a19808 & ~a19600;
assign a19812 = ~a15036 & a15018;
assign a19814 = a19812 & ~a19636;
assign a19816 = ~a15332 & a15314;
assign a19818 = a19816 & ~a19636;
assign a19820 = ~a15628 & a15610;
assign a19822 = a19820 & ~a19636;
assign a19824 = ~a15924 & a15906;
assign a19826 = a19824 & ~a19636;
assign a19828 = ~a19826 & ~a19822;
assign a19830 = a19828 & ~a19818;
assign a19832 = a19830 & ~a19814;
assign a19834 = a19832 & ~a19810;
assign a19836 = a19834 & ~a19806;
assign a19838 = a19836 & ~a19802;
assign a19840 = a19838 & ~a19798;
assign a19842 = a19840 & ~a19794;
assign a19844 = a19842 & ~a19790;
assign a19846 = a19844 & ~a19786;
assign a19848 = a19846 & ~a19782;
assign a19850 = a19848 & a19778;
assign a19852 = ~a19850 & a10878;
assign a19854 = ~a11486 & a11466;
assign a19856 = ~a11782 & a11762;
assign a19858 = ~a19856 & ~a19854;
assign a19860 = ~a12078 & a12058;
assign a19862 = ~a19860 & a19858;
assign a19864 = ~a12374 & a12354;
assign a19866 = ~a19864 & a19862;
assign a19868 = ~a12670 & a12650;
assign a19870 = a19868 & ~a19552;
assign a19872 = ~a12966 & a12946;
assign a19874 = a19872 & ~a19552;
assign a19876 = ~a13262 & a13242;
assign a19878 = a19876 & ~a19552;
assign a19880 = ~a13558 & a13538;
assign a19882 = a19880 & ~a19552;
assign a19884 = ~a13854 & a13834;
assign a19886 = a19884 & ~a19600;
assign a19888 = ~a14150 & a14130;
assign a19890 = a19888 & ~a19600;
assign a19892 = ~a14446 & a14426;
assign a19894 = a19892 & ~a19600;
assign a19896 = ~a14742 & a14722;
assign a19898 = a19896 & ~a19600;
assign a19900 = ~a15038 & a15018;
assign a19902 = a19900 & ~a19636;
assign a19904 = ~a15334 & a15314;
assign a19906 = a19904 & ~a19636;
assign a19908 = ~a15630 & a15610;
assign a19910 = a19908 & ~a19636;
assign a19912 = ~a15926 & a15906;
assign a19914 = a19912 & ~a19636;
assign a19916 = ~a19914 & ~a19910;
assign a19918 = a19916 & ~a19906;
assign a19920 = a19918 & ~a19902;
assign a19922 = a19920 & ~a19898;
assign a19924 = a19922 & ~a19894;
assign a19926 = a19924 & ~a19890;
assign a19928 = a19926 & ~a19886;
assign a19930 = a19928 & ~a19882;
assign a19932 = a19930 & ~a19878;
assign a19934 = a19932 & ~a19874;
assign a19936 = a19934 & ~a19870;
assign a19938 = a19936 & a19866;
assign a19940 = ~a19938 & a11174;
assign a19942 = ~a12950 & ~a12654;
assign a19944 = a19942 & ~a13246;
assign a19946 = a19944 & ~a13542;
assign a19948 = ~a14134 & ~a13838;
assign a19950 = a19948 & ~a14430;
assign a19952 = a19950 & ~a14726;
assign a19954 = ~a19952 & ~a19574;
assign a19956 = ~a15318 & ~a15022;
assign a19958 = a19956 & ~a15614;
assign a19960 = a19958 & ~a15910;
assign a19962 = ~a19960 & ~a19588;
assign a19964 = ~a19962 & ~a19954;
assign a19966 = a19964 & a19946;
assign a19968 = ~a19960 & ~a19534;
assign a19970 = a19968 & ~a19574;
assign a19972 = ~a19952 & ~a19544;
assign a19974 = a19972 & ~a19588;
assign a19976 = ~a19974 & ~a19970;
assign a19978 = a19976 & a19966;
assign a19980 = ~a19978 & ~a19488;
assign a19982 = ~a19946 & ~a19502;
assign a19984 = ~a19982 & ~a19590;
assign a19986 = a19984 & a19574;
assign a19988 = ~a19946 & a19578;
assign a19990 = ~a19960 & ~a19502;
assign a19992 = a19990 & ~a19588;
assign a19994 = ~a19992 & ~a19988;
assign a19996 = a19994 & a19986;
assign a19998 = ~a19996 & a19568;
assign a20000 = ~a19996 & a19604;
assign a20002 = ~a19996 & a19608;
assign a20004 = ~a19996 & a19612;
assign a20006 = ~a19946 & ~a19516;
assign a20008 = ~a20006 & ~a19626;
assign a20010 = a20008 & a19588;
assign a20012 = ~a19946 & a19620;
assign a20014 = ~a19952 & ~a19516;
assign a20016 = a20014 & ~a19574;
assign a20018 = ~a20016 & ~a20012;
assign a20020 = a20018 & a20010;
assign a20022 = ~a20020 & a19616;
assign a20024 = ~a20020 & a19640;
assign a20026 = ~a20020 & a19644;
assign a20028 = ~a20020 & a19648;
assign a20030 = ~a20028 & ~a20026;
assign a20032 = a20030 & ~a20024;
assign a20034 = a20032 & ~a20022;
assign a20036 = a20034 & ~a20004;
assign a20038 = a20036 & ~a20002;
assign a20040 = a20038 & ~a20000;
assign a20042 = a20040 & ~a19998;
assign a20044 = a20042 & ~a19980;
assign a20046 = a20044 & ~a19490;
assign a20048 = a20046 & ~a19556;
assign a20050 = a20048 & ~a19560;
assign a20052 = a20050 & ~a19564;
assign a20054 = ~a20052 & a10290;
assign a20056 = ~a19978 & ~a19690;
assign a20058 = ~a19996 & a19708;
assign a20060 = ~a19996 & a19712;
assign a20062 = ~a19996 & a19716;
assign a20064 = ~a19996 & a19720;
assign a20066 = ~a20020 & a19724;
assign a20068 = ~a20020 & a19728;
assign a20070 = ~a20020 & a19732;
assign a20072 = ~a20020 & a19736;
assign a20074 = ~a20072 & ~a20070;
assign a20076 = a20074 & ~a20068;
assign a20078 = a20076 & ~a20066;
assign a20080 = a20078 & ~a20064;
assign a20082 = a20080 & ~a20062;
assign a20084 = a20082 & ~a20060;
assign a20086 = a20084 & ~a20058;
assign a20088 = a20086 & ~a20056;
assign a20090 = a20088 & ~a19692;
assign a20092 = a20090 & ~a19696;
assign a20094 = a20092 & ~a19700;
assign a20096 = a20094 & ~a19704;
assign a20098 = ~a20096 & a10586;
assign a20100 = ~a19978 & ~a19778;
assign a20102 = ~a19996 & a19796;
assign a20104 = ~a19996 & a19800;
assign a20106 = ~a19996 & a19804;
assign a20108 = ~a19996 & a19808;
assign a20110 = ~a20020 & a19812;
assign a20112 = ~a20020 & a19816;
assign a20114 = ~a20020 & a19820;
assign a20116 = ~a20020 & a19824;
assign a20118 = ~a20116 & ~a20114;
assign a20120 = a20118 & ~a20112;
assign a20122 = a20120 & ~a20110;
assign a20124 = a20122 & ~a20108;
assign a20126 = a20124 & ~a20106;
assign a20128 = a20126 & ~a20104;
assign a20130 = a20128 & ~a20102;
assign a20132 = a20130 & ~a20100;
assign a20134 = a20132 & ~a19780;
assign a20136 = a20134 & ~a19784;
assign a20138 = a20136 & ~a19788;
assign a20140 = a20138 & ~a19792;
assign a20142 = ~a20140 & a10882;
assign a20144 = ~a19978 & ~a19866;
assign a20146 = ~a19996 & a19884;
assign a20148 = ~a19996 & a19888;
assign a20150 = ~a19996 & a19892;
assign a20152 = ~a19996 & a19896;
assign a20154 = ~a20020 & a19900;
assign a20156 = ~a20020 & a19904;
assign a20158 = ~a20020 & a19908;
assign a20160 = ~a20020 & a19912;
assign a20162 = ~a20160 & ~a20158;
assign a20164 = a20162 & ~a20156;
assign a20166 = a20164 & ~a20154;
assign a20168 = a20166 & ~a20152;
assign a20170 = a20168 & ~a20150;
assign a20172 = a20170 & ~a20148;
assign a20174 = a20172 & ~a20146;
assign a20176 = a20174 & ~a20144;
assign a20178 = a20176 & ~a19868;
assign a20180 = a20178 & ~a19872;
assign a20182 = a20180 & ~a19876;
assign a20184 = a20182 & ~a19880;
assign a20186 = ~a20184 & a11178;
assign a20188 = ~a19946 & ~a19508;
assign a20190 = ~a20188 & ~a19968;
assign a20192 = a20190 & a19952;
assign a20194 = a19962 & ~a19508;
assign a20196 = ~a19946 & ~a19522;
assign a20198 = a20196 & ~a19534;
assign a20200 = ~a20198 & ~a20194;
assign a20202 = a20200 & a20192;
assign a20204 = ~a20202 & ~a19488;
assign a20206 = ~a19952 & ~a19496;
assign a20208 = ~a20206 & ~a19536;
assign a20210 = a20208 & a19508;
assign a20212 = ~a19952 & a19524;
assign a20214 = ~a19960 & ~a19496;
assign a20216 = a20214 & ~a19534;
assign a20218 = ~a20216 & ~a20212;
assign a20220 = a20218 & a20210;
assign a20222 = ~a20220 & a19490;
assign a20224 = ~a20220 & a19556;
assign a20226 = ~a20220 & a19560;
assign a20228 = ~a20220 & a19564;
assign a20230 = ~a20014 & ~a19630;
assign a20232 = a20230 & a19534;
assign a20234 = ~a19952 & a19618;
assign a20236 = a20006 & ~a19508;
assign a20238 = ~a20236 & ~a20234;
assign a20240 = a20238 & a20232;
assign a20242 = ~a20240 & a19616;
assign a20244 = ~a20240 & a19640;
assign a20246 = ~a20240 & a19644;
assign a20248 = ~a20240 & a19648;
assign a20250 = ~a20248 & ~a20246;
assign a20252 = a20250 & ~a20244;
assign a20254 = a20252 & ~a20242;
assign a20256 = a20254 & ~a20228;
assign a20258 = a20256 & ~a20226;
assign a20260 = a20258 & ~a20224;
assign a20262 = a20260 & ~a20222;
assign a20264 = a20262 & ~a20204;
assign a20266 = a20264 & ~a19568;
assign a20268 = a20266 & ~a19604;
assign a20270 = a20268 & ~a19608;
assign a20272 = a20270 & ~a19612;
assign a20274 = ~a20272 & a10292;
assign a20276 = ~a20202 & ~a19690;
assign a20278 = ~a20220 & a19692;
assign a20280 = ~a20220 & a19696;
assign a20282 = ~a20220 & a19700;
assign a20284 = ~a20220 & a19704;
assign a20286 = ~a20240 & a19724;
assign a20288 = ~a20240 & a19728;
assign a20290 = ~a20240 & a19732;
assign a20292 = ~a20240 & a19736;
assign a20294 = ~a20292 & ~a20290;
assign a20296 = a20294 & ~a20288;
assign a20298 = a20296 & ~a20286;
assign a20300 = a20298 & ~a20284;
assign a20302 = a20300 & ~a20282;
assign a20304 = a20302 & ~a20280;
assign a20306 = a20304 & ~a20278;
assign a20308 = a20306 & ~a20276;
assign a20310 = a20308 & ~a19708;
assign a20312 = a20310 & ~a19712;
assign a20314 = a20312 & ~a19716;
assign a20316 = a20314 & ~a19720;
assign a20318 = ~a20316 & a10588;
assign a20320 = ~a20202 & ~a19778;
assign a20322 = ~a20220 & a19780;
assign a20324 = ~a20220 & a19784;
assign a20326 = ~a20220 & a19788;
assign a20328 = ~a20220 & a19792;
assign a20330 = ~a20240 & a19812;
assign a20332 = ~a20240 & a19816;
assign a20334 = ~a20240 & a19820;
assign a20336 = ~a20240 & a19824;
assign a20338 = ~a20336 & ~a20334;
assign a20340 = a20338 & ~a20332;
assign a20342 = a20340 & ~a20330;
assign a20344 = a20342 & ~a20328;
assign a20346 = a20344 & ~a20326;
assign a20348 = a20346 & ~a20324;
assign a20350 = a20348 & ~a20322;
assign a20352 = a20350 & ~a20320;
assign a20354 = a20352 & ~a19796;
assign a20356 = a20354 & ~a19800;
assign a20358 = a20356 & ~a19804;
assign a20360 = a20358 & ~a19808;
assign a20362 = ~a20360 & a10884;
assign a20364 = ~a20202 & ~a19866;
assign a20366 = ~a20220 & a19868;
assign a20368 = ~a20220 & a19872;
assign a20370 = ~a20220 & a19876;
assign a20372 = ~a20220 & a19880;
assign a20374 = ~a20240 & a19900;
assign a20376 = ~a20240 & a19904;
assign a20378 = ~a20240 & a19908;
assign a20380 = ~a20240 & a19912;
assign a20382 = ~a20380 & ~a20378;
assign a20384 = a20382 & ~a20376;
assign a20386 = a20384 & ~a20374;
assign a20388 = a20386 & ~a20372;
assign a20390 = a20388 & ~a20370;
assign a20392 = a20390 & ~a20368;
assign a20394 = a20392 & ~a20366;
assign a20396 = a20394 & ~a20364;
assign a20398 = a20396 & ~a19884;
assign a20400 = a20398 & ~a19888;
assign a20402 = a20400 & ~a19892;
assign a20404 = a20402 & ~a19896;
assign a20406 = ~a20404 & a11180;
assign a20408 = ~a20196 & ~a19972;
assign a20410 = a20408 & a19960;
assign a20412 = a19954 & ~a19522;
assign a20414 = a20188 & ~a19544;
assign a20416 = ~a20414 & ~a20412;
assign a20418 = a20416 & a20410;
assign a20420 = ~a20418 & ~a19488;
assign a20422 = ~a20214 & ~a19546;
assign a20424 = a20422 & a19522;
assign a20426 = ~a19960 & a19510;
assign a20428 = a20206 & ~a19544;
assign a20430 = ~a20428 & ~a20426;
assign a20432 = a20430 & a20424;
assign a20434 = ~a20432 & a19490;
assign a20436 = ~a20432 & a19556;
assign a20438 = ~a20432 & a19560;
assign a20440 = ~a20432 & a19564;
assign a20442 = ~a19990 & ~a19594;
assign a20444 = a20442 & a19544;
assign a20446 = ~a19960 & a19576;
assign a20448 = a19982 & ~a19522;
assign a20450 = ~a20448 & ~a20446;
assign a20452 = a20450 & a20444;
assign a20454 = ~a20452 & a19568;
assign a20456 = ~a20452 & a19604;
assign a20458 = ~a20452 & a19608;
assign a20460 = ~a20452 & a19612;
assign a20462 = ~a20460 & ~a20458;
assign a20464 = a20462 & ~a20456;
assign a20466 = a20464 & ~a20454;
assign a20468 = a20466 & ~a20440;
assign a20470 = a20468 & ~a20438;
assign a20472 = a20470 & ~a20436;
assign a20474 = a20472 & ~a20434;
assign a20476 = a20474 & ~a20420;
assign a20478 = a20476 & ~a19616;
assign a20480 = a20478 & ~a19640;
assign a20482 = a20480 & ~a19644;
assign a20484 = a20482 & ~a19648;
assign a20486 = ~a20484 & a10294;
assign a20488 = ~a20418 & ~a19690;
assign a20490 = ~a20432 & a19692;
assign a20492 = ~a20432 & a19696;
assign a20494 = ~a20432 & a19700;
assign a20496 = ~a20432 & a19704;
assign a20498 = ~a20452 & a19708;
assign a20500 = ~a20452 & a19712;
assign a20502 = ~a20452 & a19716;
assign a20504 = ~a20452 & a19720;
assign a20506 = ~a20504 & ~a20502;
assign a20508 = a20506 & ~a20500;
assign a20510 = a20508 & ~a20498;
assign a20512 = a20510 & ~a20496;
assign a20514 = a20512 & ~a20494;
assign a20516 = a20514 & ~a20492;
assign a20518 = a20516 & ~a20490;
assign a20520 = a20518 & ~a20488;
assign a20522 = a20520 & ~a19724;
assign a20524 = a20522 & ~a19728;
assign a20526 = a20524 & ~a19732;
assign a20528 = a20526 & ~a19736;
assign a20530 = ~a20528 & a10590;
assign a20532 = ~a20418 & ~a19778;
assign a20534 = ~a20432 & a19780;
assign a20536 = ~a20432 & a19784;
assign a20538 = ~a20432 & a19788;
assign a20540 = ~a20432 & a19792;
assign a20542 = ~a20452 & a19796;
assign a20544 = ~a20452 & a19800;
assign a20546 = ~a20452 & a19804;
assign a20548 = ~a20452 & a19808;
assign a20550 = ~a20548 & ~a20546;
assign a20552 = a20550 & ~a20544;
assign a20554 = a20552 & ~a20542;
assign a20556 = a20554 & ~a20540;
assign a20558 = a20556 & ~a20538;
assign a20560 = a20558 & ~a20536;
assign a20562 = a20560 & ~a20534;
assign a20564 = a20562 & ~a20532;
assign a20566 = a20564 & ~a19812;
assign a20568 = a20566 & ~a19816;
assign a20570 = a20568 & ~a19820;
assign a20572 = a20570 & ~a19824;
assign a20574 = ~a20572 & a10886;
assign a20576 = ~a20418 & ~a19866;
assign a20578 = ~a20432 & a19868;
assign a20580 = ~a20432 & a19872;
assign a20582 = ~a20432 & a19876;
assign a20584 = ~a20432 & a19880;
assign a20586 = ~a20452 & a19884;
assign a20588 = ~a20452 & a19888;
assign a20590 = ~a20452 & a19892;
assign a20592 = ~a20452 & a19896;
assign a20594 = ~a20592 & ~a20590;
assign a20596 = a20594 & ~a20588;
assign a20598 = a20596 & ~a20586;
assign a20600 = a20598 & ~a20584;
assign a20602 = a20600 & ~a20582;
assign a20604 = a20602 & ~a20580;
assign a20606 = a20604 & ~a20578;
assign a20608 = a20606 & ~a20576;
assign a20610 = a20608 & ~a19900;
assign a20612 = a20610 & ~a19904;
assign a20614 = a20612 & ~a19908;
assign a20616 = a20614 & ~a19912;
assign a20618 = ~a20616 & a11182;
assign a20620 = ~a10296 & a10286;
assign a20622 = ~a10592 & a10582;
assign a20624 = ~a20622 & ~a20620;
assign a20626 = ~a10888 & a10878;
assign a20628 = ~a20626 & a20624;
assign a20630 = ~a11184 & a11174;
assign a20632 = ~a20630 & a20628;
assign a20634 = ~a12664 & a12654;
assign a20636 = ~a10586 & ~a10290;
assign a20638 = a20636 & ~a10882;
assign a20640 = a20638 & ~a11178;
assign a20642 = ~a10588 & ~a10292;
assign a20644 = a20642 & ~a10884;
assign a20646 = a20644 & ~a11180;
assign a20648 = ~a20646 & ~a19508;
assign a20650 = ~a10590 & ~a10294;
assign a20652 = a20650 & ~a10886;
assign a20654 = a20652 & ~a11182;
assign a20656 = ~a20654 & ~a19522;
assign a20658 = ~a20656 & ~a20648;
assign a20660 = a20658 & a20640;
assign a20662 = ~a20646 & a19536;
assign a20664 = ~a20654 & a19546;
assign a20666 = ~a20664 & ~a20662;
assign a20668 = a20666 & a20660;
assign a20670 = ~a20668 & a20634;
assign a20672 = ~a12960 & a12950;
assign a20674 = a20672 & ~a20668;
assign a20676 = ~a13256 & a13246;
assign a20678 = a20676 & ~a20668;
assign a20680 = ~a13552 & a13542;
assign a20682 = a20680 & ~a20668;
assign a20684 = ~a13848 & a13838;
assign a20686 = ~a20640 & ~a19574;
assign a20688 = ~a20654 & ~a19544;
assign a20690 = ~a20688 & ~a20686;
assign a20692 = a20690 & a20646;
assign a20694 = ~a20640 & a19590;
assign a20696 = ~a20654 & a19594;
assign a20698 = ~a20696 & ~a20694;
assign a20700 = a20698 & a20692;
assign a20702 = ~a20700 & a20684;
assign a20704 = ~a14144 & a14134;
assign a20706 = a20704 & ~a20700;
assign a20708 = ~a14440 & a14430;
assign a20710 = a20708 & ~a20700;
assign a20712 = ~a14736 & a14726;
assign a20714 = a20712 & ~a20700;
assign a20716 = ~a15032 & a15022;
assign a20718 = ~a20640 & ~a19588;
assign a20720 = ~a20646 & ~a19534;
assign a20722 = ~a20720 & ~a20718;
assign a20724 = a20722 & a20654;
assign a20726 = ~a20640 & a19626;
assign a20728 = ~a20646 & a19630;
assign a20730 = ~a20728 & ~a20726;
assign a20732 = a20730 & a20724;
assign a20734 = ~a20732 & a20716;
assign a20736 = ~a15328 & a15318;
assign a20738 = a20736 & ~a20732;
assign a20740 = ~a15624 & a15614;
assign a20742 = a20740 & ~a20732;
assign a20744 = ~a15920 & a15910;
assign a20746 = a20744 & ~a20732;
assign a20748 = ~a20746 & ~a20742;
assign a20750 = a20748 & ~a20738;
assign a20752 = a20750 & ~a20734;
assign a20754 = a20752 & ~a20714;
assign a20756 = a20754 & ~a20710;
assign a20758 = a20756 & ~a20706;
assign a20760 = a20758 & ~a20702;
assign a20762 = a20760 & ~a20682;
assign a20764 = a20762 & ~a20678;
assign a20766 = a20764 & ~a20674;
assign a20768 = a20766 & ~a20670;
assign a20770 = a20768 & a20632;
assign a20772 = ~a20770 & a11466;
assign a20774 = ~a10298 & a10286;
assign a20776 = ~a10594 & a10582;
assign a20778 = ~a20776 & ~a20774;
assign a20780 = ~a10890 & a10878;
assign a20782 = ~a20780 & a20778;
assign a20784 = ~a11186 & a11174;
assign a20786 = ~a20784 & a20782;
assign a20788 = ~a12666 & a12654;
assign a20790 = a20788 & ~a20668;
assign a20792 = ~a12962 & a12950;
assign a20794 = a20792 & ~a20668;
assign a20796 = ~a13258 & a13246;
assign a20798 = a20796 & ~a20668;
assign a20800 = ~a13554 & a13542;
assign a20802 = a20800 & ~a20668;
assign a20804 = ~a13850 & a13838;
assign a20806 = a20804 & ~a20700;
assign a20808 = ~a14146 & a14134;
assign a20810 = a20808 & ~a20700;
assign a20812 = ~a14442 & a14430;
assign a20814 = a20812 & ~a20700;
assign a20816 = ~a14738 & a14726;
assign a20818 = a20816 & ~a20700;
assign a20820 = ~a15034 & a15022;
assign a20822 = a20820 & ~a20732;
assign a20824 = ~a15330 & a15318;
assign a20826 = a20824 & ~a20732;
assign a20828 = ~a15626 & a15614;
assign a20830 = a20828 & ~a20732;
assign a20832 = ~a15922 & a15910;
assign a20834 = a20832 & ~a20732;
assign a20836 = ~a20834 & ~a20830;
assign a20838 = a20836 & ~a20826;
assign a20840 = a20838 & ~a20822;
assign a20842 = a20840 & ~a20818;
assign a20844 = a20842 & ~a20814;
assign a20846 = a20844 & ~a20810;
assign a20848 = a20846 & ~a20806;
assign a20850 = a20848 & ~a20802;
assign a20852 = a20850 & ~a20798;
assign a20854 = a20852 & ~a20794;
assign a20856 = a20854 & ~a20790;
assign a20858 = a20856 & a20786;
assign a20860 = ~a20858 & a11762;
assign a20862 = ~a10300 & a10286;
assign a20864 = ~a10596 & a10582;
assign a20866 = ~a20864 & ~a20862;
assign a20868 = ~a10892 & a10878;
assign a20870 = ~a20868 & a20866;
assign a20872 = ~a11188 & a11174;
assign a20874 = ~a20872 & a20870;
assign a20876 = ~a12668 & a12654;
assign a20878 = a20876 & ~a20668;
assign a20880 = ~a12964 & a12950;
assign a20882 = a20880 & ~a20668;
assign a20884 = ~a13260 & a13246;
assign a20886 = a20884 & ~a20668;
assign a20888 = ~a13556 & a13542;
assign a20890 = a20888 & ~a20668;
assign a20892 = ~a13852 & a13838;
assign a20894 = a20892 & ~a20700;
assign a20896 = ~a14148 & a14134;
assign a20898 = a20896 & ~a20700;
assign a20900 = ~a14444 & a14430;
assign a20902 = a20900 & ~a20700;
assign a20904 = ~a14740 & a14726;
assign a20906 = a20904 & ~a20700;
assign a20908 = ~a15036 & a15022;
assign a20910 = a20908 & ~a20732;
assign a20912 = ~a15332 & a15318;
assign a20914 = a20912 & ~a20732;
assign a20916 = ~a15628 & a15614;
assign a20918 = a20916 & ~a20732;
assign a20920 = ~a15924 & a15910;
assign a20922 = a20920 & ~a20732;
assign a20924 = ~a20922 & ~a20918;
assign a20926 = a20924 & ~a20914;
assign a20928 = a20926 & ~a20910;
assign a20930 = a20928 & ~a20906;
assign a20932 = a20930 & ~a20902;
assign a20934 = a20932 & ~a20898;
assign a20936 = a20934 & ~a20894;
assign a20938 = a20936 & ~a20890;
assign a20940 = a20938 & ~a20886;
assign a20942 = a20940 & ~a20882;
assign a20944 = a20942 & ~a20878;
assign a20946 = a20944 & a20874;
assign a20948 = ~a20946 & a12058;
assign a20950 = ~a10302 & a10286;
assign a20952 = ~a10598 & a10582;
assign a20954 = ~a20952 & ~a20950;
assign a20956 = ~a10894 & a10878;
assign a20958 = ~a20956 & a20954;
assign a20960 = ~a11190 & a11174;
assign a20962 = ~a20960 & a20958;
assign a20964 = ~a12670 & a12654;
assign a20966 = a20964 & ~a20668;
assign a20968 = ~a12966 & a12950;
assign a20970 = a20968 & ~a20668;
assign a20972 = ~a13262 & a13246;
assign a20974 = a20972 & ~a20668;
assign a20976 = ~a13558 & a13542;
assign a20978 = a20976 & ~a20668;
assign a20980 = ~a13854 & a13838;
assign a20982 = a20980 & ~a20700;
assign a20984 = ~a14150 & a14134;
assign a20986 = a20984 & ~a20700;
assign a20988 = ~a14446 & a14430;
assign a20990 = a20988 & ~a20700;
assign a20992 = ~a14742 & a14726;
assign a20994 = a20992 & ~a20700;
assign a20996 = ~a15038 & a15022;
assign a20998 = a20996 & ~a20732;
assign a21000 = ~a15334 & a15318;
assign a21002 = a21000 & ~a20732;
assign a21004 = ~a15630 & a15614;
assign a21006 = a21004 & ~a20732;
assign a21008 = ~a15926 & a15910;
assign a21010 = a21008 & ~a20732;
assign a21012 = ~a21010 & ~a21006;
assign a21014 = a21012 & ~a21002;
assign a21016 = a21014 & ~a20998;
assign a21018 = a21016 & ~a20994;
assign a21020 = a21018 & ~a20990;
assign a21022 = a21020 & ~a20986;
assign a21024 = a21022 & ~a20982;
assign a21026 = a21024 & ~a20978;
assign a21028 = a21026 & ~a20974;
assign a21030 = a21028 & ~a20970;
assign a21032 = a21030 & ~a20966;
assign a21034 = a21032 & a20962;
assign a21036 = ~a21034 & a12354;
assign a21038 = ~a12946 & ~a12650;
assign a21040 = a21038 & ~a13242;
assign a21042 = a21040 & ~a13538;
assign a21044 = ~a14130 & ~a13834;
assign a21046 = a21044 & ~a14426;
assign a21048 = a21046 & ~a14722;
assign a21050 = ~a21048 & ~a19574;
assign a21052 = ~a15314 & ~a15018;
assign a21054 = a21052 & ~a15610;
assign a21056 = a21054 & ~a15906;
assign a21058 = ~a21056 & ~a19588;
assign a21060 = ~a21058 & ~a21050;
assign a21062 = a21060 & a21042;
assign a21064 = ~a21056 & ~a19534;
assign a21066 = a21064 & ~a19574;
assign a21068 = ~a21048 & ~a19544;
assign a21070 = a21068 & ~a19588;
assign a21072 = ~a21070 & ~a21066;
assign a21074 = a21072 & a21062;
assign a21076 = ~a21074 & ~a20632;
assign a21078 = ~a21042 & ~a20646;
assign a21080 = ~a21078 & ~a19590;
assign a21082 = a21080 & a19574;
assign a21084 = ~a21042 & a20688;
assign a21086 = ~a21056 & ~a20646;
assign a21088 = a21086 & ~a19588;
assign a21090 = ~a21088 & ~a21084;
assign a21092 = a21090 & a21082;
assign a21094 = ~a21092 & a20684;
assign a21096 = ~a21092 & a20704;
assign a21098 = ~a21092 & a20708;
assign a21100 = ~a21092 & a20712;
assign a21102 = ~a21042 & ~a20654;
assign a21104 = ~a21102 & ~a19626;
assign a21106 = a21104 & a19588;
assign a21108 = ~a21042 & a20720;
assign a21110 = ~a21048 & ~a20654;
assign a21112 = a21110 & ~a19574;
assign a21114 = ~a21112 & ~a21108;
assign a21116 = a21114 & a21106;
assign a21118 = ~a21116 & a20716;
assign a21120 = ~a21116 & a20736;
assign a21122 = ~a21116 & a20740;
assign a21124 = ~a21116 & a20744;
assign a21126 = ~a21124 & ~a21122;
assign a21128 = a21126 & ~a21120;
assign a21130 = a21128 & ~a21118;
assign a21132 = a21130 & ~a21100;
assign a21134 = a21132 & ~a21098;
assign a21136 = a21134 & ~a21096;
assign a21138 = a21136 & ~a21094;
assign a21140 = a21138 & ~a21076;
assign a21142 = a21140 & ~a20634;
assign a21144 = a21142 & ~a20672;
assign a21146 = a21144 & ~a20676;
assign a21148 = a21146 & ~a20680;
assign a21150 = ~a21148 & a11474;
assign a21152 = ~a21074 & ~a20786;
assign a21154 = ~a21092 & a20804;
assign a21156 = ~a21092 & a20808;
assign a21158 = ~a21092 & a20812;
assign a21160 = ~a21092 & a20816;
assign a21162 = ~a21116 & a20820;
assign a21164 = ~a21116 & a20824;
assign a21166 = ~a21116 & a20828;
assign a21168 = ~a21116 & a20832;
assign a21170 = ~a21168 & ~a21166;
assign a21172 = a21170 & ~a21164;
assign a21174 = a21172 & ~a21162;
assign a21176 = a21174 & ~a21160;
assign a21178 = a21176 & ~a21158;
assign a21180 = a21178 & ~a21156;
assign a21182 = a21180 & ~a21154;
assign a21184 = a21182 & ~a21152;
assign a21186 = a21184 & ~a20788;
assign a21188 = a21186 & ~a20792;
assign a21190 = a21188 & ~a20796;
assign a21192 = a21190 & ~a20800;
assign a21194 = ~a21192 & a11770;
assign a21196 = ~a21074 & ~a20874;
assign a21198 = ~a21092 & a20892;
assign a21200 = ~a21092 & a20896;
assign a21202 = ~a21092 & a20900;
assign a21204 = ~a21092 & a20904;
assign a21206 = ~a21116 & a20908;
assign a21208 = ~a21116 & a20912;
assign a21210 = ~a21116 & a20916;
assign a21212 = ~a21116 & a20920;
assign a21214 = ~a21212 & ~a21210;
assign a21216 = a21214 & ~a21208;
assign a21218 = a21216 & ~a21206;
assign a21220 = a21218 & ~a21204;
assign a21222 = a21220 & ~a21202;
assign a21224 = a21222 & ~a21200;
assign a21226 = a21224 & ~a21198;
assign a21228 = a21226 & ~a21196;
assign a21230 = a21228 & ~a20876;
assign a21232 = a21230 & ~a20880;
assign a21234 = a21232 & ~a20884;
assign a21236 = a21234 & ~a20888;
assign a21238 = ~a21236 & a12066;
assign a21240 = ~a21074 & ~a20962;
assign a21242 = ~a21092 & a20980;
assign a21244 = ~a21092 & a20984;
assign a21246 = ~a21092 & a20988;
assign a21248 = ~a21092 & a20992;
assign a21250 = ~a21116 & a20996;
assign a21252 = ~a21116 & a21000;
assign a21254 = ~a21116 & a21004;
assign a21256 = ~a21116 & a21008;
assign a21258 = ~a21256 & ~a21254;
assign a21260 = a21258 & ~a21252;
assign a21262 = a21260 & ~a21250;
assign a21264 = a21262 & ~a21248;
assign a21266 = a21264 & ~a21246;
assign a21268 = a21266 & ~a21244;
assign a21270 = a21268 & ~a21242;
assign a21272 = a21270 & ~a21240;
assign a21274 = a21272 & ~a20964;
assign a21276 = a21274 & ~a20968;
assign a21278 = a21276 & ~a20972;
assign a21280 = a21278 & ~a20976;
assign a21282 = ~a21280 & a12362;
assign a21284 = ~a21042 & ~a19508;
assign a21286 = ~a21284 & ~a21064;
assign a21288 = a21286 & a21048;
assign a21290 = a21058 & ~a19508;
assign a21292 = ~a21042 & ~a19522;
assign a21294 = a21292 & ~a19534;
assign a21296 = ~a21294 & ~a21290;
assign a21298 = a21296 & a21288;
assign a21300 = ~a21298 & ~a20632;
assign a21302 = ~a21048 & ~a20640;
assign a21304 = ~a21302 & ~a19536;
assign a21306 = a21304 & a19508;
assign a21308 = ~a21048 & a20656;
assign a21310 = ~a21056 & ~a20640;
assign a21312 = a21310 & ~a19534;
assign a21314 = ~a21312 & ~a21308;
assign a21316 = a21314 & a21306;
assign a21318 = ~a21316 & a20634;
assign a21320 = ~a21316 & a20672;
assign a21322 = ~a21316 & a20676;
assign a21324 = ~a21316 & a20680;
assign a21326 = ~a21110 & ~a19630;
assign a21328 = a21326 & a19534;
assign a21330 = ~a21048 & a20718;
assign a21332 = a21102 & ~a19508;
assign a21334 = ~a21332 & ~a21330;
assign a21336 = a21334 & a21328;
assign a21338 = ~a21336 & a20716;
assign a21340 = ~a21336 & a20736;
assign a21342 = ~a21336 & a20740;
assign a21344 = ~a21336 & a20744;
assign a21346 = ~a21344 & ~a21342;
assign a21348 = a21346 & ~a21340;
assign a21350 = a21348 & ~a21338;
assign a21352 = a21350 & ~a21324;
assign a21354 = a21352 & ~a21322;
assign a21356 = a21354 & ~a21320;
assign a21358 = a21356 & ~a21318;
assign a21360 = a21358 & ~a21300;
assign a21362 = a21360 & ~a20684;
assign a21364 = a21362 & ~a20704;
assign a21366 = a21364 & ~a20708;
assign a21368 = a21366 & ~a20712;
assign a21370 = ~a21368 & a11476;
assign a21372 = ~a21298 & ~a20786;
assign a21374 = ~a21316 & a20788;
assign a21376 = ~a21316 & a20792;
assign a21378 = ~a21316 & a20796;
assign a21380 = ~a21316 & a20800;
assign a21382 = ~a21336 & a20820;
assign a21384 = ~a21336 & a20824;
assign a21386 = ~a21336 & a20828;
assign a21388 = ~a21336 & a20832;
assign a21390 = ~a21388 & ~a21386;
assign a21392 = a21390 & ~a21384;
assign a21394 = a21392 & ~a21382;
assign a21396 = a21394 & ~a21380;
assign a21398 = a21396 & ~a21378;
assign a21400 = a21398 & ~a21376;
assign a21402 = a21400 & ~a21374;
assign a21404 = a21402 & ~a21372;
assign a21406 = a21404 & ~a20804;
assign a21408 = a21406 & ~a20808;
assign a21410 = a21408 & ~a20812;
assign a21412 = a21410 & ~a20816;
assign a21414 = ~a21412 & a11772;
assign a21416 = ~a21298 & ~a20874;
assign a21418 = ~a21316 & a20876;
assign a21420 = ~a21316 & a20880;
assign a21422 = ~a21316 & a20884;
assign a21424 = ~a21316 & a20888;
assign a21426 = ~a21336 & a20908;
assign a21428 = ~a21336 & a20912;
assign a21430 = ~a21336 & a20916;
assign a21432 = ~a21336 & a20920;
assign a21434 = ~a21432 & ~a21430;
assign a21436 = a21434 & ~a21428;
assign a21438 = a21436 & ~a21426;
assign a21440 = a21438 & ~a21424;
assign a21442 = a21440 & ~a21422;
assign a21444 = a21442 & ~a21420;
assign a21446 = a21444 & ~a21418;
assign a21448 = a21446 & ~a21416;
assign a21450 = a21448 & ~a20892;
assign a21452 = a21450 & ~a20896;
assign a21454 = a21452 & ~a20900;
assign a21456 = a21454 & ~a20904;
assign a21458 = ~a21456 & a12068;
assign a21460 = ~a21298 & ~a20962;
assign a21462 = ~a21316 & a20964;
assign a21464 = ~a21316 & a20968;
assign a21466 = ~a21316 & a20972;
assign a21468 = ~a21316 & a20976;
assign a21470 = ~a21336 & a20996;
assign a21472 = ~a21336 & a21000;
assign a21474 = ~a21336 & a21004;
assign a21476 = ~a21336 & a21008;
assign a21478 = ~a21476 & ~a21474;
assign a21480 = a21478 & ~a21472;
assign a21482 = a21480 & ~a21470;
assign a21484 = a21482 & ~a21468;
assign a21486 = a21484 & ~a21466;
assign a21488 = a21486 & ~a21464;
assign a21490 = a21488 & ~a21462;
assign a21492 = a21490 & ~a21460;
assign a21494 = a21492 & ~a20980;
assign a21496 = a21494 & ~a20984;
assign a21498 = a21496 & ~a20988;
assign a21500 = a21498 & ~a20992;
assign a21502 = ~a21500 & a12364;
assign a21504 = ~a21292 & ~a21068;
assign a21506 = a21504 & a21056;
assign a21508 = a21050 & ~a19522;
assign a21510 = a21284 & ~a19544;
assign a21512 = ~a21510 & ~a21508;
assign a21514 = a21512 & a21506;
assign a21516 = ~a21514 & ~a20632;
assign a21518 = ~a21310 & ~a19546;
assign a21520 = a21518 & a19522;
assign a21522 = ~a21056 & a20648;
assign a21524 = a21302 & ~a19544;
assign a21526 = ~a21524 & ~a21522;
assign a21528 = a21526 & a21520;
assign a21530 = ~a21528 & a20634;
assign a21532 = ~a21528 & a20672;
assign a21534 = ~a21528 & a20676;
assign a21536 = ~a21528 & a20680;
assign a21538 = ~a21086 & ~a19594;
assign a21540 = a21538 & a19544;
assign a21542 = ~a21056 & a20686;
assign a21544 = a21078 & ~a19522;
assign a21546 = ~a21544 & ~a21542;
assign a21548 = a21546 & a21540;
assign a21550 = ~a21548 & a20684;
assign a21552 = ~a21548 & a20704;
assign a21554 = ~a21548 & a20708;
assign a21556 = ~a21548 & a20712;
assign a21558 = ~a21556 & ~a21554;
assign a21560 = a21558 & ~a21552;
assign a21562 = a21560 & ~a21550;
assign a21564 = a21562 & ~a21536;
assign a21566 = a21564 & ~a21534;
assign a21568 = a21566 & ~a21532;
assign a21570 = a21568 & ~a21530;
assign a21572 = a21570 & ~a21516;
assign a21574 = a21572 & ~a20716;
assign a21576 = a21574 & ~a20736;
assign a21578 = a21576 & ~a20740;
assign a21580 = a21578 & ~a20744;
assign a21582 = ~a21580 & a11478;
assign a21584 = ~a21514 & ~a20786;
assign a21586 = ~a21528 & a20788;
assign a21588 = ~a21528 & a20792;
assign a21590 = ~a21528 & a20796;
assign a21592 = ~a21528 & a20800;
assign a21594 = ~a21548 & a20804;
assign a21596 = ~a21548 & a20808;
assign a21598 = ~a21548 & a20812;
assign a21600 = ~a21548 & a20816;
assign a21602 = ~a21600 & ~a21598;
assign a21604 = a21602 & ~a21596;
assign a21606 = a21604 & ~a21594;
assign a21608 = a21606 & ~a21592;
assign a21610 = a21608 & ~a21590;
assign a21612 = a21610 & ~a21588;
assign a21614 = a21612 & ~a21586;
assign a21616 = a21614 & ~a21584;
assign a21618 = a21616 & ~a20820;
assign a21620 = a21618 & ~a20824;
assign a21622 = a21620 & ~a20828;
assign a21624 = a21622 & ~a20832;
assign a21626 = ~a21624 & a11774;
assign a21628 = ~a21514 & ~a20874;
assign a21630 = ~a21528 & a20876;
assign a21632 = ~a21528 & a20880;
assign a21634 = ~a21528 & a20884;
assign a21636 = ~a21528 & a20888;
assign a21638 = ~a21548 & a20892;
assign a21640 = ~a21548 & a20896;
assign a21642 = ~a21548 & a20900;
assign a21644 = ~a21548 & a20904;
assign a21646 = ~a21644 & ~a21642;
assign a21648 = a21646 & ~a21640;
assign a21650 = a21648 & ~a21638;
assign a21652 = a21650 & ~a21636;
assign a21654 = a21652 & ~a21634;
assign a21656 = a21654 & ~a21632;
assign a21658 = a21656 & ~a21630;
assign a21660 = a21658 & ~a21628;
assign a21662 = a21660 & ~a20908;
assign a21664 = a21662 & ~a20912;
assign a21666 = a21664 & ~a20916;
assign a21668 = a21666 & ~a20920;
assign a21670 = ~a21668 & a12070;
assign a21672 = ~a21514 & ~a20962;
assign a21674 = ~a21528 & a20964;
assign a21676 = ~a21528 & a20968;
assign a21678 = ~a21528 & a20972;
assign a21680 = ~a21528 & a20976;
assign a21682 = ~a21548 & a20980;
assign a21684 = ~a21548 & a20984;
assign a21686 = ~a21548 & a20988;
assign a21688 = ~a21548 & a20992;
assign a21690 = ~a21688 & ~a21686;
assign a21692 = a21690 & ~a21684;
assign a21694 = a21692 & ~a21682;
assign a21696 = a21694 & ~a21680;
assign a21698 = a21696 & ~a21678;
assign a21700 = a21698 & ~a21676;
assign a21702 = a21700 & ~a21674;
assign a21704 = a21702 & ~a21672;
assign a21706 = a21704 & ~a20996;
assign a21708 = a21706 & ~a21000;
assign a21710 = a21708 & ~a21004;
assign a21712 = a21710 & ~a21008;
assign a21714 = ~a21712 & a12366;
assign a21716 = ~a10296 & a10290;
assign a21718 = ~a10592 & a10586;
assign a21720 = ~a21718 & ~a21716;
assign a21722 = ~a10888 & a10882;
assign a21724 = ~a21722 & a21720;
assign a21726 = ~a11184 & a11178;
assign a21728 = ~a21726 & a21724;
assign a21730 = ~a11480 & a11474;
assign a21732 = ~a10582 & ~a10286;
assign a21734 = a21732 & ~a10878;
assign a21736 = a21734 & ~a11174;
assign a21738 = ~a20646 & ~a19952;
assign a21740 = ~a20654 & ~a19960;
assign a21742 = ~a21740 & ~a21738;
assign a21744 = a21742 & a21736;
assign a21746 = ~a20646 & a19968;
assign a21748 = ~a20654 & a19972;
assign a21750 = ~a21748 & ~a21746;
assign a21752 = a21750 & a21744;
assign a21754 = ~a21752 & a21730;
assign a21756 = ~a11776 & a11770;
assign a21758 = a21756 & ~a21752;
assign a21760 = ~a12072 & a12066;
assign a21762 = a21760 & ~a21752;
assign a21764 = ~a12368 & a12362;
assign a21766 = a21764 & ~a21752;
assign a21768 = ~a13848 & a13842;
assign a21770 = ~a21736 & ~a19502;
assign a21772 = ~a21770 & ~a20688;
assign a21774 = a21772 & a20646;
assign a21776 = ~a21736 & a19578;
assign a21778 = ~a20654 & a19990;
assign a21780 = ~a21778 & ~a21776;
assign a21782 = a21780 & a21774;
assign a21784 = ~a21782 & a21768;
assign a21786 = ~a14144 & a14138;
assign a21788 = a21786 & ~a21782;
assign a21790 = ~a14440 & a14434;
assign a21792 = a21790 & ~a21782;
assign a21794 = ~a14736 & a14730;
assign a21796 = a21794 & ~a21782;
assign a21798 = ~a15032 & a15026;
assign a21800 = ~a21736 & ~a19516;
assign a21802 = ~a21800 & ~a20720;
assign a21804 = a21802 & a20654;
assign a21806 = ~a21736 & a19620;
assign a21808 = ~a20646 & a20014;
assign a21810 = ~a21808 & ~a21806;
assign a21812 = a21810 & a21804;
assign a21814 = ~a21812 & a21798;
assign a21816 = ~a15328 & a15322;
assign a21818 = a21816 & ~a21812;
assign a21820 = ~a15624 & a15618;
assign a21822 = a21820 & ~a21812;
assign a21824 = ~a15920 & a15914;
assign a21826 = a21824 & ~a21812;
assign a21828 = ~a21826 & ~a21822;
assign a21830 = a21828 & ~a21818;
assign a21832 = a21830 & ~a21814;
assign a21834 = a21832 & ~a21796;
assign a21836 = a21834 & ~a21792;
assign a21838 = a21836 & ~a21788;
assign a21840 = a21838 & ~a21784;
assign a21842 = a21840 & ~a21766;
assign a21844 = a21842 & ~a21762;
assign a21846 = a21844 & ~a21758;
assign a21848 = a21846 & ~a21754;
assign a21850 = a21848 & a21728;
assign a21852 = ~a21850 & a12650;
assign a21854 = ~a10298 & a10290;
assign a21856 = ~a10594 & a10586;
assign a21858 = ~a21856 & ~a21854;
assign a21860 = ~a10890 & a10882;
assign a21862 = ~a21860 & a21858;
assign a21864 = ~a11186 & a11178;
assign a21866 = ~a21864 & a21862;
assign a21868 = ~a11482 & a11474;
assign a21870 = a21868 & ~a21752;
assign a21872 = ~a11778 & a11770;
assign a21874 = a21872 & ~a21752;
assign a21876 = ~a12074 & a12066;
assign a21878 = a21876 & ~a21752;
assign a21880 = ~a12370 & a12362;
assign a21882 = a21880 & ~a21752;
assign a21884 = ~a13850 & a13842;
assign a21886 = a21884 & ~a21782;
assign a21888 = ~a14146 & a14138;
assign a21890 = a21888 & ~a21782;
assign a21892 = ~a14442 & a14434;
assign a21894 = a21892 & ~a21782;
assign a21896 = ~a14738 & a14730;
assign a21898 = a21896 & ~a21782;
assign a21900 = ~a15034 & a15026;
assign a21902 = a21900 & ~a21812;
assign a21904 = ~a15330 & a15322;
assign a21906 = a21904 & ~a21812;
assign a21908 = ~a15626 & a15618;
assign a21910 = a21908 & ~a21812;
assign a21912 = ~a15922 & a15914;
assign a21914 = a21912 & ~a21812;
assign a21916 = ~a21914 & ~a21910;
assign a21918 = a21916 & ~a21906;
assign a21920 = a21918 & ~a21902;
assign a21922 = a21920 & ~a21898;
assign a21924 = a21922 & ~a21894;
assign a21926 = a21924 & ~a21890;
assign a21928 = a21926 & ~a21886;
assign a21930 = a21928 & ~a21882;
assign a21932 = a21930 & ~a21878;
assign a21934 = a21932 & ~a21874;
assign a21936 = a21934 & ~a21870;
assign a21938 = a21936 & a21866;
assign a21940 = ~a21938 & a12946;
assign a21942 = ~a10300 & a10290;
assign a21944 = ~a10596 & a10586;
assign a21946 = ~a21944 & ~a21942;
assign a21948 = ~a10892 & a10882;
assign a21950 = ~a21948 & a21946;
assign a21952 = ~a11188 & a11178;
assign a21954 = ~a21952 & a21950;
assign a21956 = ~a11484 & a11474;
assign a21958 = a21956 & ~a21752;
assign a21960 = ~a11780 & a11770;
assign a21962 = a21960 & ~a21752;
assign a21964 = ~a12076 & a12066;
assign a21966 = a21964 & ~a21752;
assign a21968 = ~a12372 & a12362;
assign a21970 = a21968 & ~a21752;
assign a21972 = ~a13852 & a13842;
assign a21974 = a21972 & ~a21782;
assign a21976 = ~a14148 & a14138;
assign a21978 = a21976 & ~a21782;
assign a21980 = ~a14444 & a14434;
assign a21982 = a21980 & ~a21782;
assign a21984 = ~a14740 & a14730;
assign a21986 = a21984 & ~a21782;
assign a21988 = ~a15036 & a15026;
assign a21990 = a21988 & ~a21812;
assign a21992 = ~a15332 & a15322;
assign a21994 = a21992 & ~a21812;
assign a21996 = ~a15628 & a15618;
assign a21998 = a21996 & ~a21812;
assign a22000 = ~a15924 & a15914;
assign a22002 = a22000 & ~a21812;
assign a22004 = ~a22002 & ~a21998;
assign a22006 = a22004 & ~a21994;
assign a22008 = a22006 & ~a21990;
assign a22010 = a22008 & ~a21986;
assign a22012 = a22010 & ~a21982;
assign a22014 = a22012 & ~a21978;
assign a22016 = a22014 & ~a21974;
assign a22018 = a22016 & ~a21970;
assign a22020 = a22018 & ~a21966;
assign a22022 = a22020 & ~a21962;
assign a22024 = a22022 & ~a21958;
assign a22026 = a22024 & a21954;
assign a22028 = ~a22026 & a13242;
assign a22030 = ~a10302 & a10290;
assign a22032 = ~a10598 & a10586;
assign a22034 = ~a22032 & ~a22030;
assign a22036 = ~a10894 & a10882;
assign a22038 = ~a22036 & a22034;
assign a22040 = ~a11190 & a11178;
assign a22042 = ~a22040 & a22038;
assign a22044 = ~a11486 & a11474;
assign a22046 = a22044 & ~a21752;
assign a22048 = ~a11782 & a11770;
assign a22050 = a22048 & ~a21752;
assign a22052 = ~a12078 & a12066;
assign a22054 = a22052 & ~a21752;
assign a22056 = ~a12374 & a12362;
assign a22058 = a22056 & ~a21752;
assign a22060 = ~a13854 & a13842;
assign a22062 = a22060 & ~a21782;
assign a22064 = ~a14150 & a14138;
assign a22066 = a22064 & ~a21782;
assign a22068 = ~a14446 & a14434;
assign a22070 = a22068 & ~a21782;
assign a22072 = ~a14742 & a14730;
assign a22074 = a22072 & ~a21782;
assign a22076 = ~a15038 & a15026;
assign a22078 = a22076 & ~a21812;
assign a22080 = ~a15334 & a15322;
assign a22082 = a22080 & ~a21812;
assign a22084 = ~a15630 & a15618;
assign a22086 = a22084 & ~a21812;
assign a22088 = ~a15926 & a15914;
assign a22090 = a22088 & ~a21812;
assign a22092 = ~a22090 & ~a22086;
assign a22094 = a22092 & ~a22082;
assign a22096 = a22094 & ~a22078;
assign a22098 = a22096 & ~a22074;
assign a22100 = a22098 & ~a22070;
assign a22102 = a22100 & ~a22066;
assign a22104 = a22102 & ~a22062;
assign a22106 = a22104 & ~a22058;
assign a22108 = a22106 & ~a22054;
assign a22110 = a22108 & ~a22050;
assign a22112 = a22110 & ~a22046;
assign a22114 = a22112 & a22042;
assign a22116 = ~a22114 & a13538;
assign a22118 = ~a11762 & ~a11466;
assign a22120 = a22118 & ~a12058;
assign a22122 = a22120 & ~a12354;
assign a22124 = ~a21048 & ~a19502;
assign a22126 = ~a21056 & ~a19516;
assign a22128 = ~a22126 & ~a22124;
assign a22130 = a22128 & a22122;
assign a22132 = a21064 & ~a19502;
assign a22134 = a21068 & ~a19516;
assign a22136 = ~a22134 & ~a22132;
assign a22138 = a22136 & a22130;
assign a22140 = ~a22138 & ~a21728;
assign a22142 = ~a22122 & ~a20646;
assign a22144 = ~a22142 & ~a19578;
assign a22146 = a22144 & a19502;
assign a22148 = ~a22122 & a20688;
assign a22150 = a21086 & ~a19516;
assign a22152 = ~a22150 & ~a22148;
assign a22154 = a22152 & a22146;
assign a22156 = ~a22154 & a21768;
assign a22158 = ~a22154 & a21786;
assign a22160 = ~a22154 & a21790;
assign a22162 = ~a22154 & a21794;
assign a22164 = ~a22122 & ~a20654;
assign a22166 = ~a22164 & ~a19620;
assign a22168 = a22166 & a19516;
assign a22170 = ~a22122 & a20720;
assign a22172 = a21110 & ~a19502;
assign a22174 = ~a22172 & ~a22170;
assign a22176 = a22174 & a22168;
assign a22178 = ~a22176 & a21798;
assign a22180 = ~a22176 & a21816;
assign a22182 = ~a22176 & a21820;
assign a22184 = ~a22176 & a21824;
assign a22186 = ~a22184 & ~a22182;
assign a22188 = a22186 & ~a22180;
assign a22190 = a22188 & ~a22178;
assign a22192 = a22190 & ~a22162;
assign a22194 = a22192 & ~a22160;
assign a22196 = a22194 & ~a22158;
assign a22198 = a22196 & ~a22156;
assign a22200 = a22198 & ~a22140;
assign a22202 = a22200 & ~a21730;
assign a22204 = a22202 & ~a21756;
assign a22206 = a22204 & ~a21760;
assign a22208 = a22206 & ~a21764;
assign a22210 = ~a22208 & a12654;
assign a22212 = ~a22138 & ~a21866;
assign a22214 = ~a22154 & a21884;
assign a22216 = ~a22154 & a21888;
assign a22218 = ~a22154 & a21892;
assign a22220 = ~a22154 & a21896;
assign a22222 = ~a22176 & a21900;
assign a22224 = ~a22176 & a21904;
assign a22226 = ~a22176 & a21908;
assign a22228 = ~a22176 & a21912;
assign a22230 = ~a22228 & ~a22226;
assign a22232 = a22230 & ~a22224;
assign a22234 = a22232 & ~a22222;
assign a22236 = a22234 & ~a22220;
assign a22238 = a22236 & ~a22218;
assign a22240 = a22238 & ~a22216;
assign a22242 = a22240 & ~a22214;
assign a22244 = a22242 & ~a22212;
assign a22246 = a22244 & ~a21868;
assign a22248 = a22246 & ~a21872;
assign a22250 = a22248 & ~a21876;
assign a22252 = a22250 & ~a21880;
assign a22254 = ~a22252 & a12950;
assign a22256 = ~a22138 & ~a21954;
assign a22258 = ~a22154 & a21972;
assign a22260 = ~a22154 & a21976;
assign a22262 = ~a22154 & a21980;
assign a22264 = ~a22154 & a21984;
assign a22266 = ~a22176 & a21988;
assign a22268 = ~a22176 & a21992;
assign a22270 = ~a22176 & a21996;
assign a22272 = ~a22176 & a22000;
assign a22274 = ~a22272 & ~a22270;
assign a22276 = a22274 & ~a22268;
assign a22278 = a22276 & ~a22266;
assign a22280 = a22278 & ~a22264;
assign a22282 = a22280 & ~a22262;
assign a22284 = a22282 & ~a22260;
assign a22286 = a22284 & ~a22258;
assign a22288 = a22286 & ~a22256;
assign a22290 = a22288 & ~a21956;
assign a22292 = a22290 & ~a21960;
assign a22294 = a22292 & ~a21964;
assign a22296 = a22294 & ~a21968;
assign a22298 = ~a22296 & a13246;
assign a22300 = ~a22138 & ~a22042;
assign a22302 = ~a22154 & a22060;
assign a22304 = ~a22154 & a22064;
assign a22306 = ~a22154 & a22068;
assign a22308 = ~a22154 & a22072;
assign a22310 = ~a22176 & a22076;
assign a22312 = ~a22176 & a22080;
assign a22314 = ~a22176 & a22084;
assign a22316 = ~a22176 & a22088;
assign a22318 = ~a22316 & ~a22314;
assign a22320 = a22318 & ~a22312;
assign a22322 = a22320 & ~a22310;
assign a22324 = a22322 & ~a22308;
assign a22326 = a22324 & ~a22306;
assign a22328 = a22326 & ~a22304;
assign a22330 = a22328 & ~a22302;
assign a22332 = a22330 & ~a22300;
assign a22334 = a22332 & ~a22044;
assign a22336 = a22334 & ~a22048;
assign a22338 = a22336 & ~a22052;
assign a22340 = a22338 & ~a22056;
assign a22342 = ~a22340 & a13542;
assign a22344 = ~a22122 & ~a19952;
assign a22346 = ~a22344 & ~a21064;
assign a22348 = a22346 & a21048;
assign a22350 = a22126 & ~a19952;
assign a22352 = ~a22122 & ~a19960;
assign a22354 = a22352 & ~a19534;
assign a22356 = ~a22354 & ~a22350;
assign a22358 = a22356 & a22348;
assign a22360 = ~a22358 & ~a21728;
assign a22362 = ~a21736 & ~a21048;
assign a22364 = ~a22362 & ~a19968;
assign a22366 = a22364 & a19952;
assign a22368 = a21740 & ~a21048;
assign a22370 = ~a21736 & ~a21056;
assign a22372 = a22370 & ~a19534;
assign a22374 = ~a22372 & ~a22368;
assign a22376 = a22374 & a22366;
assign a22378 = ~a22376 & a21730;
assign a22380 = ~a22376 & a21756;
assign a22382 = ~a22376 & a21760;
assign a22384 = ~a22376 & a21764;
assign a22386 = ~a21110 & ~a20014;
assign a22388 = a22386 & a19534;
assign a22390 = a21800 & ~a21048;
assign a22392 = a22164 & ~a19952;
assign a22394 = ~a22392 & ~a22390;
assign a22396 = a22394 & a22388;
assign a22398 = ~a22396 & a21798;
assign a22400 = ~a22396 & a21816;
assign a22402 = ~a22396 & a21820;
assign a22404 = ~a22396 & a21824;
assign a22406 = ~a22404 & ~a22402;
assign a22408 = a22406 & ~a22400;
assign a22410 = a22408 & ~a22398;
assign a22412 = a22410 & ~a22384;
assign a22414 = a22412 & ~a22382;
assign a22416 = a22414 & ~a22380;
assign a22418 = a22416 & ~a22378;
assign a22420 = a22418 & ~a22360;
assign a22422 = a22420 & ~a21768;
assign a22424 = a22422 & ~a21786;
assign a22426 = a22424 & ~a21790;
assign a22428 = a22426 & ~a21794;
assign a22430 = ~a22428 & a12660;
assign a22432 = ~a22358 & ~a21866;
assign a22434 = ~a22376 & a21868;
assign a22436 = ~a22376 & a21872;
assign a22438 = ~a22376 & a21876;
assign a22440 = ~a22376 & a21880;
assign a22442 = ~a22396 & a21900;
assign a22444 = ~a22396 & a21904;
assign a22446 = ~a22396 & a21908;
assign a22448 = ~a22396 & a21912;
assign a22450 = ~a22448 & ~a22446;
assign a22452 = a22450 & ~a22444;
assign a22454 = a22452 & ~a22442;
assign a22456 = a22454 & ~a22440;
assign a22458 = a22456 & ~a22438;
assign a22460 = a22458 & ~a22436;
assign a22462 = a22460 & ~a22434;
assign a22464 = a22462 & ~a22432;
assign a22466 = a22464 & ~a21884;
assign a22468 = a22466 & ~a21888;
assign a22470 = a22468 & ~a21892;
assign a22472 = a22470 & ~a21896;
assign a22474 = ~a22472 & a12956;
assign a22476 = ~a22358 & ~a21954;
assign a22478 = ~a22376 & a21956;
assign a22480 = ~a22376 & a21960;
assign a22482 = ~a22376 & a21964;
assign a22484 = ~a22376 & a21968;
assign a22486 = ~a22396 & a21988;
assign a22488 = ~a22396 & a21992;
assign a22490 = ~a22396 & a21996;
assign a22492 = ~a22396 & a22000;
assign a22494 = ~a22492 & ~a22490;
assign a22496 = a22494 & ~a22488;
assign a22498 = a22496 & ~a22486;
assign a22500 = a22498 & ~a22484;
assign a22502 = a22500 & ~a22482;
assign a22504 = a22502 & ~a22480;
assign a22506 = a22504 & ~a22478;
assign a22508 = a22506 & ~a22476;
assign a22510 = a22508 & ~a21972;
assign a22512 = a22510 & ~a21976;
assign a22514 = a22512 & ~a21980;
assign a22516 = a22514 & ~a21984;
assign a22518 = ~a22516 & a13252;
assign a22520 = ~a22358 & ~a22042;
assign a22522 = ~a22376 & a22044;
assign a22524 = ~a22376 & a22048;
assign a22526 = ~a22376 & a22052;
assign a22528 = ~a22376 & a22056;
assign a22530 = ~a22396 & a22076;
assign a22532 = ~a22396 & a22080;
assign a22534 = ~a22396 & a22084;
assign a22536 = ~a22396 & a22088;
assign a22538 = ~a22536 & ~a22534;
assign a22540 = a22538 & ~a22532;
assign a22542 = a22540 & ~a22530;
assign a22544 = a22542 & ~a22528;
assign a22546 = a22544 & ~a22526;
assign a22548 = a22546 & ~a22524;
assign a22550 = a22548 & ~a22522;
assign a22552 = a22550 & ~a22520;
assign a22554 = a22552 & ~a22060;
assign a22556 = a22554 & ~a22064;
assign a22558 = a22556 & ~a22068;
assign a22560 = a22558 & ~a22072;
assign a22562 = ~a22560 & a13548;
assign a22564 = ~a22352 & ~a21068;
assign a22566 = a22564 & a21056;
assign a22568 = a22124 & ~a19960;
assign a22570 = a22344 & ~a19544;
assign a22572 = ~a22570 & ~a22568;
assign a22574 = a22572 & a22566;
assign a22576 = ~a22574 & ~a21728;
assign a22578 = ~a22370 & ~a19972;
assign a22580 = a22578 & a19960;
assign a22582 = a21738 & ~a21056;
assign a22584 = a22362 & ~a19544;
assign a22586 = ~a22584 & ~a22582;
assign a22588 = a22586 & a22580;
assign a22590 = ~a22588 & a21730;
assign a22592 = ~a22588 & a21756;
assign a22594 = ~a22588 & a21760;
assign a22596 = ~a22588 & a21764;
assign a22598 = ~a21086 & ~a19990;
assign a22600 = a22598 & a19544;
assign a22602 = a21770 & ~a21056;
assign a22604 = a22142 & ~a19960;
assign a22606 = ~a22604 & ~a22602;
assign a22608 = a22606 & a22600;
assign a22610 = ~a22608 & a21768;
assign a22612 = ~a22608 & a21786;
assign a22614 = ~a22608 & a21790;
assign a22616 = ~a22608 & a21794;
assign a22618 = ~a22616 & ~a22614;
assign a22620 = a22618 & ~a22612;
assign a22622 = a22620 & ~a22610;
assign a22624 = a22622 & ~a22596;
assign a22626 = a22624 & ~a22594;
assign a22628 = a22626 & ~a22592;
assign a22630 = a22628 & ~a22590;
assign a22632 = a22630 & ~a22576;
assign a22634 = a22632 & ~a21798;
assign a22636 = a22634 & ~a21816;
assign a22638 = a22636 & ~a21820;
assign a22640 = a22638 & ~a21824;
assign a22642 = ~a22640 & a12662;
assign a22644 = ~a22574 & ~a21866;
assign a22646 = ~a22588 & a21868;
assign a22648 = ~a22588 & a21872;
assign a22650 = ~a22588 & a21876;
assign a22652 = ~a22588 & a21880;
assign a22654 = ~a22608 & a21884;
assign a22656 = ~a22608 & a21888;
assign a22658 = ~a22608 & a21892;
assign a22660 = ~a22608 & a21896;
assign a22662 = ~a22660 & ~a22658;
assign a22664 = a22662 & ~a22656;
assign a22666 = a22664 & ~a22654;
assign a22668 = a22666 & ~a22652;
assign a22670 = a22668 & ~a22650;
assign a22672 = a22670 & ~a22648;
assign a22674 = a22672 & ~a22646;
assign a22676 = a22674 & ~a22644;
assign a22678 = a22676 & ~a21900;
assign a22680 = a22678 & ~a21904;
assign a22682 = a22680 & ~a21908;
assign a22684 = a22682 & ~a21912;
assign a22686 = ~a22684 & a12958;
assign a22688 = ~a22574 & ~a21954;
assign a22690 = ~a22588 & a21956;
assign a22692 = ~a22588 & a21960;
assign a22694 = ~a22588 & a21964;
assign a22696 = ~a22588 & a21968;
assign a22698 = ~a22608 & a21972;
assign a22700 = ~a22608 & a21976;
assign a22702 = ~a22608 & a21980;
assign a22704 = ~a22608 & a21984;
assign a22706 = ~a22704 & ~a22702;
assign a22708 = a22706 & ~a22700;
assign a22710 = a22708 & ~a22698;
assign a22712 = a22710 & ~a22696;
assign a22714 = a22712 & ~a22694;
assign a22716 = a22714 & ~a22692;
assign a22718 = a22716 & ~a22690;
assign a22720 = a22718 & ~a22688;
assign a22722 = a22720 & ~a21988;
assign a22724 = a22722 & ~a21992;
assign a22726 = a22724 & ~a21996;
assign a22728 = a22726 & ~a22000;
assign a22730 = ~a22728 & a13254;
assign a22732 = ~a22574 & ~a22042;
assign a22734 = ~a22588 & a22044;
assign a22736 = ~a22588 & a22048;
assign a22738 = ~a22588 & a22052;
assign a22740 = ~a22588 & a22056;
assign a22742 = ~a22608 & a22060;
assign a22744 = ~a22608 & a22064;
assign a22746 = ~a22608 & a22068;
assign a22748 = ~a22608 & a22072;
assign a22750 = ~a22748 & ~a22746;
assign a22752 = a22750 & ~a22744;
assign a22754 = a22752 & ~a22742;
assign a22756 = a22754 & ~a22740;
assign a22758 = a22756 & ~a22738;
assign a22760 = a22758 & ~a22736;
assign a22762 = a22760 & ~a22734;
assign a22764 = a22762 & ~a22732;
assign a22766 = a22764 & ~a22076;
assign a22768 = a22766 & ~a22080;
assign a22770 = a22768 & ~a22084;
assign a22772 = a22770 & ~a22088;
assign a22774 = ~a22772 & a13550;
assign a22776 = ~a10296 & a10292;
assign a22778 = ~a10592 & a10588;
assign a22780 = ~a22778 & ~a22776;
assign a22782 = ~a10888 & a10884;
assign a22784 = ~a22782 & a22780;
assign a22786 = ~a11184 & a11180;
assign a22788 = ~a22786 & a22784;
assign a22790 = ~a11480 & a11476;
assign a22792 = ~a20640 & ~a19946;
assign a22794 = ~a22792 & ~a21740;
assign a22796 = a22794 & a21736;
assign a22798 = ~a20640 & a19962;
assign a22800 = ~a20654 & a20196;
assign a22802 = ~a22800 & ~a22798;
assign a22804 = a22802 & a22796;
assign a22806 = ~a22804 & a22790;
assign a22808 = ~a11776 & a11772;
assign a22810 = a22808 & ~a22804;
assign a22812 = ~a12072 & a12068;
assign a22814 = a22812 & ~a22804;
assign a22816 = ~a12368 & a12364;
assign a22818 = a22816 & ~a22804;
assign a22820 = ~a12664 & a12660;
assign a22822 = ~a21736 & ~a19496;
assign a22824 = ~a22822 & ~a20656;
assign a22826 = a22824 & a20640;
assign a22828 = ~a21736 & a19524;
assign a22830 = ~a20654 & a20214;
assign a22832 = ~a22830 & ~a22828;
assign a22834 = a22832 & a22826;
assign a22836 = ~a22834 & a22820;
assign a22838 = ~a12960 & a12956;
assign a22840 = a22838 & ~a22834;
assign a22842 = ~a13256 & a13252;
assign a22844 = a22842 & ~a22834;
assign a22846 = ~a13552 & a13548;
assign a22848 = a22846 & ~a22834;
assign a22850 = ~a15032 & a15028;
assign a22852 = ~a21800 & ~a20718;
assign a22854 = a22852 & a20654;
assign a22856 = ~a21736 & a19618;
assign a22858 = ~a20640 & a20006;
assign a22860 = ~a22858 & ~a22856;
assign a22862 = a22860 & a22854;
assign a22864 = ~a22862 & a22850;
assign a22866 = ~a15328 & a15324;
assign a22868 = a22866 & ~a22862;
assign a22870 = ~a15624 & a15620;
assign a22872 = a22870 & ~a22862;
assign a22874 = ~a15920 & a15916;
assign a22876 = a22874 & ~a22862;
assign a22878 = ~a22876 & ~a22872;
assign a22880 = a22878 & ~a22868;
assign a22882 = a22880 & ~a22864;
assign a22884 = a22882 & ~a22848;
assign a22886 = a22884 & ~a22844;
assign a22888 = a22886 & ~a22840;
assign a22890 = a22888 & ~a22836;
assign a22892 = a22890 & ~a22818;
assign a22894 = a22892 & ~a22814;
assign a22896 = a22894 & ~a22810;
assign a22898 = a22896 & ~a22806;
assign a22900 = a22898 & a22788;
assign a22902 = ~a22900 & a13834;
assign a22904 = ~a10298 & a10292;
assign a22906 = ~a10594 & a10588;
assign a22908 = ~a22906 & ~a22904;
assign a22910 = ~a10890 & a10884;
assign a22912 = ~a22910 & a22908;
assign a22914 = ~a11186 & a11180;
assign a22916 = ~a22914 & a22912;
assign a22918 = ~a11482 & a11476;
assign a22920 = a22918 & ~a22804;
assign a22922 = ~a11778 & a11772;
assign a22924 = a22922 & ~a22804;
assign a22926 = ~a12074 & a12068;
assign a22928 = a22926 & ~a22804;
assign a22930 = ~a12370 & a12364;
assign a22932 = a22930 & ~a22804;
assign a22934 = ~a12666 & a12660;
assign a22936 = a22934 & ~a22834;
assign a22938 = ~a12962 & a12956;
assign a22940 = a22938 & ~a22834;
assign a22942 = ~a13258 & a13252;
assign a22944 = a22942 & ~a22834;
assign a22946 = ~a13554 & a13548;
assign a22948 = a22946 & ~a22834;
assign a22950 = ~a15034 & a15028;
assign a22952 = a22950 & ~a22862;
assign a22954 = ~a15330 & a15324;
assign a22956 = a22954 & ~a22862;
assign a22958 = ~a15626 & a15620;
assign a22960 = a22958 & ~a22862;
assign a22962 = ~a15922 & a15916;
assign a22964 = a22962 & ~a22862;
assign a22966 = ~a22964 & ~a22960;
assign a22968 = a22966 & ~a22956;
assign a22970 = a22968 & ~a22952;
assign a22972 = a22970 & ~a22948;
assign a22974 = a22972 & ~a22944;
assign a22976 = a22974 & ~a22940;
assign a22978 = a22976 & ~a22936;
assign a22980 = a22978 & ~a22932;
assign a22982 = a22980 & ~a22928;
assign a22984 = a22982 & ~a22924;
assign a22986 = a22984 & ~a22920;
assign a22988 = a22986 & a22916;
assign a22990 = ~a22988 & a14130;
assign a22992 = ~a10300 & a10292;
assign a22994 = ~a10596 & a10588;
assign a22996 = ~a22994 & ~a22992;
assign a22998 = ~a10892 & a10884;
assign a23000 = ~a22998 & a22996;
assign a23002 = ~a11188 & a11180;
assign a23004 = ~a23002 & a23000;
assign a23006 = ~a11484 & a11476;
assign a23008 = a23006 & ~a22804;
assign a23010 = ~a11780 & a11772;
assign a23012 = a23010 & ~a22804;
assign a23014 = ~a12076 & a12068;
assign a23016 = a23014 & ~a22804;
assign a23018 = ~a12372 & a12364;
assign a23020 = a23018 & ~a22804;
assign a23022 = ~a12668 & a12660;
assign a23024 = a23022 & ~a22834;
assign a23026 = ~a12964 & a12956;
assign a23028 = a23026 & ~a22834;
assign a23030 = ~a13260 & a13252;
assign a23032 = a23030 & ~a22834;
assign a23034 = ~a13556 & a13548;
assign a23036 = a23034 & ~a22834;
assign a23038 = ~a15036 & a15028;
assign a23040 = a23038 & ~a22862;
assign a23042 = ~a15332 & a15324;
assign a23044 = a23042 & ~a22862;
assign a23046 = ~a15628 & a15620;
assign a23048 = a23046 & ~a22862;
assign a23050 = ~a15924 & a15916;
assign a23052 = a23050 & ~a22862;
assign a23054 = ~a23052 & ~a23048;
assign a23056 = a23054 & ~a23044;
assign a23058 = a23056 & ~a23040;
assign a23060 = a23058 & ~a23036;
assign a23062 = a23060 & ~a23032;
assign a23064 = a23062 & ~a23028;
assign a23066 = a23064 & ~a23024;
assign a23068 = a23066 & ~a23020;
assign a23070 = a23068 & ~a23016;
assign a23072 = a23070 & ~a23012;
assign a23074 = a23072 & ~a23008;
assign a23076 = a23074 & a23004;
assign a23078 = ~a23076 & a14426;
assign a23080 = ~a10302 & a10292;
assign a23082 = ~a10598 & a10588;
assign a23084 = ~a23082 & ~a23080;
assign a23086 = ~a10894 & a10884;
assign a23088 = ~a23086 & a23084;
assign a23090 = ~a11190 & a11180;
assign a23092 = ~a23090 & a23088;
assign a23094 = ~a11486 & a11476;
assign a23096 = a23094 & ~a22804;
assign a23098 = ~a11782 & a11772;
assign a23100 = a23098 & ~a22804;
assign a23102 = ~a12078 & a12068;
assign a23104 = a23102 & ~a22804;
assign a23106 = ~a12374 & a12364;
assign a23108 = a23106 & ~a22804;
assign a23110 = ~a12670 & a12660;
assign a23112 = a23110 & ~a22834;
assign a23114 = ~a12966 & a12956;
assign a23116 = a23114 & ~a22834;
assign a23118 = ~a13262 & a13252;
assign a23120 = a23118 & ~a22834;
assign a23122 = ~a13558 & a13548;
assign a23124 = a23122 & ~a22834;
assign a23126 = ~a15038 & a15028;
assign a23128 = a23126 & ~a22862;
assign a23130 = ~a15334 & a15324;
assign a23132 = a23130 & ~a22862;
assign a23134 = ~a15630 & a15620;
assign a23136 = a23134 & ~a22862;
assign a23138 = ~a15926 & a15916;
assign a23140 = a23138 & ~a22862;
assign a23142 = ~a23140 & ~a23136;
assign a23144 = a23142 & ~a23132;
assign a23146 = a23144 & ~a23128;
assign a23148 = a23146 & ~a23124;
assign a23150 = a23148 & ~a23120;
assign a23152 = a23150 & ~a23116;
assign a23154 = a23152 & ~a23112;
assign a23156 = a23154 & ~a23108;
assign a23158 = a23156 & ~a23104;
assign a23160 = a23158 & ~a23100;
assign a23162 = a23160 & ~a23096;
assign a23164 = a23162 & a23092;
assign a23166 = ~a23164 & a14722;
assign a23168 = ~a21042 & ~a19496;
assign a23170 = ~a23168 & ~a22126;
assign a23172 = a23170 & a22122;
assign a23174 = a21058 & ~a19496;
assign a23176 = a21292 & ~a19516;
assign a23178 = ~a23176 & ~a23174;
assign a23180 = a23178 & a23172;
assign a23182 = ~a23180 & ~a22788;
assign a23184 = ~a22122 & ~a20640;
assign a23186 = ~a23184 & ~a19524;
assign a23188 = a23186 & a19496;
assign a23190 = ~a22122 & a20656;
assign a23192 = a21310 & ~a19516;
assign a23194 = ~a23192 & ~a23190;
assign a23196 = a23194 & a23188;
assign a23198 = ~a23196 & a22820;
assign a23200 = ~a23196 & a22838;
assign a23202 = ~a23196 & a22842;
assign a23204 = ~a23196 & a22846;
assign a23206 = ~a22164 & ~a19618;
assign a23208 = a23206 & a19516;
assign a23210 = ~a22122 & a20718;
assign a23212 = a21102 & ~a19496;
assign a23214 = ~a23212 & ~a23210;
assign a23216 = a23214 & a23208;
assign a23218 = ~a23216 & a22850;
assign a23220 = ~a23216 & a22866;
assign a23222 = ~a23216 & a22870;
assign a23224 = ~a23216 & a22874;
assign a23226 = ~a23224 & ~a23222;
assign a23228 = a23226 & ~a23220;
assign a23230 = a23228 & ~a23218;
assign a23232 = a23230 & ~a23204;
assign a23234 = a23232 & ~a23202;
assign a23236 = a23234 & ~a23200;
assign a23238 = a23236 & ~a23198;
assign a23240 = a23238 & ~a23182;
assign a23242 = a23240 & ~a22790;
assign a23244 = a23242 & ~a22808;
assign a23246 = a23244 & ~a22812;
assign a23248 = a23246 & ~a22816;
assign a23250 = ~a23248 & a13838;
assign a23252 = ~a23180 & ~a22916;
assign a23254 = ~a23196 & a22934;
assign a23256 = ~a23196 & a22938;
assign a23258 = ~a23196 & a22942;
assign a23260 = ~a23196 & a22946;
assign a23262 = ~a23216 & a22950;
assign a23264 = ~a23216 & a22954;
assign a23266 = ~a23216 & a22958;
assign a23268 = ~a23216 & a22962;
assign a23270 = ~a23268 & ~a23266;
assign a23272 = a23270 & ~a23264;
assign a23274 = a23272 & ~a23262;
assign a23276 = a23274 & ~a23260;
assign a23278 = a23276 & ~a23258;
assign a23280 = a23278 & ~a23256;
assign a23282 = a23280 & ~a23254;
assign a23284 = a23282 & ~a23252;
assign a23286 = a23284 & ~a22918;
assign a23288 = a23286 & ~a22922;
assign a23290 = a23288 & ~a22926;
assign a23292 = a23290 & ~a22930;
assign a23294 = ~a23292 & a14134;
assign a23296 = ~a23180 & ~a23004;
assign a23298 = ~a23196 & a23022;
assign a23300 = ~a23196 & a23026;
assign a23302 = ~a23196 & a23030;
assign a23304 = ~a23196 & a23034;
assign a23306 = ~a23216 & a23038;
assign a23308 = ~a23216 & a23042;
assign a23310 = ~a23216 & a23046;
assign a23312 = ~a23216 & a23050;
assign a23314 = ~a23312 & ~a23310;
assign a23316 = a23314 & ~a23308;
assign a23318 = a23316 & ~a23306;
assign a23320 = a23318 & ~a23304;
assign a23322 = a23320 & ~a23302;
assign a23324 = a23322 & ~a23300;
assign a23326 = a23324 & ~a23298;
assign a23328 = a23326 & ~a23296;
assign a23330 = a23328 & ~a23006;
assign a23332 = a23330 & ~a23010;
assign a23334 = a23332 & ~a23014;
assign a23336 = a23334 & ~a23018;
assign a23338 = ~a23336 & a14430;
assign a23340 = ~a23180 & ~a23092;
assign a23342 = ~a23196 & a23110;
assign a23344 = ~a23196 & a23114;
assign a23346 = ~a23196 & a23118;
assign a23348 = ~a23196 & a23122;
assign a23350 = ~a23216 & a23126;
assign a23352 = ~a23216 & a23130;
assign a23354 = ~a23216 & a23134;
assign a23356 = ~a23216 & a23138;
assign a23358 = ~a23356 & ~a23354;
assign a23360 = a23358 & ~a23352;
assign a23362 = a23360 & ~a23350;
assign a23364 = a23362 & ~a23348;
assign a23366 = a23364 & ~a23346;
assign a23368 = a23366 & ~a23344;
assign a23370 = a23368 & ~a23342;
assign a23372 = a23370 & ~a23340;
assign a23374 = a23372 & ~a23094;
assign a23376 = a23374 & ~a23098;
assign a23378 = a23376 & ~a23102;
assign a23380 = a23378 & ~a23106;
assign a23382 = ~a23380 & a14726;
assign a23384 = ~a22122 & ~a19946;
assign a23386 = ~a23384 & ~a21058;
assign a23388 = a23386 & a21042;
assign a23390 = a22126 & ~a19946;
assign a23392 = a22352 & ~a19588;
assign a23394 = ~a23392 & ~a23390;
assign a23396 = a23394 & a23388;
assign a23398 = ~a23396 & ~a22788;
assign a23400 = ~a21736 & ~a21042;
assign a23402 = ~a23400 & ~a19962;
assign a23404 = a23402 & a19946;
assign a23406 = a21740 & ~a21042;
assign a23408 = a22370 & ~a19588;
assign a23410 = ~a23408 & ~a23406;
assign a23412 = a23410 & a23404;
assign a23414 = ~a23412 & a22790;
assign a23416 = ~a23412 & a22808;
assign a23418 = ~a23412 & a22812;
assign a23420 = ~a23412 & a22816;
assign a23422 = ~a21102 & ~a20006;
assign a23424 = a23422 & a19588;
assign a23426 = a21800 & ~a21042;
assign a23428 = a22164 & ~a19946;
assign a23430 = ~a23428 & ~a23426;
assign a23432 = a23430 & a23424;
assign a23434 = ~a23432 & a22850;
assign a23436 = ~a23432 & a22866;
assign a23438 = ~a23432 & a22870;
assign a23440 = ~a23432 & a22874;
assign a23442 = ~a23440 & ~a23438;
assign a23444 = a23442 & ~a23436;
assign a23446 = a23444 & ~a23434;
assign a23448 = a23446 & ~a23420;
assign a23450 = a23448 & ~a23418;
assign a23452 = a23450 & ~a23416;
assign a23454 = a23452 & ~a23414;
assign a23456 = a23454 & ~a23398;
assign a23458 = a23456 & ~a22820;
assign a23460 = a23458 & ~a22838;
assign a23462 = a23460 & ~a22842;
assign a23464 = a23462 & ~a22846;
assign a23466 = ~a23464 & a13842;
assign a23468 = ~a23396 & ~a22916;
assign a23470 = ~a23412 & a22918;
assign a23472 = ~a23412 & a22922;
assign a23474 = ~a23412 & a22926;
assign a23476 = ~a23412 & a22930;
assign a23478 = ~a23432 & a22950;
assign a23480 = ~a23432 & a22954;
assign a23482 = ~a23432 & a22958;
assign a23484 = ~a23432 & a22962;
assign a23486 = ~a23484 & ~a23482;
assign a23488 = a23486 & ~a23480;
assign a23490 = a23488 & ~a23478;
assign a23492 = a23490 & ~a23476;
assign a23494 = a23492 & ~a23474;
assign a23496 = a23494 & ~a23472;
assign a23498 = a23496 & ~a23470;
assign a23500 = a23498 & ~a23468;
assign a23502 = a23500 & ~a22934;
assign a23504 = a23502 & ~a22938;
assign a23506 = a23504 & ~a22942;
assign a23508 = a23506 & ~a22946;
assign a23510 = ~a23508 & a14138;
assign a23512 = ~a23396 & ~a23004;
assign a23514 = ~a23412 & a23006;
assign a23516 = ~a23412 & a23010;
assign a23518 = ~a23412 & a23014;
assign a23520 = ~a23412 & a23018;
assign a23522 = ~a23432 & a23038;
assign a23524 = ~a23432 & a23042;
assign a23526 = ~a23432 & a23046;
assign a23528 = ~a23432 & a23050;
assign a23530 = ~a23528 & ~a23526;
assign a23532 = a23530 & ~a23524;
assign a23534 = a23532 & ~a23522;
assign a23536 = a23534 & ~a23520;
assign a23538 = a23536 & ~a23518;
assign a23540 = a23538 & ~a23516;
assign a23542 = a23540 & ~a23514;
assign a23544 = a23542 & ~a23512;
assign a23546 = a23544 & ~a23022;
assign a23548 = a23546 & ~a23026;
assign a23550 = a23548 & ~a23030;
assign a23552 = a23550 & ~a23034;
assign a23554 = ~a23552 & a14434;
assign a23556 = ~a23396 & ~a23092;
assign a23558 = ~a23412 & a23094;
assign a23560 = ~a23412 & a23098;
assign a23562 = ~a23412 & a23102;
assign a23564 = ~a23412 & a23106;
assign a23566 = ~a23432 & a23126;
assign a23568 = ~a23432 & a23130;
assign a23570 = ~a23432 & a23134;
assign a23572 = ~a23432 & a23138;
assign a23574 = ~a23572 & ~a23570;
assign a23576 = a23574 & ~a23568;
assign a23578 = a23576 & ~a23566;
assign a23580 = a23578 & ~a23564;
assign a23582 = a23580 & ~a23562;
assign a23584 = a23582 & ~a23560;
assign a23586 = a23584 & ~a23558;
assign a23588 = a23586 & ~a23556;
assign a23590 = a23588 & ~a23110;
assign a23592 = a23590 & ~a23114;
assign a23594 = a23592 & ~a23118;
assign a23596 = a23594 & ~a23122;
assign a23598 = ~a23596 & a14730;
assign a23600 = ~a22352 & ~a21292;
assign a23602 = a23600 & a21056;
assign a23604 = a23168 & ~a19960;
assign a23606 = a23384 & ~a19522;
assign a23608 = ~a23606 & ~a23604;
assign a23610 = a23608 & a23602;
assign a23612 = ~a23610 & ~a22788;
assign a23614 = ~a22370 & ~a20196;
assign a23616 = a23614 & a19960;
assign a23618 = a22792 & ~a21056;
assign a23620 = a23400 & ~a19522;
assign a23622 = ~a23620 & ~a23618;
assign a23624 = a23622 & a23616;
assign a23626 = ~a23624 & a22790;
assign a23628 = ~a23624 & a22808;
assign a23630 = ~a23624 & a22812;
assign a23632 = ~a23624 & a22816;
assign a23634 = ~a21310 & ~a20214;
assign a23636 = a23634 & a19522;
assign a23638 = a22822 & ~a21056;
assign a23640 = a23184 & ~a19960;
assign a23642 = ~a23640 & ~a23638;
assign a23644 = a23642 & a23636;
assign a23646 = ~a23644 & a22820;
assign a23648 = ~a23644 & a22838;
assign a23650 = ~a23644 & a22842;
assign a23652 = ~a23644 & a22846;
assign a23654 = ~a23652 & ~a23650;
assign a23656 = a23654 & ~a23648;
assign a23658 = a23656 & ~a23646;
assign a23660 = a23658 & ~a23632;
assign a23662 = a23660 & ~a23630;
assign a23664 = a23662 & ~a23628;
assign a23666 = a23664 & ~a23626;
assign a23668 = a23666 & ~a23612;
assign a23670 = a23668 & ~a22850;
assign a23672 = a23670 & ~a22866;
assign a23674 = a23672 & ~a22870;
assign a23676 = a23674 & ~a22874;
assign a23678 = ~a23676 & a13846;
assign a23680 = ~a23610 & ~a22916;
assign a23682 = ~a23624 & a22918;
assign a23684 = ~a23624 & a22922;
assign a23686 = ~a23624 & a22926;
assign a23688 = ~a23624 & a22930;
assign a23690 = ~a23644 & a22934;
assign a23692 = ~a23644 & a22938;
assign a23694 = ~a23644 & a22942;
assign a23696 = ~a23644 & a22946;
assign a23698 = ~a23696 & ~a23694;
assign a23700 = a23698 & ~a23692;
assign a23702 = a23700 & ~a23690;
assign a23704 = a23702 & ~a23688;
assign a23706 = a23704 & ~a23686;
assign a23708 = a23706 & ~a23684;
assign a23710 = a23708 & ~a23682;
assign a23712 = a23710 & ~a23680;
assign a23714 = a23712 & ~a22950;
assign a23716 = a23714 & ~a22954;
assign a23718 = a23716 & ~a22958;
assign a23720 = a23718 & ~a22962;
assign a23722 = ~a23720 & a14142;
assign a23724 = ~a23610 & ~a23004;
assign a23726 = ~a23624 & a23006;
assign a23728 = ~a23624 & a23010;
assign a23730 = ~a23624 & a23014;
assign a23732 = ~a23624 & a23018;
assign a23734 = ~a23644 & a23022;
assign a23736 = ~a23644 & a23026;
assign a23738 = ~a23644 & a23030;
assign a23740 = ~a23644 & a23034;
assign a23742 = ~a23740 & ~a23738;
assign a23744 = a23742 & ~a23736;
assign a23746 = a23744 & ~a23734;
assign a23748 = a23746 & ~a23732;
assign a23750 = a23748 & ~a23730;
assign a23752 = a23750 & ~a23728;
assign a23754 = a23752 & ~a23726;
assign a23756 = a23754 & ~a23724;
assign a23758 = a23756 & ~a23038;
assign a23760 = a23758 & ~a23042;
assign a23762 = a23760 & ~a23046;
assign a23764 = a23762 & ~a23050;
assign a23766 = ~a23764 & a14438;
assign a23768 = ~a23610 & ~a23092;
assign a23770 = ~a23624 & a23094;
assign a23772 = ~a23624 & a23098;
assign a23774 = ~a23624 & a23102;
assign a23776 = ~a23624 & a23106;
assign a23778 = ~a23644 & a23110;
assign a23780 = ~a23644 & a23114;
assign a23782 = ~a23644 & a23118;
assign a23784 = ~a23644 & a23122;
assign a23786 = ~a23784 & ~a23782;
assign a23788 = a23786 & ~a23780;
assign a23790 = a23788 & ~a23778;
assign a23792 = a23790 & ~a23776;
assign a23794 = a23792 & ~a23774;
assign a23796 = a23794 & ~a23772;
assign a23798 = a23796 & ~a23770;
assign a23800 = a23798 & ~a23768;
assign a23802 = a23800 & ~a23126;
assign a23804 = a23802 & ~a23130;
assign a23806 = a23804 & ~a23134;
assign a23808 = a23806 & ~a23138;
assign a23810 = ~a23808 & a14734;
assign a23812 = ~a10296 & a10294;
assign a23814 = ~a10592 & a10590;
assign a23816 = ~a23814 & ~a23812;
assign a23818 = ~a10888 & a10886;
assign a23820 = ~a23818 & a23816;
assign a23822 = ~a11184 & a11182;
assign a23824 = ~a23822 & a23820;
assign a23826 = ~a11480 & a11478;
assign a23828 = ~a22792 & ~a21738;
assign a23830 = a23828 & a21736;
assign a23832 = ~a20640 & a19954;
assign a23834 = ~a20646 & a20188;
assign a23836 = ~a23834 & ~a23832;
assign a23838 = a23836 & a23830;
assign a23840 = ~a23838 & a23826;
assign a23842 = ~a11776 & a11774;
assign a23844 = a23842 & ~a23838;
assign a23846 = ~a12072 & a12070;
assign a23848 = a23846 & ~a23838;
assign a23850 = ~a12368 & a12366;
assign a23852 = a23850 & ~a23838;
assign a23854 = ~a12664 & a12662;
assign a23856 = ~a22822 & ~a20648;
assign a23858 = a23856 & a20640;
assign a23860 = ~a21736 & a19510;
assign a23862 = ~a20646 & a20206;
assign a23864 = ~a23862 & ~a23860;
assign a23866 = a23864 & a23858;
assign a23868 = ~a23866 & a23854;
assign a23870 = ~a12960 & a12958;
assign a23872 = a23870 & ~a23866;
assign a23874 = ~a13256 & a13254;
assign a23876 = a23874 & ~a23866;
assign a23878 = ~a13552 & a13550;
assign a23880 = a23878 & ~a23866;
assign a23882 = ~a13848 & a13846;
assign a23884 = ~a21770 & ~a20686;
assign a23886 = a23884 & a20646;
assign a23888 = ~a21736 & a19576;
assign a23890 = ~a20640 & a19982;
assign a23892 = ~a23890 & ~a23888;
assign a23894 = a23892 & a23886;
assign a23896 = ~a23894 & a23882;
assign a23898 = ~a14144 & a14142;
assign a23900 = a23898 & ~a23894;
assign a23902 = ~a14440 & a14438;
assign a23904 = a23902 & ~a23894;
assign a23906 = ~a14736 & a14734;
assign a23908 = a23906 & ~a23894;
assign a23910 = ~a23908 & ~a23904;
assign a23912 = a23910 & ~a23900;
assign a23914 = a23912 & ~a23896;
assign a23916 = a23914 & ~a23880;
assign a23918 = a23916 & ~a23876;
assign a23920 = a23918 & ~a23872;
assign a23922 = a23920 & ~a23868;
assign a23924 = a23922 & ~a23852;
assign a23926 = a23924 & ~a23848;
assign a23928 = a23926 & ~a23844;
assign a23930 = a23928 & ~a23840;
assign a23932 = a23930 & a23824;
assign a23934 = ~a23932 & a15018;
assign a23936 = ~a10298 & a10294;
assign a23938 = ~a10594 & a10590;
assign a23940 = ~a23938 & ~a23936;
assign a23942 = ~a10890 & a10886;
assign a23944 = ~a23942 & a23940;
assign a23946 = ~a11186 & a11182;
assign a23948 = ~a23946 & a23944;
assign a23950 = ~a11482 & a11478;
assign a23952 = a23950 & ~a23838;
assign a23954 = ~a11778 & a11774;
assign a23956 = a23954 & ~a23838;
assign a23958 = ~a12074 & a12070;
assign a23960 = a23958 & ~a23838;
assign a23962 = ~a12370 & a12366;
assign a23964 = a23962 & ~a23838;
assign a23966 = ~a12666 & a12662;
assign a23968 = a23966 & ~a23866;
assign a23970 = ~a12962 & a12958;
assign a23972 = a23970 & ~a23866;
assign a23974 = ~a13258 & a13254;
assign a23976 = a23974 & ~a23866;
assign a23978 = ~a13554 & a13550;
assign a23980 = a23978 & ~a23866;
assign a23982 = ~a13850 & a13846;
assign a23984 = a23982 & ~a23894;
assign a23986 = ~a14146 & a14142;
assign a23988 = a23986 & ~a23894;
assign a23990 = ~a14442 & a14438;
assign a23992 = a23990 & ~a23894;
assign a23994 = ~a14738 & a14734;
assign a23996 = a23994 & ~a23894;
assign a23998 = ~a23996 & ~a23992;
assign a24000 = a23998 & ~a23988;
assign a24002 = a24000 & ~a23984;
assign a24004 = a24002 & ~a23980;
assign a24006 = a24004 & ~a23976;
assign a24008 = a24006 & ~a23972;
assign a24010 = a24008 & ~a23968;
assign a24012 = a24010 & ~a23964;
assign a24014 = a24012 & ~a23960;
assign a24016 = a24014 & ~a23956;
assign a24018 = a24016 & ~a23952;
assign a24020 = a24018 & a23948;
assign a24022 = ~a24020 & a15314;
assign a24024 = ~a10300 & a10294;
assign a24026 = ~a10596 & a10590;
assign a24028 = ~a24026 & ~a24024;
assign a24030 = ~a10892 & a10886;
assign a24032 = ~a24030 & a24028;
assign a24034 = ~a11188 & a11182;
assign a24036 = ~a24034 & a24032;
assign a24038 = ~a11484 & a11478;
assign a24040 = a24038 & ~a23838;
assign a24042 = ~a11780 & a11774;
assign a24044 = a24042 & ~a23838;
assign a24046 = ~a12076 & a12070;
assign a24048 = a24046 & ~a23838;
assign a24050 = ~a12372 & a12366;
assign a24052 = a24050 & ~a23838;
assign a24054 = ~a12668 & a12662;
assign a24056 = a24054 & ~a23866;
assign a24058 = ~a12964 & a12958;
assign a24060 = a24058 & ~a23866;
assign a24062 = ~a13260 & a13254;
assign a24064 = a24062 & ~a23866;
assign a24066 = ~a13556 & a13550;
assign a24068 = a24066 & ~a23866;
assign a24070 = ~a13852 & a13846;
assign a24072 = a24070 & ~a23894;
assign a24074 = ~a14148 & a14142;
assign a24076 = a24074 & ~a23894;
assign a24078 = ~a14444 & a14438;
assign a24080 = a24078 & ~a23894;
assign a24082 = ~a14740 & a14734;
assign a24084 = a24082 & ~a23894;
assign a24086 = ~a24084 & ~a24080;
assign a24088 = a24086 & ~a24076;
assign a24090 = a24088 & ~a24072;
assign a24092 = a24090 & ~a24068;
assign a24094 = a24092 & ~a24064;
assign a24096 = a24094 & ~a24060;
assign a24098 = a24096 & ~a24056;
assign a24100 = a24098 & ~a24052;
assign a24102 = a24100 & ~a24048;
assign a24104 = a24102 & ~a24044;
assign a24106 = a24104 & ~a24040;
assign a24108 = a24106 & a24036;
assign a24110 = ~a24108 & a15610;
assign a24112 = ~a10302 & a10294;
assign a24114 = ~a10598 & a10590;
assign a24116 = ~a24114 & ~a24112;
assign a24118 = ~a10894 & a10886;
assign a24120 = ~a24118 & a24116;
assign a24122 = ~a11190 & a11182;
assign a24124 = ~a24122 & a24120;
assign a24126 = ~a11486 & a11478;
assign a24128 = a24126 & ~a23838;
assign a24130 = ~a11782 & a11774;
assign a24132 = a24130 & ~a23838;
assign a24134 = ~a12078 & a12070;
assign a24136 = a24134 & ~a23838;
assign a24138 = ~a12374 & a12366;
assign a24140 = a24138 & ~a23838;
assign a24142 = ~a12670 & a12662;
assign a24144 = a24142 & ~a23866;
assign a24146 = ~a12966 & a12958;
assign a24148 = a24146 & ~a23866;
assign a24150 = ~a13262 & a13254;
assign a24152 = a24150 & ~a23866;
assign a24154 = ~a13558 & a13550;
assign a24156 = a24154 & ~a23866;
assign a24158 = ~a13854 & a13846;
assign a24160 = a24158 & ~a23894;
assign a24162 = ~a14150 & a14142;
assign a24164 = a24162 & ~a23894;
assign a24166 = ~a14446 & a14438;
assign a24168 = a24166 & ~a23894;
assign a24170 = ~a14742 & a14734;
assign a24172 = a24170 & ~a23894;
assign a24174 = ~a24172 & ~a24168;
assign a24176 = a24174 & ~a24164;
assign a24178 = a24176 & ~a24160;
assign a24180 = a24178 & ~a24156;
assign a24182 = a24180 & ~a24152;
assign a24184 = a24182 & ~a24148;
assign a24186 = a24184 & ~a24144;
assign a24188 = a24186 & ~a24140;
assign a24190 = a24188 & ~a24136;
assign a24192 = a24190 & ~a24132;
assign a24194 = a24192 & ~a24128;
assign a24196 = a24194 & a24124;
assign a24198 = ~a24196 & a15906;
assign a24200 = ~a23168 & ~a22124;
assign a24202 = a24200 & a22122;
assign a24204 = a21050 & ~a19496;
assign a24206 = a21284 & ~a19502;
assign a24208 = ~a24206 & ~a24204;
assign a24210 = a24208 & a24202;
assign a24212 = ~a24210 & ~a23824;
assign a24214 = ~a23184 & ~a19510;
assign a24216 = a24214 & a19496;
assign a24218 = ~a22122 & a20648;
assign a24220 = a21302 & ~a19502;
assign a24222 = ~a24220 & ~a24218;
assign a24224 = a24222 & a24216;
assign a24226 = ~a24224 & a23854;
assign a24228 = ~a24224 & a23870;
assign a24230 = ~a24224 & a23874;
assign a24232 = ~a24224 & a23878;
assign a24234 = ~a22142 & ~a19576;
assign a24236 = a24234 & a19502;
assign a24238 = ~a22122 & a20686;
assign a24240 = a21078 & ~a19496;
assign a24242 = ~a24240 & ~a24238;
assign a24244 = a24242 & a24236;
assign a24246 = ~a24244 & a23882;
assign a24248 = ~a24244 & a23898;
assign a24250 = ~a24244 & a23902;
assign a24252 = ~a24244 & a23906;
assign a24254 = ~a24252 & ~a24250;
assign a24256 = a24254 & ~a24248;
assign a24258 = a24256 & ~a24246;
assign a24260 = a24258 & ~a24232;
assign a24262 = a24260 & ~a24230;
assign a24264 = a24262 & ~a24228;
assign a24266 = a24264 & ~a24226;
assign a24268 = a24266 & ~a24212;
assign a24270 = a24268 & ~a23826;
assign a24272 = a24270 & ~a23842;
assign a24274 = a24272 & ~a23846;
assign a24276 = a24274 & ~a23850;
assign a24278 = ~a24276 & a15022;
assign a24280 = ~a24210 & ~a23948;
assign a24282 = ~a24224 & a23966;
assign a24284 = ~a24224 & a23970;
assign a24286 = ~a24224 & a23974;
assign a24288 = ~a24224 & a23978;
assign a24290 = ~a24244 & a23982;
assign a24292 = ~a24244 & a23986;
assign a24294 = ~a24244 & a23990;
assign a24296 = ~a24244 & a23994;
assign a24298 = ~a24296 & ~a24294;
assign a24300 = a24298 & ~a24292;
assign a24302 = a24300 & ~a24290;
assign a24304 = a24302 & ~a24288;
assign a24306 = a24304 & ~a24286;
assign a24308 = a24306 & ~a24284;
assign a24310 = a24308 & ~a24282;
assign a24312 = a24310 & ~a24280;
assign a24314 = a24312 & ~a23950;
assign a24316 = a24314 & ~a23954;
assign a24318 = a24316 & ~a23958;
assign a24320 = a24318 & ~a23962;
assign a24322 = ~a24320 & a15318;
assign a24324 = ~a24210 & ~a24036;
assign a24326 = ~a24224 & a24054;
assign a24328 = ~a24224 & a24058;
assign a24330 = ~a24224 & a24062;
assign a24332 = ~a24224 & a24066;
assign a24334 = ~a24244 & a24070;
assign a24336 = ~a24244 & a24074;
assign a24338 = ~a24244 & a24078;
assign a24340 = ~a24244 & a24082;
assign a24342 = ~a24340 & ~a24338;
assign a24344 = a24342 & ~a24336;
assign a24346 = a24344 & ~a24334;
assign a24348 = a24346 & ~a24332;
assign a24350 = a24348 & ~a24330;
assign a24352 = a24350 & ~a24328;
assign a24354 = a24352 & ~a24326;
assign a24356 = a24354 & ~a24324;
assign a24358 = a24356 & ~a24038;
assign a24360 = a24358 & ~a24042;
assign a24362 = a24360 & ~a24046;
assign a24364 = a24362 & ~a24050;
assign a24366 = ~a24364 & a15614;
assign a24368 = ~a24210 & ~a24124;
assign a24370 = ~a24224 & a24142;
assign a24372 = ~a24224 & a24146;
assign a24374 = ~a24224 & a24150;
assign a24376 = ~a24224 & a24154;
assign a24378 = ~a24244 & a24158;
assign a24380 = ~a24244 & a24162;
assign a24382 = ~a24244 & a24166;
assign a24384 = ~a24244 & a24170;
assign a24386 = ~a24384 & ~a24382;
assign a24388 = a24386 & ~a24380;
assign a24390 = a24388 & ~a24378;
assign a24392 = a24390 & ~a24376;
assign a24394 = a24392 & ~a24374;
assign a24396 = a24394 & ~a24372;
assign a24398 = a24396 & ~a24370;
assign a24400 = a24398 & ~a24368;
assign a24402 = a24400 & ~a24126;
assign a24404 = a24402 & ~a24130;
assign a24406 = a24404 & ~a24134;
assign a24408 = a24406 & ~a24138;
assign a24410 = ~a24408 & a15910;
assign a24412 = ~a23384 & ~a21050;
assign a24414 = a24412 & a21042;
assign a24416 = a22124 & ~a19946;
assign a24418 = a22344 & ~a19574;
assign a24420 = ~a24418 & ~a24416;
assign a24422 = a24420 & a24414;
assign a24424 = ~a24422 & ~a23824;
assign a24426 = ~a23400 & ~a19954;
assign a24428 = a24426 & a19946;
assign a24430 = a21738 & ~a21042;
assign a24432 = a22362 & ~a19574;
assign a24434 = ~a24432 & ~a24430;
assign a24436 = a24434 & a24428;
assign a24438 = ~a24436 & a23826;
assign a24440 = ~a24436 & a23842;
assign a24442 = ~a24436 & a23846;
assign a24444 = ~a24436 & a23850;
assign a24446 = ~a21078 & ~a19982;
assign a24448 = a24446 & a19574;
assign a24450 = a21770 & ~a21042;
assign a24452 = a22142 & ~a19946;
assign a24454 = ~a24452 & ~a24450;
assign a24456 = a24454 & a24448;
assign a24458 = ~a24456 & a23882;
assign a24460 = ~a24456 & a23898;
assign a24462 = ~a24456 & a23902;
assign a24464 = ~a24456 & a23906;
assign a24466 = ~a24464 & ~a24462;
assign a24468 = a24466 & ~a24460;
assign a24470 = a24468 & ~a24458;
assign a24472 = a24470 & ~a24444;
assign a24474 = a24472 & ~a24442;
assign a24476 = a24474 & ~a24440;
assign a24478 = a24476 & ~a24438;
assign a24480 = a24478 & ~a24424;
assign a24482 = a24480 & ~a23854;
assign a24484 = a24482 & ~a23870;
assign a24486 = a24484 & ~a23874;
assign a24488 = a24486 & ~a23878;
assign a24490 = ~a24488 & a15026;
assign a24492 = ~a24422 & ~a23948;
assign a24494 = ~a24436 & a23950;
assign a24496 = ~a24436 & a23954;
assign a24498 = ~a24436 & a23958;
assign a24500 = ~a24436 & a23962;
assign a24502 = ~a24456 & a23982;
assign a24504 = ~a24456 & a23986;
assign a24506 = ~a24456 & a23990;
assign a24508 = ~a24456 & a23994;
assign a24510 = ~a24508 & ~a24506;
assign a24512 = a24510 & ~a24504;
assign a24514 = a24512 & ~a24502;
assign a24516 = a24514 & ~a24500;
assign a24518 = a24516 & ~a24498;
assign a24520 = a24518 & ~a24496;
assign a24522 = a24520 & ~a24494;
assign a24524 = a24522 & ~a24492;
assign a24526 = a24524 & ~a23966;
assign a24528 = a24526 & ~a23970;
assign a24530 = a24528 & ~a23974;
assign a24532 = a24530 & ~a23978;
assign a24534 = ~a24532 & a15322;
assign a24536 = ~a24422 & ~a24036;
assign a24538 = ~a24436 & a24038;
assign a24540 = ~a24436 & a24042;
assign a24542 = ~a24436 & a24046;
assign a24544 = ~a24436 & a24050;
assign a24546 = ~a24456 & a24070;
assign a24548 = ~a24456 & a24074;
assign a24550 = ~a24456 & a24078;
assign a24552 = ~a24456 & a24082;
assign a24554 = ~a24552 & ~a24550;
assign a24556 = a24554 & ~a24548;
assign a24558 = a24556 & ~a24546;
assign a24560 = a24558 & ~a24544;
assign a24562 = a24560 & ~a24542;
assign a24564 = a24562 & ~a24540;
assign a24566 = a24564 & ~a24538;
assign a24568 = a24566 & ~a24536;
assign a24570 = a24568 & ~a24054;
assign a24572 = a24570 & ~a24058;
assign a24574 = a24572 & ~a24062;
assign a24576 = a24574 & ~a24066;
assign a24578 = ~a24576 & a15618;
assign a24580 = ~a24422 & ~a24124;
assign a24582 = ~a24436 & a24126;
assign a24584 = ~a24436 & a24130;
assign a24586 = ~a24436 & a24134;
assign a24588 = ~a24436 & a24138;
assign a24590 = ~a24456 & a24158;
assign a24592 = ~a24456 & a24162;
assign a24594 = ~a24456 & a24166;
assign a24596 = ~a24456 & a24170;
assign a24598 = ~a24596 & ~a24594;
assign a24600 = a24598 & ~a24592;
assign a24602 = a24600 & ~a24590;
assign a24604 = a24602 & ~a24588;
assign a24606 = a24604 & ~a24586;
assign a24608 = a24606 & ~a24584;
assign a24610 = a24608 & ~a24582;
assign a24612 = a24610 & ~a24580;
assign a24614 = a24612 & ~a24142;
assign a24616 = a24614 & ~a24146;
assign a24618 = a24616 & ~a24150;
assign a24620 = a24618 & ~a24154;
assign a24622 = ~a24620 & a15914;
assign a24624 = ~a22344 & ~a21284;
assign a24626 = a24624 & a21048;
assign a24628 = a23168 & ~a19952;
assign a24630 = a23384 & ~a19508;
assign a24632 = ~a24630 & ~a24628;
assign a24634 = a24632 & a24626;
assign a24636 = ~a24634 & ~a23824;
assign a24638 = ~a22362 & ~a20188;
assign a24640 = a24638 & a19952;
assign a24642 = a22792 & ~a21048;
assign a24644 = a23400 & ~a19508;
assign a24646 = ~a24644 & ~a24642;
assign a24648 = a24646 & a24640;
assign a24650 = ~a24648 & a23826;
assign a24652 = ~a24648 & a23842;
assign a24654 = ~a24648 & a23846;
assign a24656 = ~a24648 & a23850;
assign a24658 = ~a21302 & ~a20206;
assign a24660 = a24658 & a19508;
assign a24662 = a22822 & ~a21048;
assign a24664 = a23184 & ~a19952;
assign a24666 = ~a24664 & ~a24662;
assign a24668 = a24666 & a24660;
assign a24670 = ~a24668 & a23854;
assign a24672 = ~a24668 & a23870;
assign a24674 = ~a24668 & a23874;
assign a24676 = ~a24668 & a23878;
assign a24678 = ~a24676 & ~a24674;
assign a24680 = a24678 & ~a24672;
assign a24682 = a24680 & ~a24670;
assign a24684 = a24682 & ~a24656;
assign a24686 = a24684 & ~a24654;
assign a24688 = a24686 & ~a24652;
assign a24690 = a24688 & ~a24650;
assign a24692 = a24690 & ~a24636;
assign a24694 = a24692 & ~a23882;
assign a24696 = a24694 & ~a23898;
assign a24698 = a24696 & ~a23902;
assign a24700 = a24698 & ~a23906;
assign a24702 = ~a24700 & a15028;
assign a24704 = ~a24634 & ~a23948;
assign a24706 = ~a24648 & a23950;
assign a24708 = ~a24648 & a23954;
assign a24710 = ~a24648 & a23958;
assign a24712 = ~a24648 & a23962;
assign a24714 = ~a24668 & a23966;
assign a24716 = ~a24668 & a23970;
assign a24718 = ~a24668 & a23974;
assign a24720 = ~a24668 & a23978;
assign a24722 = ~a24720 & ~a24718;
assign a24724 = a24722 & ~a24716;
assign a24726 = a24724 & ~a24714;
assign a24728 = a24726 & ~a24712;
assign a24730 = a24728 & ~a24710;
assign a24732 = a24730 & ~a24708;
assign a24734 = a24732 & ~a24706;
assign a24736 = a24734 & ~a24704;
assign a24738 = a24736 & ~a23982;
assign a24740 = a24738 & ~a23986;
assign a24742 = a24740 & ~a23990;
assign a24744 = a24742 & ~a23994;
assign a24746 = ~a24744 & a15324;
assign a24748 = ~a24634 & ~a24036;
assign a24750 = ~a24648 & a24038;
assign a24752 = ~a24648 & a24042;
assign a24754 = ~a24648 & a24046;
assign a24756 = ~a24648 & a24050;
assign a24758 = ~a24668 & a24054;
assign a24760 = ~a24668 & a24058;
assign a24762 = ~a24668 & a24062;
assign a24764 = ~a24668 & a24066;
assign a24766 = ~a24764 & ~a24762;
assign a24768 = a24766 & ~a24760;
assign a24770 = a24768 & ~a24758;
assign a24772 = a24770 & ~a24756;
assign a24774 = a24772 & ~a24754;
assign a24776 = a24774 & ~a24752;
assign a24778 = a24776 & ~a24750;
assign a24780 = a24778 & ~a24748;
assign a24782 = a24780 & ~a24070;
assign a24784 = a24782 & ~a24074;
assign a24786 = a24784 & ~a24078;
assign a24788 = a24786 & ~a24082;
assign a24790 = ~a24788 & a15620;
assign a24792 = ~a24634 & ~a24124;
assign a24794 = ~a24648 & a24126;
assign a24796 = ~a24648 & a24130;
assign a24798 = ~a24648 & a24134;
assign a24800 = ~a24648 & a24138;
assign a24802 = ~a24668 & a24142;
assign a24804 = ~a24668 & a24146;
assign a24806 = ~a24668 & a24150;
assign a24808 = ~a24668 & a24154;
assign a24810 = ~a24808 & ~a24806;
assign a24812 = a24810 & ~a24804;
assign a24814 = a24812 & ~a24802;
assign a24816 = a24814 & ~a24800;
assign a24818 = a24816 & ~a24798;
assign a24820 = a24818 & ~a24796;
assign a24822 = a24820 & ~a24794;
assign a24824 = a24822 & ~a24792;
assign a24826 = a24824 & ~a24158;
assign a24828 = a24826 & ~a24162;
assign a24830 = a24828 & ~a24166;
assign a24832 = a24830 & ~a24170;
assign a24834 = ~a24832 & a15916;
assign a24836 = ~a20640 & ~a19964;
assign a24838 = ~a20646 & ~a20190;
assign a24840 = ~a20654 & ~a20408;
assign a24842 = ~a20640 & ~a19976;
assign a24844 = ~a20646 & ~a20200;
assign a24846 = ~a20654 & ~a20416;
assign a24848 = ~a24846 & ~a24844;
assign a24850 = a24848 & ~a24842;
assign a24852 = a24850 & ~a24840;
assign a24854 = a24852 & ~a24838;
assign a24856 = a24854 & ~a24836;
assign a24858 = a24856 & a23828;
assign a24860 = a24858 & ~a21740;
assign a24862 = a24860 & a21736;
assign a24864 = ~a22122 & ~a20658;
assign a24866 = ~a21304 & ~a19502;
assign a24868 = ~a21518 & ~a19516;
assign a24870 = ~a22122 & ~a20666;
assign a24872 = ~a21314 & ~a19502;
assign a24874 = ~a21526 & ~a19516;
assign a24876 = ~a24874 & ~a24872;
assign a24878 = a24876 & ~a24870;
assign a24880 = a24878 & ~a24868;
assign a24882 = a24880 & ~a24866;
assign a24884 = a24882 & ~a24864;
assign a24886 = a24884 & a24214;
assign a24888 = a24886 & ~a19524;
assign a24890 = a24888 & a19496;
assign a24892 = ~a21772 & ~a21042;
assign a24894 = ~a22144 & ~a19946;
assign a24896 = ~a22598 & ~a19588;
assign a24898 = ~a21780 & ~a21042;
assign a24900 = ~a22152 & ~a19946;
assign a24902 = ~a22606 & ~a19588;
assign a24904 = ~a24902 & ~a24900;
assign a24906 = a24904 & ~a24898;
assign a24908 = a24906 & ~a24896;
assign a24910 = a24908 & ~a24894;
assign a24912 = a24910 & ~a24892;
assign a24914 = a24912 & a24446;
assign a24916 = a24914 & ~a19590;
assign a24918 = a24916 & a19574;
assign a24920 = ~a22852 & ~a21048;
assign a24922 = ~a23206 & ~a19952;
assign a24924 = ~a23422 & ~a19508;
assign a24926 = ~a22860 & ~a21048;
assign a24928 = ~a23214 & ~a19952;
assign a24930 = ~a23430 & ~a19508;
assign a24932 = ~a24930 & ~a24928;
assign a24934 = a24932 & ~a24926;
assign a24936 = a24934 & ~a24924;
assign a24938 = a24936 & ~a24922;
assign a24940 = a24938 & ~a24920;
assign a24942 = a24940 & a22386;
assign a24944 = a24942 & ~a19630;
assign a24946 = a24944 & a19534;
assign a24948 = a10278 & l938;
assign a24950 = ~a10278 & ~l938;
assign a24952 = ~a24950 & ~a24948;
assign a24954 = a10574 & l952;
assign a24956 = ~a10574 & ~l952;
assign a24958 = ~a24956 & ~a24954;
assign a24960 = a10870 & l966;
assign a24962 = ~a10870 & ~l966;
assign a24964 = ~a24962 & ~a24960;
assign a24966 = a11166 & l980;
assign a24968 = ~a11166 & ~l980;
assign a24970 = ~a24968 & ~a24966;
assign a24972 = a11462 & l1022;
assign a24974 = ~a11462 & ~l1022;
assign a24976 = ~a24974 & ~a24972;
assign a24978 = a11758 & l1036;
assign a24980 = ~a11758 & ~l1036;
assign a24982 = ~a24980 & ~a24978;
assign a24984 = a12054 & l1050;
assign a24986 = ~a12054 & ~l1050;
assign a24988 = ~a24986 & ~a24984;
assign a24990 = a12350 & l1064;
assign a24992 = ~a12350 & ~l1064;
assign a24994 = ~a24992 & ~a24990;
assign a24996 = a12646 & l1106;
assign a24998 = ~a12646 & ~l1106;
assign a25000 = ~a24998 & ~a24996;
assign a25002 = a12942 & l1120;
assign a25004 = ~a12942 & ~l1120;
assign a25006 = ~a25004 & ~a25002;
assign a25008 = a13238 & l1134;
assign a25010 = ~a13238 & ~l1134;
assign a25012 = ~a25010 & ~a25008;
assign a25014 = a13534 & l1148;
assign a25016 = ~a13534 & ~l1148;
assign a25018 = ~a25016 & ~a25014;
assign a25020 = a13830 & l1190;
assign a25022 = ~a13830 & ~l1190;
assign a25024 = ~a25022 & ~a25020;
assign a25026 = a14126 & l1204;
assign a25028 = ~a14126 & ~l1204;
assign a25030 = ~a25028 & ~a25026;
assign a25032 = a14422 & l1218;
assign a25034 = ~a14422 & ~l1218;
assign a25036 = ~a25034 & ~a25032;
assign a25038 = a14718 & l1232;
assign a25040 = ~a14718 & ~l1232;
assign a25042 = ~a25040 & ~a25038;
assign a25044 = a15014 & l1274;
assign a25046 = ~a15014 & ~l1274;
assign a25048 = ~a25046 & ~a25044;
assign a25050 = a15310 & l1288;
assign a25052 = ~a15310 & ~l1288;
assign a25054 = ~a25052 & ~a25050;
assign a25056 = a15606 & l1302;
assign a25058 = ~a15606 & ~l1302;
assign a25060 = ~a25058 & ~a25056;
assign a25062 = a15902 & l1316;
assign a25064 = ~a15902 & ~l1316;
assign a25066 = ~a25064 & ~a25062;
assign a25068 = ~l1360 & ~l936;
assign a25070 = l1360 & l936;
assign a25072 = ~a25070 & ~a25068;
assign a25074 = ~l1358 & l934;
assign a25076 = l1358 & ~l934;
assign a25078 = ~a25076 & ~a25074;
assign a25080 = ~l1364 & ~l942;
assign a25082 = l1364 & l942;
assign a25084 = ~a25082 & ~a25080;
assign a25086 = ~l1362 & l940;
assign a25088 = l1362 & ~l940;
assign a25090 = ~a25088 & ~a25086;
assign a25092 = ~l1368 & ~l950;
assign a25094 = l1368 & l950;
assign a25096 = ~a25094 & ~a25092;
assign a25098 = ~l1366 & l948;
assign a25100 = l1366 & ~l948;
assign a25102 = ~a25100 & ~a25098;
assign a25104 = ~l1372 & ~l956;
assign a25106 = l1372 & l956;
assign a25108 = ~a25106 & ~a25104;
assign a25110 = ~l1370 & l954;
assign a25112 = l1370 & ~l954;
assign a25114 = ~a25112 & ~a25110;
assign a25116 = ~l1376 & ~l964;
assign a25118 = l1376 & l964;
assign a25120 = ~a25118 & ~a25116;
assign a25122 = ~l1374 & l962;
assign a25124 = l1374 & ~l962;
assign a25126 = ~a25124 & ~a25122;
assign a25128 = ~l1380 & ~l970;
assign a25130 = l1380 & l970;
assign a25132 = ~a25130 & ~a25128;
assign a25134 = ~l1378 & l968;
assign a25136 = l1378 & ~l968;
assign a25138 = ~a25136 & ~a25134;
assign a25140 = ~l1384 & ~l978;
assign a25142 = l1384 & l978;
assign a25144 = ~a25142 & ~a25140;
assign a25146 = ~l1382 & l976;
assign a25148 = l1382 & ~l976;
assign a25150 = ~a25148 & ~a25146;
assign a25152 = ~l1388 & ~l984;
assign a25154 = l1388 & l984;
assign a25156 = ~a25154 & ~a25152;
assign a25158 = ~l1386 & l982;
assign a25160 = l1386 & ~l982;
assign a25162 = ~a25160 & ~a25158;
assign a25164 = ~l1394 & ~l990;
assign a25166 = l1394 & l990;
assign a25168 = ~a25166 & ~a25164;
assign a25170 = ~l1392 & l988;
assign a25172 = l1392 & ~l988;
assign a25174 = ~a25172 & ~a25170;
assign a25176 = ~l1390 & l986;
assign a25178 = l1390 & ~l986;
assign a25180 = ~a25178 & ~a25176;
assign a25182 = ~l1396 & l992;
assign a25184 = l1396 & ~l992;
assign a25186 = ~a25184 & ~a25182;
assign a25188 = ~l1400 & l996;
assign a25190 = l1400 & ~l996;
assign a25192 = ~a25190 & ~a25188;
assign a25194 = ~l1398 & l994;
assign a25196 = l1398 & ~l994;
assign a25198 = ~a25196 & ~a25194;
assign a25200 = ~l1402 & l1000;
assign a25202 = l1402 & ~l1000;
assign a25204 = ~a25202 & ~a25200;
assign a25206 = ~l1404 & l1002;
assign a25208 = l1404 & ~l1002;
assign a25210 = ~a25208 & ~a25206;
assign a25212 = ~l1414 & l1012;
assign a25214 = l1414 & ~l1012;
assign a25216 = ~a25214 & ~a25212;
assign a25218 = ~l1412 & l1010;
assign a25220 = l1412 & ~l1010;
assign a25222 = ~a25220 & ~a25218;
assign a25224 = ~l1410 & l1008;
assign a25226 = l1410 & ~l1008;
assign a25228 = ~a25226 & ~a25224;
assign a25230 = ~l1408 & l1006;
assign a25232 = l1408 & ~l1006;
assign a25234 = ~a25232 & ~a25230;
assign a25236 = ~l1406 & l1004;
assign a25238 = l1406 & ~l1004;
assign a25240 = ~a25238 & ~a25236;
assign a25242 = ~l1418 & ~l1020;
assign a25244 = l1418 & l1020;
assign a25246 = ~a25244 & ~a25242;
assign a25248 = ~l1416 & l1018;
assign a25250 = l1416 & ~l1018;
assign a25252 = ~a25250 & ~a25248;
assign a25254 = ~l1422 & ~l1026;
assign a25256 = l1422 & l1026;
assign a25258 = ~a25256 & ~a25254;
assign a25260 = ~l1420 & l1024;
assign a25262 = l1420 & ~l1024;
assign a25264 = ~a25262 & ~a25260;
assign a25266 = ~l1426 & ~l1034;
assign a25268 = l1426 & l1034;
assign a25270 = ~a25268 & ~a25266;
assign a25272 = ~l1424 & l1032;
assign a25274 = l1424 & ~l1032;
assign a25276 = ~a25274 & ~a25272;
assign a25278 = ~l1430 & ~l1040;
assign a25280 = l1430 & l1040;
assign a25282 = ~a25280 & ~a25278;
assign a25284 = ~l1428 & l1038;
assign a25286 = l1428 & ~l1038;
assign a25288 = ~a25286 & ~a25284;
assign a25290 = ~l1434 & ~l1048;
assign a25292 = l1434 & l1048;
assign a25294 = ~a25292 & ~a25290;
assign a25296 = ~l1432 & l1046;
assign a25298 = l1432 & ~l1046;
assign a25300 = ~a25298 & ~a25296;
assign a25302 = ~l1438 & ~l1054;
assign a25304 = l1438 & l1054;
assign a25306 = ~a25304 & ~a25302;
assign a25308 = ~l1436 & l1052;
assign a25310 = l1436 & ~l1052;
assign a25312 = ~a25310 & ~a25308;
assign a25314 = ~l1442 & ~l1062;
assign a25316 = l1442 & l1062;
assign a25318 = ~a25316 & ~a25314;
assign a25320 = ~l1440 & l1060;
assign a25322 = l1440 & ~l1060;
assign a25324 = ~a25322 & ~a25320;
assign a25326 = ~l1446 & ~l1068;
assign a25328 = l1446 & l1068;
assign a25330 = ~a25328 & ~a25326;
assign a25332 = ~l1444 & l1066;
assign a25334 = l1444 & ~l1066;
assign a25336 = ~a25334 & ~a25332;
assign a25338 = ~l1452 & ~l1074;
assign a25340 = l1452 & l1074;
assign a25342 = ~a25340 & ~a25338;
assign a25344 = ~l1450 & l1072;
assign a25346 = l1450 & ~l1072;
assign a25348 = ~a25346 & ~a25344;
assign a25350 = ~l1448 & l1070;
assign a25352 = l1448 & ~l1070;
assign a25354 = ~a25352 & ~a25350;
assign a25356 = ~l1454 & l1076;
assign a25358 = l1454 & ~l1076;
assign a25360 = ~a25358 & ~a25356;
assign a25362 = ~l1458 & l1080;
assign a25364 = l1458 & ~l1080;
assign a25366 = ~a25364 & ~a25362;
assign a25368 = ~l1456 & l1078;
assign a25370 = l1456 & ~l1078;
assign a25372 = ~a25370 & ~a25368;
assign a25374 = ~l1460 & l1084;
assign a25376 = l1460 & ~l1084;
assign a25378 = ~a25376 & ~a25374;
assign a25380 = ~l1462 & l1086;
assign a25382 = l1462 & ~l1086;
assign a25384 = ~a25382 & ~a25380;
assign a25386 = ~l1472 & l1096;
assign a25388 = l1472 & ~l1096;
assign a25390 = ~a25388 & ~a25386;
assign a25392 = ~l1470 & l1094;
assign a25394 = l1470 & ~l1094;
assign a25396 = ~a25394 & ~a25392;
assign a25398 = ~l1468 & l1092;
assign a25400 = l1468 & ~l1092;
assign a25402 = ~a25400 & ~a25398;
assign a25404 = ~l1466 & l1090;
assign a25406 = l1466 & ~l1090;
assign a25408 = ~a25406 & ~a25404;
assign a25410 = ~l1464 & l1088;
assign a25412 = l1464 & ~l1088;
assign a25414 = ~a25412 & ~a25410;
assign a25416 = ~l1476 & ~l1104;
assign a25418 = l1476 & l1104;
assign a25420 = ~a25418 & ~a25416;
assign a25422 = ~l1474 & l1102;
assign a25424 = l1474 & ~l1102;
assign a25426 = ~a25424 & ~a25422;
assign a25428 = ~l1480 & ~l1110;
assign a25430 = l1480 & l1110;
assign a25432 = ~a25430 & ~a25428;
assign a25434 = ~l1478 & l1108;
assign a25436 = l1478 & ~l1108;
assign a25438 = ~a25436 & ~a25434;
assign a25440 = ~l1484 & ~l1118;
assign a25442 = l1484 & l1118;
assign a25444 = ~a25442 & ~a25440;
assign a25446 = ~l1482 & l1116;
assign a25448 = l1482 & ~l1116;
assign a25450 = ~a25448 & ~a25446;
assign a25452 = ~l1488 & ~l1124;
assign a25454 = l1488 & l1124;
assign a25456 = ~a25454 & ~a25452;
assign a25458 = ~l1486 & l1122;
assign a25460 = l1486 & ~l1122;
assign a25462 = ~a25460 & ~a25458;
assign a25464 = ~l1492 & ~l1132;
assign a25466 = l1492 & l1132;
assign a25468 = ~a25466 & ~a25464;
assign a25470 = ~l1490 & l1130;
assign a25472 = l1490 & ~l1130;
assign a25474 = ~a25472 & ~a25470;
assign a25476 = ~l1496 & ~l1138;
assign a25478 = l1496 & l1138;
assign a25480 = ~a25478 & ~a25476;
assign a25482 = ~l1494 & l1136;
assign a25484 = l1494 & ~l1136;
assign a25486 = ~a25484 & ~a25482;
assign a25488 = ~l1500 & ~l1146;
assign a25490 = l1500 & l1146;
assign a25492 = ~a25490 & ~a25488;
assign a25494 = ~l1498 & l1144;
assign a25496 = l1498 & ~l1144;
assign a25498 = ~a25496 & ~a25494;
assign a25500 = ~l1504 & ~l1152;
assign a25502 = l1504 & l1152;
assign a25504 = ~a25502 & ~a25500;
assign a25506 = ~l1502 & l1150;
assign a25508 = l1502 & ~l1150;
assign a25510 = ~a25508 & ~a25506;
assign a25512 = ~l1510 & ~l1158;
assign a25514 = l1510 & l1158;
assign a25516 = ~a25514 & ~a25512;
assign a25518 = ~l1508 & l1156;
assign a25520 = l1508 & ~l1156;
assign a25522 = ~a25520 & ~a25518;
assign a25524 = ~l1506 & l1154;
assign a25526 = l1506 & ~l1154;
assign a25528 = ~a25526 & ~a25524;
assign a25530 = ~l1512 & l1160;
assign a25532 = l1512 & ~l1160;
assign a25534 = ~a25532 & ~a25530;
assign a25536 = ~l1516 & l1164;
assign a25538 = l1516 & ~l1164;
assign a25540 = ~a25538 & ~a25536;
assign a25542 = ~l1514 & l1162;
assign a25544 = l1514 & ~l1162;
assign a25546 = ~a25544 & ~a25542;
assign a25548 = ~l1518 & l1168;
assign a25550 = l1518 & ~l1168;
assign a25552 = ~a25550 & ~a25548;
assign a25554 = ~l1520 & l1170;
assign a25556 = l1520 & ~l1170;
assign a25558 = ~a25556 & ~a25554;
assign a25560 = ~l1530 & l1180;
assign a25562 = l1530 & ~l1180;
assign a25564 = ~a25562 & ~a25560;
assign a25566 = ~l1528 & l1178;
assign a25568 = l1528 & ~l1178;
assign a25570 = ~a25568 & ~a25566;
assign a25572 = ~l1526 & l1176;
assign a25574 = l1526 & ~l1176;
assign a25576 = ~a25574 & ~a25572;
assign a25578 = ~l1524 & l1174;
assign a25580 = l1524 & ~l1174;
assign a25582 = ~a25580 & ~a25578;
assign a25584 = ~l1522 & l1172;
assign a25586 = l1522 & ~l1172;
assign a25588 = ~a25586 & ~a25584;
assign a25590 = ~l1534 & ~l1188;
assign a25592 = l1534 & l1188;
assign a25594 = ~a25592 & ~a25590;
assign a25596 = ~l1532 & l1186;
assign a25598 = l1532 & ~l1186;
assign a25600 = ~a25598 & ~a25596;
assign a25602 = ~l1538 & ~l1194;
assign a25604 = l1538 & l1194;
assign a25606 = ~a25604 & ~a25602;
assign a25608 = ~l1536 & l1192;
assign a25610 = l1536 & ~l1192;
assign a25612 = ~a25610 & ~a25608;
assign a25614 = ~l1542 & ~l1202;
assign a25616 = l1542 & l1202;
assign a25618 = ~a25616 & ~a25614;
assign a25620 = ~l1540 & l1200;
assign a25622 = l1540 & ~l1200;
assign a25624 = ~a25622 & ~a25620;
assign a25626 = ~l1546 & ~l1208;
assign a25628 = l1546 & l1208;
assign a25630 = ~a25628 & ~a25626;
assign a25632 = ~l1544 & l1206;
assign a25634 = l1544 & ~l1206;
assign a25636 = ~a25634 & ~a25632;
assign a25638 = ~l1550 & ~l1216;
assign a25640 = l1550 & l1216;
assign a25642 = ~a25640 & ~a25638;
assign a25644 = ~l1548 & l1214;
assign a25646 = l1548 & ~l1214;
assign a25648 = ~a25646 & ~a25644;
assign a25650 = ~l1554 & ~l1222;
assign a25652 = l1554 & l1222;
assign a25654 = ~a25652 & ~a25650;
assign a25656 = ~l1552 & l1220;
assign a25658 = l1552 & ~l1220;
assign a25660 = ~a25658 & ~a25656;
assign a25662 = ~l1558 & ~l1230;
assign a25664 = l1558 & l1230;
assign a25666 = ~a25664 & ~a25662;
assign a25668 = ~l1556 & l1228;
assign a25670 = l1556 & ~l1228;
assign a25672 = ~a25670 & ~a25668;
assign a25674 = ~l1562 & ~l1236;
assign a25676 = l1562 & l1236;
assign a25678 = ~a25676 & ~a25674;
assign a25680 = ~l1560 & l1234;
assign a25682 = l1560 & ~l1234;
assign a25684 = ~a25682 & ~a25680;
assign a25686 = ~l1568 & ~l1242;
assign a25688 = l1568 & l1242;
assign a25690 = ~a25688 & ~a25686;
assign a25692 = ~l1566 & l1240;
assign a25694 = l1566 & ~l1240;
assign a25696 = ~a25694 & ~a25692;
assign a25698 = ~l1564 & l1238;
assign a25700 = l1564 & ~l1238;
assign a25702 = ~a25700 & ~a25698;
assign a25704 = ~l1570 & l1244;
assign a25706 = l1570 & ~l1244;
assign a25708 = ~a25706 & ~a25704;
assign a25710 = ~l1574 & l1248;
assign a25712 = l1574 & ~l1248;
assign a25714 = ~a25712 & ~a25710;
assign a25716 = ~l1572 & l1246;
assign a25718 = l1572 & ~l1246;
assign a25720 = ~a25718 & ~a25716;
assign a25722 = ~l1576 & l1252;
assign a25724 = l1576 & ~l1252;
assign a25726 = ~a25724 & ~a25722;
assign a25728 = ~l1578 & l1254;
assign a25730 = l1578 & ~l1254;
assign a25732 = ~a25730 & ~a25728;
assign a25734 = ~l1588 & l1264;
assign a25736 = l1588 & ~l1264;
assign a25738 = ~a25736 & ~a25734;
assign a25740 = ~l1586 & l1262;
assign a25742 = l1586 & ~l1262;
assign a25744 = ~a25742 & ~a25740;
assign a25746 = ~l1584 & l1260;
assign a25748 = l1584 & ~l1260;
assign a25750 = ~a25748 & ~a25746;
assign a25752 = ~l1582 & l1258;
assign a25754 = l1582 & ~l1258;
assign a25756 = ~a25754 & ~a25752;
assign a25758 = ~l1580 & l1256;
assign a25760 = l1580 & ~l1256;
assign a25762 = ~a25760 & ~a25758;
assign a25764 = ~l1592 & ~l1272;
assign a25766 = l1592 & l1272;
assign a25768 = ~a25766 & ~a25764;
assign a25770 = ~l1590 & l1270;
assign a25772 = l1590 & ~l1270;
assign a25774 = ~a25772 & ~a25770;
assign a25776 = ~l1596 & ~l1278;
assign a25778 = l1596 & l1278;
assign a25780 = ~a25778 & ~a25776;
assign a25782 = ~l1594 & l1276;
assign a25784 = l1594 & ~l1276;
assign a25786 = ~a25784 & ~a25782;
assign a25788 = ~l1600 & ~l1286;
assign a25790 = l1600 & l1286;
assign a25792 = ~a25790 & ~a25788;
assign a25794 = ~l1598 & l1284;
assign a25796 = l1598 & ~l1284;
assign a25798 = ~a25796 & ~a25794;
assign a25800 = ~l1604 & ~l1292;
assign a25802 = l1604 & l1292;
assign a25804 = ~a25802 & ~a25800;
assign a25806 = ~l1602 & l1290;
assign a25808 = l1602 & ~l1290;
assign a25810 = ~a25808 & ~a25806;
assign a25812 = ~l1608 & ~l1300;
assign a25814 = l1608 & l1300;
assign a25816 = ~a25814 & ~a25812;
assign a25818 = ~l1606 & l1298;
assign a25820 = l1606 & ~l1298;
assign a25822 = ~a25820 & ~a25818;
assign a25824 = ~l1612 & ~l1306;
assign a25826 = l1612 & l1306;
assign a25828 = ~a25826 & ~a25824;
assign a25830 = ~l1610 & l1304;
assign a25832 = l1610 & ~l1304;
assign a25834 = ~a25832 & ~a25830;
assign a25836 = ~l1616 & ~l1314;
assign a25838 = l1616 & l1314;
assign a25840 = ~a25838 & ~a25836;
assign a25842 = ~l1614 & l1312;
assign a25844 = l1614 & ~l1312;
assign a25846 = ~a25844 & ~a25842;
assign a25848 = ~l1620 & ~l1320;
assign a25850 = l1620 & l1320;
assign a25852 = ~a25850 & ~a25848;
assign a25854 = ~l1618 & l1318;
assign a25856 = l1618 & ~l1318;
assign a25858 = ~a25856 & ~a25854;
assign a25860 = ~l1624 & l1324;
assign a25862 = l1624 & ~l1324;
assign a25864 = ~a25862 & ~a25860;
assign a25866 = ~l1622 & l1322;
assign a25868 = l1622 & ~l1322;
assign a25870 = ~a25868 & ~a25866;
assign a25872 = ~l1628 & l1328;
assign a25874 = l1628 & ~l1328;
assign a25876 = ~a25874 & ~a25872;
assign a25878 = ~l1632 & l1332;
assign a25880 = l1632 & ~l1332;
assign a25882 = ~a25880 & ~a25878;
assign a25884 = ~l1630 & l1330;
assign a25886 = l1630 & ~l1330;
assign a25888 = ~a25886 & ~a25884;
assign a25890 = ~l1634 & l1336;
assign a25892 = l1634 & ~l1336;
assign a25894 = ~a25892 & ~a25890;
assign a25896 = ~l1636 & l1338;
assign a25898 = l1636 & ~l1338;
assign a25900 = ~a25898 & ~a25896;
assign a25902 = ~l1646 & l1348;
assign a25904 = l1646 & ~l1348;
assign a25906 = ~a25904 & ~a25902;
assign a25908 = ~l1644 & l1346;
assign a25910 = l1644 & ~l1346;
assign a25912 = ~a25910 & ~a25908;
assign a25914 = ~l1642 & l1344;
assign a25916 = l1642 & ~l1344;
assign a25918 = ~a25916 & ~a25914;
assign a25920 = ~l1640 & l1342;
assign a25922 = l1640 & ~l1342;
assign a25924 = ~a25922 & ~a25920;
assign a25926 = ~l1638 & l1340;
assign a25928 = l1638 & ~l1340;
assign a25930 = ~a25928 & ~a25926;
assign a25932 = ~l1648 & l1350;
assign a25934 = l1648 & ~l1350;
assign a25936 = ~a25934 & ~a25932;
assign a25938 = l1650 & ~l1352;
assign a25940 = ~l1650 & l1352;
assign a25942 = ~a25940 & ~a25938;
assign a25944 = l1652 & ~l1354;
assign a25946 = ~l1652 & l1354;
assign a25948 = ~a25946 & ~a25944;
assign a25950 = l1654 & ~l1356;
assign a25952 = ~l1654 & l1356;
assign a25954 = ~a25952 & ~a25950;
assign a25956 = a25954 & a25948;
assign a25958 = a25956 & a25942;
assign a25960 = a25958 & a25936;
assign a25962 = a25960 & a25930;
assign a25964 = a25962 & a25924;
assign a25966 = a25964 & a25918;
assign a25968 = a25966 & a25912;
assign a25970 = a25968 & a25906;
assign a25972 = a25970 & a25900;
assign a25974 = a25972 & a25894;
assign a25976 = a25974 & a25888;
assign a25978 = a25976 & a25882;
assign a25980 = a25978 & a25876;
assign a25982 = a25980 & a25870;
assign a25984 = a25982 & a25864;
assign a25986 = ~l1626 & ~l1326;
assign a25988 = l1626 & l1326;
assign a25990 = ~a25988 & ~a25986;
assign a25992 = a25990 & a25984;
assign a25994 = a25992 & a25858;
assign a25996 = a25994 & a25852;
assign a25998 = a25996 & a25846;
assign a26000 = a25998 & a25840;
assign a26002 = a26000 & a25834;
assign a26004 = a26002 & a25828;
assign a26006 = a26004 & a25822;
assign a26008 = a26006 & a25816;
assign a26010 = a26008 & a25810;
assign a26012 = a26010 & a25804;
assign a26014 = a26012 & a25798;
assign a26016 = a26014 & a25792;
assign a26018 = a26016 & a25786;
assign a26020 = a26018 & a25780;
assign a26022 = a26020 & a25774;
assign a26024 = a26022 & a25768;
assign a26026 = a26024 & a25762;
assign a26028 = a26026 & a25756;
assign a26030 = a26028 & a25750;
assign a26032 = a26030 & a25744;
assign a26034 = a26032 & a25738;
assign a26036 = a26034 & a25732;
assign a26038 = a26036 & a25726;
assign a26040 = a26038 & a25720;
assign a26042 = a26040 & a25714;
assign a26044 = a26042 & a25708;
assign a26046 = a26044 & a25702;
assign a26048 = a26046 & a25696;
assign a26050 = a26048 & a25690;
assign a26052 = a26050 & a25684;
assign a26054 = a26052 & a25678;
assign a26056 = a26054 & a25672;
assign a26058 = a26056 & a25666;
assign a26060 = a26058 & a25660;
assign a26062 = a26060 & a25654;
assign a26064 = a26062 & a25648;
assign a26066 = a26064 & a25642;
assign a26068 = a26066 & a25636;
assign a26070 = a26068 & a25630;
assign a26072 = a26070 & a25624;
assign a26074 = a26072 & a25618;
assign a26076 = a26074 & a25612;
assign a26078 = a26076 & a25606;
assign a26080 = a26078 & a25600;
assign a26082 = a26080 & a25594;
assign a26084 = a26082 & a25588;
assign a26086 = a26084 & a25582;
assign a26088 = a26086 & a25576;
assign a26090 = a26088 & a25570;
assign a26092 = a26090 & a25564;
assign a26094 = a26092 & a25558;
assign a26096 = a26094 & a25552;
assign a26098 = a26096 & a25546;
assign a26100 = a26098 & a25540;
assign a26102 = a26100 & a25534;
assign a26104 = a26102 & a25528;
assign a26106 = a26104 & a25522;
assign a26108 = a26106 & a25516;
assign a26110 = a26108 & a25510;
assign a26112 = a26110 & a25504;
assign a26114 = a26112 & a25498;
assign a26116 = a26114 & a25492;
assign a26118 = a26116 & a25486;
assign a26120 = a26118 & a25480;
assign a26122 = a26120 & a25474;
assign a26124 = a26122 & a25468;
assign a26126 = a26124 & a25462;
assign a26128 = a26126 & a25456;
assign a26130 = a26128 & a25450;
assign a26132 = a26130 & a25444;
assign a26134 = a26132 & a25438;
assign a26136 = a26134 & a25432;
assign a26138 = a26136 & a25426;
assign a26140 = a26138 & a25420;
assign a26142 = a26140 & a25414;
assign a26144 = a26142 & a25408;
assign a26146 = a26144 & a25402;
assign a26148 = a26146 & a25396;
assign a26150 = a26148 & a25390;
assign a26152 = a26150 & a25384;
assign a26154 = a26152 & a25378;
assign a26156 = a26154 & a25372;
assign a26158 = a26156 & a25366;
assign a26160 = a26158 & a25360;
assign a26162 = a26160 & a25354;
assign a26164 = a26162 & a25348;
assign a26166 = a26164 & a25342;
assign a26168 = a26166 & a25336;
assign a26170 = a26168 & a25330;
assign a26172 = a26170 & a25324;
assign a26174 = a26172 & a25318;
assign a26176 = a26174 & a25312;
assign a26178 = a26176 & a25306;
assign a26180 = a26178 & a25300;
assign a26182 = a26180 & a25294;
assign a26184 = a26182 & a25288;
assign a26186 = a26184 & a25282;
assign a26188 = a26186 & a25276;
assign a26190 = a26188 & a25270;
assign a26192 = a26190 & a25264;
assign a26194 = a26192 & a25258;
assign a26196 = a26194 & a25252;
assign a26198 = a26196 & a25246;
assign a26200 = a26198 & a25240;
assign a26202 = a26200 & a25234;
assign a26204 = a26202 & a25228;
assign a26206 = a26204 & a25222;
assign a26208 = a26206 & a25216;
assign a26210 = a26208 & a25210;
assign a26212 = a26210 & a25204;
assign a26214 = a26212 & a25198;
assign a26216 = a26214 & a25192;
assign a26218 = a26216 & a25186;
assign a26220 = a26218 & a25180;
assign a26222 = a26220 & a25174;
assign a26224 = a26222 & a25168;
assign a26226 = a26224 & a25162;
assign a26228 = a26226 & a25156;
assign a26230 = a26228 & a25150;
assign a26232 = a26230 & a25144;
assign a26234 = a26232 & a25138;
assign a26236 = a26234 & a25132;
assign a26238 = a26236 & a25126;
assign a26240 = a26238 & a25120;
assign a26242 = a26240 & a25114;
assign a26244 = a26242 & a25108;
assign a26246 = a26244 & a25102;
assign a26248 = a26246 & a25096;
assign a26250 = a26248 & a25090;
assign a26252 = a26250 & a25084;
assign a26254 = a26252 & a25078;
assign a26256 = a26254 & a25072;
assign a26258 = a26256 & l1664;
assign a26260 = a26258 & l1656;
assign a26262 = a26260 & l1658;
assign a26264 = a26262 & l1660;
assign a26266 = ~a26264 & i718;
assign a26268 = ~a26266 & a25066;
assign a26270 = a26268 & a25060;
assign a26272 = a26270 & a25054;
assign a26274 = a26272 & a25048;
assign a26276 = a26274 & a25042;
assign a26278 = a26276 & a25036;
assign a26280 = a26278 & a25030;
assign a26282 = a26280 & a25024;
assign a26284 = a26282 & a25018;
assign a26286 = a26284 & a25012;
assign a26288 = a26286 & a25006;
assign a26290 = a26288 & a25000;
assign a26292 = a26290 & a24994;
assign a26294 = a26292 & a24988;
assign a26296 = a26294 & a24982;
assign a26298 = a26296 & a24976;
assign a26300 = a26298 & a24970;
assign a26302 = a26300 & a24964;
assign a26304 = a26302 & a24958;
assign a26306 = a26304 & a24952;
assign a26308 = a26306 & ~a24946;
assign a26310 = a26308 & ~a24918;
assign a26312 = a26310 & ~a24890;
assign a26314 = a26312 & ~a24862;
assign a26316 = a26314 & ~a24834;
assign a26318 = a26316 & ~a24790;
assign a26320 = a26318 & ~a24746;
assign a26322 = a26320 & ~a24702;
assign a26324 = a26322 & ~a24622;
assign a26326 = a26324 & ~a24578;
assign a26328 = a26326 & ~a24534;
assign a26330 = a26328 & ~a24490;
assign a26332 = a26330 & ~a24410;
assign a26334 = a26332 & ~a24366;
assign a26336 = a26334 & ~a24322;
assign a26338 = a26336 & ~a24278;
assign a26340 = a26338 & ~a24198;
assign a26342 = a26340 & ~a24110;
assign a26344 = a26342 & ~a24022;
assign a26346 = a26344 & ~a23934;
assign a26348 = a26346 & ~a23810;
assign a26350 = a26348 & ~a23766;
assign a26352 = a26350 & ~a23722;
assign a26354 = a26352 & ~a23678;
assign a26356 = a26354 & ~a23598;
assign a26358 = a26356 & ~a23554;
assign a26360 = a26358 & ~a23510;
assign a26362 = a26360 & ~a23466;
assign a26364 = a26362 & ~a23382;
assign a26366 = a26364 & ~a23338;
assign a26368 = a26366 & ~a23294;
assign a26370 = a26368 & ~a23250;
assign a26372 = a26370 & ~a23166;
assign a26374 = a26372 & ~a23078;
assign a26376 = a26374 & ~a22990;
assign a26378 = a26376 & ~a22902;
assign a26380 = a26378 & ~a22774;
assign a26382 = a26380 & ~a22730;
assign a26384 = a26382 & ~a22686;
assign a26386 = a26384 & ~a22642;
assign a26388 = a26386 & ~a22562;
assign a26390 = a26388 & ~a22518;
assign a26392 = a26390 & ~a22474;
assign a26394 = a26392 & ~a22430;
assign a26396 = a26394 & ~a22342;
assign a26398 = a26396 & ~a22298;
assign a26400 = a26398 & ~a22254;
assign a26402 = a26400 & ~a22210;
assign a26404 = a26402 & ~a22116;
assign a26406 = a26404 & ~a22028;
assign a26408 = a26406 & ~a21940;
assign a26410 = a26408 & ~a21852;
assign a26412 = a26410 & ~a21714;
assign a26414 = a26412 & ~a21670;
assign a26416 = a26414 & ~a21626;
assign a26418 = a26416 & ~a21582;
assign a26420 = a26418 & ~a21502;
assign a26422 = a26420 & ~a21458;
assign a26424 = a26422 & ~a21414;
assign a26426 = a26424 & ~a21370;
assign a26428 = a26426 & ~a21282;
assign a26430 = a26428 & ~a21238;
assign a26432 = a26430 & ~a21194;
assign a26434 = a26432 & ~a21150;
assign a26436 = a26434 & ~a21036;
assign a26438 = a26436 & ~a20948;
assign a26440 = a26438 & ~a20860;
assign a26442 = a26440 & ~a20772;
assign a26444 = a26442 & ~a20618;
assign a26446 = a26444 & ~a20574;
assign a26448 = a26446 & ~a20530;
assign a26450 = a26448 & ~a20486;
assign a26452 = a26450 & ~a20406;
assign a26454 = a26452 & ~a20362;
assign a26456 = a26454 & ~a20318;
assign a26458 = a26456 & ~a20274;
assign a26460 = a26458 & ~a20186;
assign a26462 = a26460 & ~a20142;
assign a26464 = a26462 & ~a20098;
assign a26466 = a26464 & ~a20054;
assign a26468 = a26466 & ~a19940;
assign a26470 = a26468 & ~a19852;
assign a26472 = a26470 & ~a19764;
assign a26474 = a26472 & ~a19676;
assign a26476 = a26474 & a19474;
assign a26478 = a26476 & ~a15918;
assign a26480 = a26478 & a19310;
assign a26482 = a26480 & ~a15622;
assign a26484 = a26482 & a19146;
assign a26486 = a26484 & ~a15326;
assign a26488 = a26486 & a18982;
assign a26490 = a26488 & ~a15030;
assign a26492 = a26490 & a18818;
assign a26494 = a26492 & ~a14732;
assign a26496 = a26494 & a18654;
assign a26498 = a26496 & ~a14436;
assign a26500 = a26498 & a18490;
assign a26502 = a26500 & ~a14140;
assign a26504 = a26502 & a18326;
assign a26506 = a26504 & ~a13844;
assign a26508 = a26506 & a18162;
assign a26510 = a26508 & ~a13546;
assign a26512 = a26510 & a17998;
assign a26514 = a26512 & ~a13250;
assign a26516 = a26514 & a17834;
assign a26518 = a26516 & ~a12954;
assign a26520 = a26518 & a17670;
assign a26522 = a26520 & ~a12658;
assign a26524 = a26522 & a17506;
assign a26526 = a26524 & ~a12358;
assign a26528 = a26526 & a17342;
assign a26530 = a26528 & ~a12062;
assign a26532 = a26530 & a17178;
assign a26534 = a26532 & ~a11766;
assign a26536 = a26534 & a17014;
assign a26538 = a26536 & ~a11470;
assign a26540 = a26538 & a16850;
assign a26542 = a26540 & ~a11170;
assign a26544 = a26542 & a16686;
assign a26546 = a26544 & ~a10874;
assign a26548 = a26546 & a16522;
assign a26550 = a26548 & ~a10578;
assign a26552 = a26550 & a16358;
assign a26554 = a26552 & ~a10282;
assign a26556 = a26554 & ~a16194;
assign a26558 = a26556 & ~a15898;
assign a26560 = a26558 & ~a15602;
assign a26562 = a26560 & ~a15306;
assign a26564 = a26562 & ~a15010;
assign a26566 = a26564 & ~a14714;
assign a26568 = a26566 & ~a14418;
assign a26570 = a26568 & ~a14122;
assign a26572 = a26570 & ~a13826;
assign a26574 = a26572 & ~a13530;
assign a26576 = a26574 & ~a13234;
assign a26578 = a26576 & ~a12938;
assign a26580 = a26578 & ~a12642;
assign a26582 = a26580 & ~a12346;
assign a26584 = a26582 & ~a12050;
assign a26586 = a26584 & ~a11754;
assign a26588 = a26586 & ~a11458;
assign a26590 = a26588 & ~a11162;
assign a26592 = a26590 & ~a10866;
assign a26594 = a26592 & ~a10570;
assign a26596 = a26594 & ~a10274;
assign a26598 = a26596 & ~a10160;
assign a26600 = a26598 & ~a10152;
assign a26602 = a26600 & ~a10148;
assign a26604 = a26602 & ~a10146;
assign a26606 = a26604 & ~a10144;
assign a26608 = a26606 & ~a10142;
assign a26610 = a26608 & ~a10140;
assign a26612 = a26610 & ~a10132;
assign a26614 = a26612 & ~a10128;
assign a26616 = a26614 & ~a10126;
assign a26618 = a26616 & ~a10124;
assign a26620 = a26618 & ~a10122;
assign a26622 = a26620 & ~a10120;
assign a26624 = a26622 & ~a10112;
assign a26626 = a26624 & ~a10108;
assign a26628 = a26626 & ~a10106;
assign a26630 = a26628 & ~a10104;
assign a26632 = a26630 & ~a10102;
assign a26634 = a26632 & ~a10100;
assign a26636 = a26634 & ~a10092;
assign a26638 = a26636 & ~a10088;
assign a26640 = a26638 & ~a10086;
assign a26642 = a26640 & ~a10084;
assign a26644 = a26642 & ~a10082;
assign a26646 = a26644 & ~a10080;
assign a26648 = a26646 & ~a10072;
assign a26650 = a26648 & ~a10068;
assign a26652 = a26650 & ~a10066;
assign a26654 = a26652 & ~a10064;
assign a26656 = a26654 & ~a10062;
assign a26658 = a26656 & ~a10060;
assign a26660 = a26658 & ~a10056;
assign a26662 = a26660 & ~a10054;
assign a26664 = a26662 & ~a10052;
assign a26666 = a26664 & ~a10050;
assign a26668 = a26666 & ~a10048;
assign a26670 = a26668 & ~a10046;
assign a26672 = a26670 & ~a10044;
assign a26674 = a26672 & ~a10042;
assign a26676 = a26674 & ~a10040;
assign a26678 = a26676 & ~a10038;
assign a26680 = a26678 & ~a10034;
assign a26682 = a26680 & ~a10032;
assign a26684 = a26682 & ~a10030;
assign a26686 = a26684 & ~a10028;
assign a26688 = a26686 & ~a10026;
assign a26690 = a26688 & ~a10024;
assign a26692 = a26690 & ~a10022;
assign a26694 = a26692 & ~a10020;
assign a26696 = a26694 & ~a10018;
assign a26698 = a26696 & ~a10016;
assign a26700 = a26698 & ~a10012;
assign a26702 = a26700 & ~a10010;
assign a26704 = a26702 & ~a10008;
assign a26706 = a26704 & ~a10006;
assign a26708 = a26706 & ~a10004;
assign a26710 = a26708 & ~a10002;
assign a26712 = a26710 & ~a10000;
assign a26714 = a26712 & ~a9998;
assign a26716 = a26714 & ~a9996;
assign a26718 = a26716 & ~a9994;
assign a26720 = a26718 & ~a9990;
assign a26722 = a26720 & ~a9988;
assign a26724 = a26722 & ~a9986;
assign a26726 = a26724 & ~a9984;
assign a26728 = a26726 & ~a9982;
assign a26730 = a26728 & ~a9980;
assign a26732 = a26730 & ~a9978;
assign a26734 = a26732 & ~a9976;
assign a26736 = a26734 & ~a9974;
assign a26738 = a26736 & ~a9972;
assign a26740 = a26738 & ~a9968;
assign a26742 = a26740 & ~a9966;
assign a26744 = a26742 & ~a9964;
assign a26746 = a26744 & ~a9962;
assign a26748 = a26746 & ~a9960;
assign a26750 = a26748 & ~a9958;
assign a26752 = a26750 & ~a9956;
assign a26754 = a26752 & ~a9954;
assign a26756 = a26754 & ~a9952;
assign a26758 = a26756 & ~a9950;
assign a26760 = a26758 & ~a9948;
assign a26762 = a26760 & ~a9946;
assign a26764 = a26762 & ~a9944;
assign a26766 = a26764 & ~a9942;
assign a26768 = a26766 & ~a9940;
assign a26770 = a26768 & ~a9938;
assign a26772 = a26770 & ~a9936;
assign a26774 = a26772 & ~a9934;
assign a26776 = a26774 & ~a9932;
assign a26778 = a26776 & ~a9930;
assign a26780 = a26778 & ~a9928;
assign a26782 = a26780 & ~a9926;
assign a26784 = a26782 & ~a9924;
assign a26786 = a26784 & ~a9922;
assign a26788 = a26786 & ~a9920;
assign a26790 = a26788 & ~a9918;
assign a26792 = a26790 & ~a9916;
assign a26794 = a26792 & ~a9914;
assign a26796 = a26794 & ~a9912;
assign a26798 = a26796 & l1676;
assign a26800 = a26798 & a9910;
assign a26804 = a26798 & i718;
assign p0 = a26804;

assert property (~p0);

endmodule
