module m6s18 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76;

output p0;

wire na854,na882,na900,na912,na934,na952,na970,na876,na964,na946,na928,na906,a894,na978,na1380,
na1396,na1408,na1390,na1402,na1420,na1448,na1466,na1484,na1502,na1520,na1538,na1556,na1574,na1606,na1618,
na1630,na1654,na1706,na1720,na1754,na1776,na1794,na1812,na1830,na1848,na1866,na1882,na1894,na1912,na1948,
na1988,na2004,na2016,na2034,na2078,na2090,na2108,na2126,na2142,na2160,na2172,na2194,na2210,na2222,na2238,
na2250,na2268,na2286,na2304,na1374,na2298,na2280,na2262,na2244,na2318,na2232,na2312,na2216,na2332,na2204,
na2346,na2360,na2326,na2354,na2340,na2188,na2166,na2154,na2136,na2378,na2400,na2120,na2394,na2418,na2372,
na2412,na2102,na2084,na2442,na2454,na2466,na2478,na2490,na2502,na2520,na2536,na2072,na2530,na2514,na2548,
na2496,na2560,na2542,na2572,na2554,na2584,na2566,na2596,na2578,na2608,na2590,na2622,na2602,na2634,na2616,
na2646,na2628,na2658,na2640,na2670,na2652,na2664,na2484,na2472,na2460,na2448,na2436,na2028,na2010,na2688,
na1998,na2710,na2682,na2704,na2760,na2790,na2816,na2836,na1982,na2830,na2848,na2810,na2842,na2784,na2754,
na1942,na1906,na1888,na1876,na1860,na1842,na1824,na1806,na1788,na2898,na2924,na2950,na2972,na2990,na3012,
na3034,na3056,na3078,na1770,na3072,na3050,na3028,na3006,na2984,na2966,na2944,na2918,na2892,na1748,na1714,
na1700,na1648,na1624,na1612,na1600,na1568,na1550,na1532,na1514,na1496,na1478,na1460,na1442,na1414,na972,
na3096,na3114,na3132,na3150,na848,na3144,na3126,na3108,a3090,na3156,na3530,na3546,na3550,na3540,na3562,
na3580,na3598,na3616,na3634,na3652,na3670,na3688,na3706,na3734,na3746,na3796,na3808,na3832,na3872,na3884,
na3902,na3920,na3938,na3956,na3974,na3992,na4008,na4042,na4076,na4092,na4098,na4116,na4156,na4168,na4186,
na4202,na4220,na4232,na4254,na4270,na4276,na4292,na4298,na4316,na4334,na4352,na3524,na4346,na4328,na4310,
na4366,na4286,na4360,na4380,na4264,na4394,na4408,na4374,na4402,na4388,na4248,na4226,na4214,na4196,na4426,
na4448,na4180,na4442,na4466,na4420,na4460,na4162,na4472,na4488,na4494,na4500,na4506,na4518,na4538,na4556,
na4150,na4550,na4532,na4568,na4512,na4580,na4562,na4592,na4574,na4604,na4586,na4616,na4598,na4628,na4610,
na4640,na4622,na4652,na4634,na4664,na4646,na4676,na4658,na4688,na4670,na4682,na4482,na4110,na4706,na4086,
na4728,na4700,na4722,na4770,na4798,na4824,na4844,na4070,na4838,na4850,na4818,na4792,na4764,na4036,na4002,
na3986,na3968,na3950,na3932,na3914,na4900,na4926,na4952,na4974,na4992,na5014,na5036,na5058,na5080,na3896,
na5074,na5052,na5030,na5008,na4986,na4968,na4946,na4920,na4894,na3878,na3866,na3826,na3802,na3790,na3740,
na3728,na3700,na3682,na3664,na3646,na3628,na3610,na3592,na3574,na3556,c1,a822,a824,a826,a828,
a830,a832,a834,a836,a838,a840,a842,a844,a846,a848,a850,a852,a854,a856,a858,
a860,a862,a864,a866,a868,a870,a872,a874,a876,a878,a880,a882,a884,a886,a888,
a890,a892,a896,a898,a900,a902,a904,a906,a908,a910,a912,a914,a916,a918,a920,
a922,a924,a926,a928,a930,a932,a934,a936,a938,a940,a942,a944,a946,a948,a950,
a952,a954,a956,a958,a960,a962,a964,a966,a968,a970,a972,a974,a976,a978,a980,
a982,a984,a986,a988,a990,a992,a994,a996,a998,a1000,a1002,a1004,a1006,a1008,a1010,
a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,a1038,a1040,
a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,a1062,a1064,a1066,a1068,a1070,
a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,a1092,a1094,a1096,a1098,a1100,
a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,a1124,a1126,a1128,a1130,
a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,a1154,a1156,a1158,a1160,
a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,a1178,a1180,a1182,a1184,a1186,a1188,a1190,
a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,a1218,a1220,
a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,a1248,a1250,
a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,a1268,a1270,a1272,a1274,a1276,a1278,a1280,
a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,a1310,
a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,a1334,a1336,a1338,a1340,
a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,a1368,a1370,
a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,a1388,a1390,a1392,a1394,a1396,a1398,a1400,
a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1426,a1428,a1430,
a1432,a1434,a1436,a1438,a1440,a1442,a1444,a1446,a1448,a1450,a1452,a1454,a1456,a1458,a1460,
a1462,a1464,a1466,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1482,a1484,a1486,a1488,a1490,
a1492,a1494,a1496,a1498,a1500,a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,a1518,a1520,
a1522,a1524,a1526,a1528,a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,a1548,a1550,
a1552,a1554,a1556,a1558,a1560,a1562,a1564,a1566,a1568,a1570,a1572,a1574,a1576,a1578,a1580,
a1582,a1584,a1586,a1588,a1590,a1592,a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,a1610,
a1612,a1614,a1616,a1618,a1620,a1622,a1624,a1626,a1628,a1630,a1632,a1634,a1636,a1638,a1640,
a1642,a1644,a1646,a1648,a1650,a1652,a1654,a1656,a1658,a1660,a1662,a1664,a1666,a1668,a1670,
a1672,a1674,a1676,a1678,a1680,a1682,a1684,a1686,a1688,a1690,a1692,a1694,a1696,a1698,a1700,
a1702,a1704,a1706,a1708,a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,
a1732,a1734,a1736,a1738,a1740,a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,a1758,a1760,
a1762,a1764,a1766,a1768,a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,a1790,
a1792,a1794,a1796,a1798,a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,
a1822,a1824,a1826,a1828,a1830,a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,a1848,a1850,
a1852,a1854,a1856,a1858,a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,
a1882,a1884,a1886,a1888,a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,a1910,
a1912,a1914,a1916,a1918,a1920,a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,a1938,a1940,
a1942,a1944,a1946,a1948,a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,
a1972,a1974,a1976,a1978,a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,a1998,a2000,
a2002,a2004,a2006,a2008,a2010,a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,a2030,
a2032,a2034,a2036,a2038,a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,a2058,a2060,
a2062,a2064,a2066,a2068,a2070,a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,a2090,
a2092,a2094,a2096,a2098,a2100,a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,a2120,
a2122,a2124,a2126,a2128,a2130,a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,
a2152,a2154,a2156,a2158,a2160,a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,a2178,a2180,
a2182,a2184,a2186,a2188,a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,a2208,a2210,
a2212,a2214,a2216,a2218,a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,a2238,a2240,
a2242,a2244,a2246,a2248,a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,a2268,a2270,
a2272,a2274,a2276,a2278,a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,a2298,a2300,
a2302,a2304,a2306,a2308,a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,a2328,a2330,
a2332,a2334,a2336,a2338,a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,a2358,a2360,
a2362,a2364,a2366,a2368,a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,a2388,a2390,
a2392,a2394,a2396,a2398,a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,a2420,
a2422,a2424,a2426,a2428,a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,a2448,a2450,
a2452,a2454,a2456,a2458,a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,a2478,a2480,
a2482,a2484,a2486,a2488,a2490,a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,a2508,a2510,
a2512,a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,a2540,
a2542,a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,
a2572,a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,
a2602,a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,a2630,
a2632,a2634,a2636,a2638,a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,
a2662,a2664,a2666,a2668,a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,
a2692,a2694,a2696,a2698,a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,a2718,a2720,
a2722,a2724,a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,
a2752,a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,
a2782,a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,a2810,
a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,a2840,
a2842,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,a2870,
a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,a2900,
a2902,a2904,a2906,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2930,
a2932,a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,a2960,
a2962,a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,a2988,a2990,
a2992,a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,
a3022,a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,a3048,a3050,
a3052,a3054,a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,a3078,a3080,
a3082,a3084,a3086,a3088,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,a3112,
a3114,a3116,a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,a3142,
a3144,a3146,a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,a3172,
a3174,a3176,a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3200,a3202,
a3204,a3206,a3208,a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,a3228,a3230,a3232,
a3234,a3236,a3238,a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,a3262,
a3264,a3266,a3268,a3270,a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,a3288,a3290,a3292,
a3294,a3296,a3298,a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,
a3324,a3326,a3328,a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,
a3354,a3356,a3358,a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3382,
a3384,a3386,a3388,a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,a3408,a3410,a3412,
a3414,a3416,a3418,a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,a3438,a3440,a3442,
a3444,a3446,a3448,a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,a3468,a3470,a3472,
a3474,a3476,a3478,a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,a3498,a3500,a3502,
a3504,a3506,a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,a3528,a3530,a3532,
a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,a3558,a3560,a3562,
a3564,a3566,a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,a3588,a3590,a3592,
a3594,a3596,a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,a3618,a3620,a3622,
a3624,a3626,a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3648,a3650,a3652,
a3654,a3656,a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,a3678,a3680,a3682,
a3684,a3686,a3688,a3690,a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,a3712,
a3714,a3716,a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,a3738,a3740,a3742,
a3744,a3746,a3748,a3750,a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,a3768,a3770,a3772,
a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,a3798,a3800,a3802,
a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,a3828,a3830,a3832,
a3834,a3836,a3838,a3840,a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,a3858,a3860,a3862,
a3864,a3866,a3868,a3870,a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,a3888,a3890,a3892,
a3894,a3896,a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,a3918,a3920,a3922,
a3924,a3926,a3928,a3930,a3932,a3934,a3936,a3938,a3940,a3942,a3944,a3946,a3948,a3950,a3952,
a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,a3978,a3980,a3982,
a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,a4008,a4010,a4012,
a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,a4038,a4040,a4042,
a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,a4068,a4070,a4072,
a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,a4096,a4098,a4100,a4102,
a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4124,a4126,a4128,a4130,a4132,
a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,a4152,a4154,a4156,a4158,a4160,a4162,
a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,a4184,a4186,a4188,a4190,a4192,
a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,a4214,a4216,a4218,a4220,a4222,
a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,a4244,a4246,a4248,a4250,a4252,
a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,a4274,a4276,a4278,a4280,a4282,
a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,a4306,a4308,a4310,a4312,
a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,a4334,a4336,a4338,a4340,a4342,
a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,a4368,a4370,a4372,
a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,a4394,a4396,a4398,a4400,a4402,
a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,a4432,
a4434,a4436,a4438,a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,a4458,a4460,a4462,
a4464,a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4482,a4484,a4486,a4488,a4490,a4492,
a4494,a4496,a4498,a4500,a4502,a4504,a4506,a4508,a4510,a4512,a4514,a4516,a4518,a4520,a4522,
a4524,a4526,a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,
a4554,a4556,a4558,a4560,a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,a4578,a4580,a4582,
a4584,a4586,a4588,a4590,a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,a4612,
a4614,a4616,a4618,a4620,a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,a4642,
a4644,a4646,a4648,a4650,a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,a4672,
a4674,a4676,a4678,a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,a4696,a4698,a4700,a4702,
a4704,a4706,a4708,a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,a4726,a4728,a4730,a4732,
a4734,a4736,a4738,a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,a4756,a4758,a4760,a4762,
a4764,a4766,a4768,a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4784,a4786,a4788,a4790,a4792,
a4794,a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,a4818,a4820,a4822,
a4824,a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,a4844,a4846,a4848,a4850,a4852,
a4854,a4856,a4858,a4860,a4862,a4864,a4866,a4868,a4870,a4872,a4874,a4876,a4878,a4880,a4882,
a4884,a4886,a4888,a4890,a4892,a4894,a4896,a4898,a4900,a4902,a4904,a4906,a4908,a4910,a4912,
a4914,a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,a4938,a4940,a4942,
a4944,a4946,a4948,a4950,a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,a4968,a4970,a4972,
a4974,a4976,a4978,a4980,a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,a4998,a5000,a5002,
a5004,a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,a5028,a5030,a5032,
a5034,a5036,a5038,a5040,a5042,a5044,a5046,a5048,a5050,a5052,a5054,a5056,a5058,a5060,a5062,
a5064,a5066,a5068,a5070,a5072,a5074,a5076,a5078,a5080,p0;

reg l78,l80,l82,l84,l86,l88,l90,l92,l94,l96,l98,l100,l102,l104,l106,
l108,l110,l112,l114,l116,l118,l120,l122,l124,l126,l128,l130,l132,l134,l136,
l138,l140,l142,l144,l146,l148,l150,l152,l154,l156,l158,l160,l162,l164,l166,
l168,l170,l172,l174,l176,l178,l180,l182,l184,l186,l188,l190,l192,l194,l196,
l198,l200,l202,l204,l206,l208,l210,l212,l214,l216,l218,l220,l222,l224,l226,
l228,l230,l232,l234,l236,l238,l240,l242,l244,l246,l248,l250,l252,l254,l256,
l258,l260,l262,l264,l266,l268,l270,l272,l274,l276,l278,l280,l282,l284,l286,
l288,l290,l292,l294,l296,l298,l300,l302,l304,l306,l308,l310,l312,l314,l316,
l318,l320,l322,l324,l326,l328,l330,l332,l334,l336,l338,l340,l342,l344,l346,
l348,l350,l352,l354,l356,l358,l360,l362,l364,l366,l368,l370,l372,l374,l376,
l378,l380,l382,l384,l386,l388,l390,l392,l394,l396,l398,l400,l402,l404,l406,
l408,l410,l412,l414,l416,l418,l420,l422,l424,l426,l428,l430,l432,l434,l436,
l438,l440,l442,l444,l446,l448,l450,l452,l454,l456,l458,l460,l462,l464,l466,
l468,l470,l472,l474,l476,l478,l480,l482,l484,l486,l488,l490,l492,l494,l496,
l498,l500,l502,l504,l506,l508,l510,l512,l514,l516,l518,l520,l522,l524,l526,
l528,l530,l532,l534,l536,l538,l540,l542,l544,l546,l548,l550,l552,l554,l556,
l558,l560,l562,l564,l566,l568,l570,l572,l574,l576,l578,l580,l582,l584,l586,
l588,l590,l592,l594,l596,l598,l600,l602,l604,l606,l608,l610,l612,l614,l616,
l618,l620,l622,l624,l626,l628,l630,l632,l634,l636,l638,l640,l642,l644,l646,
l648,l650,l652,l654,l656,l658,l660,l662,l664,l666,l668,l670,l672,l674,l676,
l678,l680,l682,l684,l686,l688,l690,l692,l694,l696,l698,l700,l702,l704,l706,
l708,l710,l712,l714,l716,l718,l720,l722,l724,l726,l728,l730,l732,l734,l736,
l738,l740,l742,l744,l746,l748,l750,l752,l754,l756,l758,l760,l762,l764,l766,
l768,l770,l772,l774,l776,l778,l780,l782,l784,l786,l788,l790,l792,l794,l796,
l798,l800,l802,l804,l806,l808,l810,l812,l814,l816,l818,l820;

initial
begin
   l78 = 0;
   l80 = 0;
   l82 = 0;
   l84 = 0;
   l86 = 0;
   l88 = 0;
   l90 = 0;
   l92 = 0;
   l94 = 0;
   l96 = 0;
   l98 = 0;
   l100 = 0;
   l102 = 0;
   l104 = 0;
   l106 = 0;
   l108 = 0;
   l110 = 0;
   l112 = 0;
   l114 = 0;
   l116 = 0;
   l118 = 0;
   l120 = 0;
   l122 = 0;
   l124 = 0;
   l126 = 0;
   l128 = 0;
   l130 = 0;
   l132 = 0;
   l134 = 0;
   l136 = 0;
   l138 = 0;
   l140 = 0;
   l142 = 0;
   l144 = 0;
   l146 = 0;
   l148 = 0;
   l150 = 0;
   l152 = 0;
   l154 = 0;
   l156 = 0;
   l158 = 0;
   l160 = 0;
   l162 = 0;
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 0;
   l176 = 0;
   l178 = 0;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
   l392 = 0;
   l394 = 0;
   l396 = 0;
   l398 = 0;
   l400 = 0;
   l402 = 0;
   l404 = 0;
   l406 = 0;
   l408 = 0;
   l410 = 0;
   l412 = 0;
   l414 = 0;
   l416 = 0;
   l418 = 0;
   l420 = 0;
   l422 = 0;
   l424 = 0;
   l426 = 0;
   l428 = 0;
   l430 = 0;
   l432 = 0;
   l434 = 0;
   l436 = 0;
   l438 = 0;
   l440 = 0;
   l442 = 0;
   l444 = 0;
   l446 = 0;
   l448 = 0;
   l450 = 0;
   l452 = 0;
   l454 = 0;
   l456 = 0;
   l458 = 0;
   l460 = 0;
   l462 = 0;
   l464 = 0;
   l466 = 0;
   l468 = 0;
   l470 = 0;
   l472 = 0;
   l474 = 0;
   l476 = 0;
   l478 = 0;
   l480 = 0;
   l482 = 0;
   l484 = 0;
   l486 = 0;
   l488 = 0;
   l490 = 0;
   l492 = 0;
   l494 = 0;
   l496 = 0;
   l498 = 0;
   l500 = 0;
   l502 = 0;
   l504 = 0;
   l506 = 0;
   l508 = 0;
   l510 = 0;
   l512 = 0;
   l514 = 0;
   l516 = 0;
   l518 = 0;
   l520 = 0;
   l522 = 0;
   l524 = 0;
   l526 = 0;
   l528 = 0;
   l530 = 0;
   l532 = 0;
   l534 = 0;
   l536 = 0;
   l538 = 0;
   l540 = 0;
   l542 = 0;
   l544 = 0;
   l546 = 0;
   l548 = 0;
   l550 = 0;
   l552 = 0;
   l554 = 0;
   l556 = 0;
   l558 = 0;
   l560 = 0;
   l562 = 0;
   l564 = 0;
   l566 = 0;
   l568 = 0;
   l570 = 0;
   l572 = 0;
   l574 = 0;
   l576 = 0;
   l578 = 0;
   l580 = 0;
   l582 = 0;
   l584 = 0;
   l586 = 0;
   l588 = 0;
   l590 = 0;
   l592 = 0;
   l594 = 0;
   l596 = 0;
   l598 = 0;
   l600 = 0;
   l602 = 0;
   l604 = 0;
   l606 = 0;
   l608 = 0;
   l610 = 0;
   l612 = 0;
   l614 = 0;
   l616 = 0;
   l618 = 0;
   l620 = 0;
   l622 = 0;
   l624 = 0;
   l626 = 0;
   l628 = 0;
   l630 = 0;
   l632 = 0;
   l634 = 0;
   l636 = 0;
   l638 = 0;
   l640 = 0;
   l642 = 0;
   l644 = 0;
   l646 = 0;
   l648 = 0;
   l650 = 0;
   l652 = 0;
   l654 = 0;
   l656 = 0;
   l658 = 0;
   l660 = 0;
   l662 = 0;
   l664 = 0;
   l666 = 0;
   l668 = 0;
   l670 = 0;
   l672 = 0;
   l674 = 0;
   l676 = 0;
   l678 = 0;
   l680 = 0;
   l682 = 0;
   l684 = 0;
   l686 = 0;
   l688 = 0;
   l690 = 0;
   l692 = 0;
   l694 = 0;
   l696 = 0;
   l698 = 0;
   l700 = 0;
   l702 = 0;
   l704 = 0;
   l706 = 0;
   l708 = 0;
   l710 = 0;
   l712 = 0;
   l714 = 0;
   l716 = 0;
   l718 = 0;
   l720 = 0;
   l722 = 0;
   l724 = 0;
   l726 = 0;
   l728 = 0;
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
   l802 = 0;
   l804 = 0;
   l806 = 0;
   l808 = 0;
   l810 = 0;
   l812 = 0;
   l814 = 0;
   l816 = 0;
   l818 = 0;
   l820 = 0;
end

always @(posedge na854)
   l78 <= na854;

always @(posedge na882)
   l80 <= na882;

always @(posedge na900)
   l82 <= na900;

always @(posedge na912)
   l84 <= na912;

always @(posedge i2)
   l86 <= i2;

always @(posedge na934)
   l88 <= na934;

always @(posedge na952)
   l90 <= na952;

always @(posedge na970)
   l92 <= na970;

always @(posedge na876)
   l94 <= na876;

always @(posedge na964)
   l96 <= na964;

always @(posedge na946)
   l98 <= na946;

always @(posedge na928)
   l100 <= na928;

always @(posedge na906)
   l102 <= na906;

always @(posedge a894)
   l104 <= a894;

always @(posedge na978)
   l106 <= na978;

always @(posedge na1380)
   l108 <= na1380;

always @(posedge na1396)
   l110 <= na1396;

always @(posedge na1408)
   l112 <= na1408;

always @(posedge na1390)
   l114 <= na1390;

always @(posedge na1402)
   l116 <= na1402;

always @(posedge na1420)
   l118 <= na1420;

always @(posedge na1448)
   l120 <= na1448;

always @(posedge na1466)
   l122 <= na1466;

always @(posedge na1484)
   l124 <= na1484;

always @(posedge na1502)
   l126 <= na1502;

always @(posedge na1520)
   l128 <= na1520;

always @(posedge na1538)
   l130 <= na1538;

always @(posedge na1556)
   l132 <= na1556;

always @(posedge na1574)
   l134 <= na1574;

always @(posedge na1606)
   l136 <= na1606;

always @(posedge na1618)
   l138 <= na1618;

always @(posedge na1630)
   l140 <= na1630;

always @(posedge na1654)
   l142 <= na1654;

always @(posedge na1706)
   l144 <= na1706;

always @(posedge na1720)
   l146 <= na1720;

always @(posedge na1754)
   l148 <= na1754;

always @(posedge na1776)
   l150 <= na1776;

always @(posedge na1794)
   l152 <= na1794;

always @(posedge na1812)
   l154 <= na1812;

always @(posedge na1830)
   l156 <= na1830;

always @(posedge na1848)
   l158 <= na1848;

always @(posedge na1866)
   l160 <= na1866;

always @(posedge na1882)
   l162 <= na1882;

always @(posedge na1894)
   l164 <= na1894;

always @(posedge na1912)
   l166 <= na1912;

always @(posedge na1948)
   l168 <= na1948;

always @(posedge na1988)
   l170 <= na1988;

always @(posedge na2004)
   l172 <= na2004;

always @(posedge na2016)
   l174 <= na2016;

always @(posedge na2034)
   l176 <= na2034;

always @(posedge na2078)
   l178 <= na2078;

always @(posedge na2090)
   l180 <= na2090;

always @(posedge na2108)
   l182 <= na2108;

always @(posedge na2126)
   l184 <= na2126;

always @(posedge na2142)
   l186 <= na2142;

always @(posedge na2160)
   l188 <= na2160;

always @(posedge na2172)
   l190 <= na2172;

always @(posedge na2194)
   l192 <= na2194;

always @(posedge na2210)
   l194 <= na2210;

always @(posedge na2222)
   l196 <= na2222;

always @(posedge na2238)
   l198 <= na2238;

always @(posedge na2250)
   l200 <= na2250;

always @(posedge na2268)
   l202 <= na2268;

always @(posedge na2286)
   l204 <= na2286;

always @(posedge na2304)
   l206 <= na2304;

always @(posedge na1374)
   l208 <= na1374;

always @(posedge na2298)
   l210 <= na2298;

always @(posedge na2280)
   l212 <= na2280;

always @(posedge na2262)
   l214 <= na2262;

always @(posedge na2244)
   l216 <= na2244;

always @(posedge na2318)
   l218 <= na2318;

always @(posedge na2232)
   l220 <= na2232;

always @(posedge na2312)
   l222 <= na2312;

always @(posedge na2216)
   l224 <= na2216;

always @(posedge na2332)
   l226 <= na2332;

always @(posedge na2204)
   l228 <= na2204;

always @(posedge na2346)
   l230 <= na2346;

always @(posedge na2360)
   l232 <= na2360;

always @(posedge na2326)
   l234 <= na2326;

always @(posedge na2354)
   l236 <= na2354;

always @(posedge na2340)
   l238 <= na2340;

always @(posedge na2188)
   l240 <= na2188;

always @(posedge na2166)
   l242 <= na2166;

always @(posedge na2154)
   l244 <= na2154;

always @(posedge na2136)
   l246 <= na2136;

always @(posedge na2378)
   l248 <= na2378;

always @(posedge na2400)
   l250 <= na2400;

always @(posedge na2120)
   l252 <= na2120;

always @(posedge na2394)
   l254 <= na2394;

always @(posedge na2418)
   l256 <= na2418;

always @(posedge na2372)
   l258 <= na2372;

always @(posedge na2412)
   l260 <= na2412;

always @(posedge na2102)
   l262 <= na2102;

always @(posedge na2084)
   l264 <= na2084;

always @(posedge na2442)
   l266 <= na2442;

always @(posedge na2454)
   l268 <= na2454;

always @(posedge na2466)
   l270 <= na2466;

always @(posedge na2478)
   l272 <= na2478;

always @(posedge na2490)
   l274 <= na2490;

always @(posedge na2502)
   l276 <= na2502;

always @(posedge na2520)
   l278 <= na2520;

always @(posedge na2536)
   l280 <= na2536;

always @(posedge na2072)
   l282 <= na2072;

always @(posedge na2530)
   l284 <= na2530;

always @(posedge na2514)
   l286 <= na2514;

always @(posedge na2548)
   l288 <= na2548;

always @(posedge na2496)
   l290 <= na2496;

always @(posedge na2560)
   l292 <= na2560;

always @(posedge na2542)
   l294 <= na2542;

always @(posedge na2572)
   l296 <= na2572;

always @(posedge na2554)
   l298 <= na2554;

always @(posedge na2584)
   l300 <= na2584;

always @(posedge na2566)
   l302 <= na2566;

always @(posedge na2596)
   l304 <= na2596;

always @(posedge na2578)
   l306 <= na2578;

always @(posedge na2608)
   l308 <= na2608;

always @(posedge na2590)
   l310 <= na2590;

always @(posedge na2622)
   l312 <= na2622;

always @(posedge na2602)
   l314 <= na2602;

always @(posedge na2634)
   l316 <= na2634;

always @(posedge na2616)
   l318 <= na2616;

always @(posedge na2646)
   l320 <= na2646;

always @(posedge na2628)
   l322 <= na2628;

always @(posedge na2658)
   l324 <= na2658;

always @(posedge na2640)
   l326 <= na2640;

always @(posedge na2670)
   l328 <= na2670;

always @(posedge na2652)
   l330 <= na2652;

always @(posedge na2664)
   l332 <= na2664;

always @(posedge na2484)
   l334 <= na2484;

always @(posedge na2472)
   l336 <= na2472;

always @(posedge na2460)
   l338 <= na2460;

always @(posedge na2448)
   l340 <= na2448;

always @(posedge na2436)
   l342 <= na2436;

always @(posedge na2028)
   l344 <= na2028;

always @(posedge na2010)
   l346 <= na2010;

always @(posedge na2688)
   l348 <= na2688;

always @(posedge na1998)
   l350 <= na1998;

always @(posedge na2710)
   l352 <= na2710;

always @(posedge na2682)
   l354 <= na2682;

always @(posedge na2704)
   l356 <= na2704;

always @(posedge na2760)
   l358 <= na2760;

always @(posedge na2790)
   l360 <= na2790;

always @(posedge na2816)
   l362 <= na2816;

always @(posedge na2836)
   l364 <= na2836;

always @(posedge na1982)
   l366 <= na1982;

always @(posedge na2830)
   l368 <= na2830;

always @(posedge na2848)
   l370 <= na2848;

always @(posedge na2810)
   l372 <= na2810;

always @(posedge na2842)
   l374 <= na2842;

always @(posedge na2784)
   l376 <= na2784;

always @(posedge na2754)
   l378 <= na2754;

always @(posedge na1942)
   l380 <= na1942;

always @(posedge na1906)
   l382 <= na1906;

always @(posedge na1888)
   l384 <= na1888;

always @(posedge na1876)
   l386 <= na1876;

always @(posedge na1860)
   l388 <= na1860;

always @(posedge na1842)
   l390 <= na1842;

always @(posedge na1824)
   l392 <= na1824;

always @(posedge na1806)
   l394 <= na1806;

always @(posedge na1788)
   l396 <= na1788;

always @(posedge na2898)
   l398 <= na2898;

always @(posedge na2924)
   l400 <= na2924;

always @(posedge na2950)
   l402 <= na2950;

always @(posedge na2972)
   l404 <= na2972;

always @(posedge na2990)
   l406 <= na2990;

always @(posedge na3012)
   l408 <= na3012;

always @(posedge na3034)
   l410 <= na3034;

always @(posedge na3056)
   l412 <= na3056;

always @(posedge na3078)
   l414 <= na3078;

always @(posedge na1770)
   l416 <= na1770;

always @(posedge na3072)
   l418 <= na3072;

always @(posedge na3050)
   l420 <= na3050;

always @(posedge na3028)
   l422 <= na3028;

always @(posedge na3006)
   l424 <= na3006;

always @(posedge na2984)
   l426 <= na2984;

always @(posedge na2966)
   l428 <= na2966;

always @(posedge na2944)
   l430 <= na2944;

always @(posedge na2918)
   l432 <= na2918;

always @(posedge na2892)
   l434 <= na2892;

always @(posedge na1748)
   l436 <= na1748;

always @(posedge na1714)
   l438 <= na1714;

always @(posedge na1700)
   l440 <= na1700;

always @(posedge na1648)
   l442 <= na1648;

always @(posedge na1624)
   l444 <= na1624;

always @(posedge na1612)
   l446 <= na1612;

always @(posedge na1600)
   l448 <= na1600;

always @(posedge na1568)
   l450 <= na1568;

always @(posedge na1550)
   l452 <= na1550;

always @(posedge na1532)
   l454 <= na1532;

always @(posedge na1514)
   l456 <= na1514;

always @(posedge na1496)
   l458 <= na1496;

always @(posedge na1478)
   l460 <= na1478;

always @(posedge na1460)
   l462 <= na1460;

always @(posedge na1442)
   l464 <= na1442;

always @(posedge na1414)
   l466 <= na1414;

always @(posedge na972)
   l468 <= na972;

always @(posedge na3096)
   l470 <= na3096;

always @(posedge na3114)
   l472 <= na3114;

always @(posedge na3132)
   l474 <= na3132;

always @(posedge na3150)
   l476 <= na3150;

always @(posedge na848)
   l478 <= na848;

always @(posedge na3144)
   l480 <= na3144;

always @(posedge na3126)
   l482 <= na3126;

always @(posedge na3108)
   l484 <= na3108;

always @(posedge a3090)
   l486 <= a3090;

always @(posedge na3156)
   l488 <= na3156;

always @(posedge na3530)
   l490 <= na3530;

always @(posedge na3546)
   l492 <= na3546;

always @(posedge na3550)
   l494 <= na3550;

always @(posedge na3540)
   l496 <= na3540;

always @(posedge na3562)
   l498 <= na3562;

always @(posedge na3580)
   l500 <= na3580;

always @(posedge na3598)
   l502 <= na3598;

always @(posedge na3616)
   l504 <= na3616;

always @(posedge na3634)
   l506 <= na3634;

always @(posedge na3652)
   l508 <= na3652;

always @(posedge na3670)
   l510 <= na3670;

always @(posedge na3688)
   l512 <= na3688;

always @(posedge na3706)
   l514 <= na3706;

always @(posedge na3734)
   l516 <= na3734;

always @(posedge na3746)
   l518 <= na3746;

always @(posedge na3796)
   l520 <= na3796;

always @(posedge na3808)
   l522 <= na3808;

always @(posedge na3832)
   l524 <= na3832;

always @(posedge na3872)
   l526 <= na3872;

always @(posedge na3884)
   l528 <= na3884;

always @(posedge na3902)
   l530 <= na3902;

always @(posedge na3920)
   l532 <= na3920;

always @(posedge na3938)
   l534 <= na3938;

always @(posedge na3956)
   l536 <= na3956;

always @(posedge na3974)
   l538 <= na3974;

always @(posedge na3992)
   l540 <= na3992;

always @(posedge na4008)
   l542 <= na4008;

always @(posedge na4042)
   l544 <= na4042;

always @(posedge na4076)
   l546 <= na4076;

always @(posedge na4092)
   l548 <= na4092;

always @(posedge na4098)
   l550 <= na4098;

always @(posedge na4116)
   l552 <= na4116;

always @(posedge na4156)
   l554 <= na4156;

always @(posedge na4168)
   l556 <= na4168;

always @(posedge na4186)
   l558 <= na4186;

always @(posedge na4202)
   l560 <= na4202;

always @(posedge na4220)
   l562 <= na4220;

always @(posedge na4232)
   l564 <= na4232;

always @(posedge na4254)
   l566 <= na4254;

always @(posedge na4270)
   l568 <= na4270;

always @(posedge na4276)
   l570 <= na4276;

always @(posedge na4292)
   l572 <= na4292;

always @(posedge na4298)
   l574 <= na4298;

always @(posedge na4316)
   l576 <= na4316;

always @(posedge na4334)
   l578 <= na4334;

always @(posedge na4352)
   l580 <= na4352;

always @(posedge na3524)
   l582 <= na3524;

always @(posedge na4346)
   l584 <= na4346;

always @(posedge na4328)
   l586 <= na4328;

always @(posedge na4310)
   l588 <= na4310;

always @(posedge na4366)
   l590 <= na4366;

always @(posedge na4286)
   l592 <= na4286;

always @(posedge na4360)
   l594 <= na4360;

always @(posedge na4380)
   l596 <= na4380;

always @(posedge na4264)
   l598 <= na4264;

always @(posedge na4394)
   l600 <= na4394;

always @(posedge na4408)
   l602 <= na4408;

always @(posedge na4374)
   l604 <= na4374;

always @(posedge na4402)
   l606 <= na4402;

always @(posedge na4388)
   l608 <= na4388;

always @(posedge na4248)
   l610 <= na4248;

always @(posedge na4226)
   l612 <= na4226;

always @(posedge na4214)
   l614 <= na4214;

always @(posedge na4196)
   l616 <= na4196;

always @(posedge na4426)
   l618 <= na4426;

always @(posedge na4448)
   l620 <= na4448;

always @(posedge na4180)
   l622 <= na4180;

always @(posedge na4442)
   l624 <= na4442;

always @(posedge na4466)
   l626 <= na4466;

always @(posedge na4420)
   l628 <= na4420;

always @(posedge na4460)
   l630 <= na4460;

always @(posedge na4162)
   l632 <= na4162;

always @(posedge na4472)
   l634 <= na4472;

always @(posedge na4488)
   l636 <= na4488;

always @(posedge na4494)
   l638 <= na4494;

always @(posedge na4500)
   l640 <= na4500;

always @(posedge na4506)
   l642 <= na4506;

always @(posedge na4518)
   l644 <= na4518;

always @(posedge na4538)
   l646 <= na4538;

always @(posedge na4556)
   l648 <= na4556;

always @(posedge na4150)
   l650 <= na4150;

always @(posedge na4550)
   l652 <= na4550;

always @(posedge na4532)
   l654 <= na4532;

always @(posedge na4568)
   l656 <= na4568;

always @(posedge na4512)
   l658 <= na4512;

always @(posedge na4580)
   l660 <= na4580;

always @(posedge na4562)
   l662 <= na4562;

always @(posedge na4592)
   l664 <= na4592;

always @(posedge na4574)
   l666 <= na4574;

always @(posedge na4604)
   l668 <= na4604;

always @(posedge na4586)
   l670 <= na4586;

always @(posedge na4616)
   l672 <= na4616;

always @(posedge na4598)
   l674 <= na4598;

always @(posedge na4628)
   l676 <= na4628;

always @(posedge na4610)
   l678 <= na4610;

always @(posedge na4640)
   l680 <= na4640;

always @(posedge na4622)
   l682 <= na4622;

always @(posedge na4652)
   l684 <= na4652;

always @(posedge na4634)
   l686 <= na4634;

always @(posedge na4664)
   l688 <= na4664;

always @(posedge na4646)
   l690 <= na4646;

always @(posedge na4676)
   l692 <= na4676;

always @(posedge na4658)
   l694 <= na4658;

always @(posedge na4688)
   l696 <= na4688;

always @(posedge na4670)
   l698 <= na4670;

always @(posedge na4682)
   l700 <= na4682;

always @(posedge na4482)
   l702 <= na4482;

always @(posedge na4110)
   l704 <= na4110;

always @(posedge na4706)
   l706 <= na4706;

always @(posedge na4086)
   l708 <= na4086;

always @(posedge na4728)
   l710 <= na4728;

always @(posedge na4700)
   l712 <= na4700;

always @(posedge na4722)
   l714 <= na4722;

always @(posedge na4770)
   l716 <= na4770;

always @(posedge na4798)
   l718 <= na4798;

always @(posedge na4824)
   l720 <= na4824;

always @(posedge na4844)
   l722 <= na4844;

always @(posedge na4070)
   l724 <= na4070;

always @(posedge na4838)
   l726 <= na4838;

always @(posedge na4850)
   l728 <= na4850;

always @(posedge na4818)
   l730 <= na4818;

always @(posedge na4792)
   l732 <= na4792;

always @(posedge na4764)
   l734 <= na4764;

always @(posedge na4036)
   l736 <= na4036;

always @(posedge na4002)
   l738 <= na4002;

always @(posedge na3986)
   l740 <= na3986;

always @(posedge na3968)
   l742 <= na3968;

always @(posedge na3950)
   l744 <= na3950;

always @(posedge na3932)
   l746 <= na3932;

always @(posedge na3914)
   l748 <= na3914;

always @(posedge na4900)
   l750 <= na4900;

always @(posedge na4926)
   l752 <= na4926;

always @(posedge na4952)
   l754 <= na4952;

always @(posedge na4974)
   l756 <= na4974;

always @(posedge na4992)
   l758 <= na4992;

always @(posedge na5014)
   l760 <= na5014;

always @(posedge na5036)
   l762 <= na5036;

always @(posedge na5058)
   l764 <= na5058;

always @(posedge na5080)
   l766 <= na5080;

always @(posedge na3896)
   l768 <= na3896;

always @(posedge na5074)
   l770 <= na5074;

always @(posedge na5052)
   l772 <= na5052;

always @(posedge na5030)
   l774 <= na5030;

always @(posedge na5008)
   l776 <= na5008;

always @(posedge na4986)
   l778 <= na4986;

always @(posedge na4968)
   l780 <= na4968;

always @(posedge na4946)
   l782 <= na4946;

always @(posedge na4920)
   l784 <= na4920;

always @(posedge na4894)
   l786 <= na4894;

always @(posedge na3878)
   l788 <= na3878;

always @(posedge na3866)
   l790 <= na3866;

always @(posedge na3826)
   l792 <= na3826;

always @(posedge na3802)
   l794 <= na3802;

always @(posedge na3790)
   l796 <= na3790;

always @(posedge na3740)
   l798 <= na3740;

always @(posedge na3728)
   l800 <= na3728;

always @(posedge na3700)
   l802 <= na3700;

always @(posedge na3682)
   l804 <= na3682;

always @(posedge na3664)
   l806 <= na3664;

always @(posedge na3646)
   l808 <= na3646;

always @(posedge na3628)
   l810 <= na3628;

always @(posedge na3610)
   l812 <= na3610;

always @(posedge na3592)
   l814 <= na3592;

always @(posedge na3574)
   l816 <= na3574;

always @(posedge na3556)
   l818 <= na3556;

always @(posedge c1)
   l820 <= c1;


assign na854 = ~a854;
assign na882 = ~a882;
assign na900 = ~a900;
assign na912 = ~a912;
assign na934 = ~a934;
assign na952 = ~a952;
assign na970 = ~a970;
assign na876 = ~a876;
assign na964 = ~a964;
assign na946 = ~a946;
assign na928 = ~a928;
assign na906 = ~a906;
assign a894 = ~a892 & ~a884;
assign na978 = ~a978;
assign na1380 = ~a1380;
assign na1396 = ~a1396;
assign na1408 = ~a1408;
assign na1390 = ~a1390;
assign na1402 = ~a1402;
assign na1420 = ~a1420;
assign na1448 = ~a1448;
assign na1466 = ~a1466;
assign na1484 = ~a1484;
assign na1502 = ~a1502;
assign na1520 = ~a1520;
assign na1538 = ~a1538;
assign na1556 = ~a1556;
assign na1574 = ~a1574;
assign na1606 = ~a1606;
assign na1618 = ~a1618;
assign na1630 = ~a1630;
assign na1654 = ~a1654;
assign na1706 = ~a1706;
assign na1720 = ~a1720;
assign na1754 = ~a1754;
assign na1776 = ~a1776;
assign na1794 = ~a1794;
assign na1812 = ~a1812;
assign na1830 = ~a1830;
assign na1848 = ~a1848;
assign na1866 = ~a1866;
assign na1882 = ~a1882;
assign na1894 = ~a1894;
assign na1912 = ~a1912;
assign na1948 = ~a1948;
assign na1988 = ~a1988;
assign na2004 = ~a2004;
assign na2016 = ~a2016;
assign na2034 = ~a2034;
assign na2078 = ~a2078;
assign na2090 = ~a2090;
assign na2108 = ~a2108;
assign na2126 = ~a2126;
assign na2142 = ~a2142;
assign na2160 = ~a2160;
assign na2172 = ~a2172;
assign na2194 = ~a2194;
assign na2210 = ~a2210;
assign na2222 = ~a2222;
assign na2238 = ~a2238;
assign na2250 = ~a2250;
assign na2268 = ~a2268;
assign na2286 = ~a2286;
assign na2304 = ~a2304;
assign na1374 = ~a1374;
assign na2298 = ~a2298;
assign na2280 = ~a2280;
assign na2262 = ~a2262;
assign na2244 = ~a2244;
assign na2318 = ~a2318;
assign na2232 = ~a2232;
assign na2312 = ~a2312;
assign na2216 = ~a2216;
assign na2332 = ~a2332;
assign na2204 = ~a2204;
assign na2346 = ~a2346;
assign na2360 = ~a2360;
assign na2326 = ~a2326;
assign na2354 = ~a2354;
assign na2340 = ~a2340;
assign na2188 = ~a2188;
assign na2166 = ~a2166;
assign na2154 = ~a2154;
assign na2136 = ~a2136;
assign na2378 = ~a2378;
assign na2400 = ~a2400;
assign na2120 = ~a2120;
assign na2394 = ~a2394;
assign na2418 = ~a2418;
assign na2372 = ~a2372;
assign na2412 = ~a2412;
assign na2102 = ~a2102;
assign na2084 = ~a2084;
assign na2442 = ~a2442;
assign na2454 = ~a2454;
assign na2466 = ~a2466;
assign na2478 = ~a2478;
assign na2490 = ~a2490;
assign na2502 = ~a2502;
assign na2520 = ~a2520;
assign na2536 = ~a2536;
assign na2072 = ~a2072;
assign na2530 = ~a2530;
assign na2514 = ~a2514;
assign na2548 = ~a2548;
assign na2496 = ~a2496;
assign na2560 = ~a2560;
assign na2542 = ~a2542;
assign na2572 = ~a2572;
assign na2554 = ~a2554;
assign na2584 = ~a2584;
assign na2566 = ~a2566;
assign na2596 = ~a2596;
assign na2578 = ~a2578;
assign na2608 = ~a2608;
assign na2590 = ~a2590;
assign na2622 = ~a2622;
assign na2602 = ~a2602;
assign na2634 = ~a2634;
assign na2616 = ~a2616;
assign na2646 = ~a2646;
assign na2628 = ~a2628;
assign na2658 = ~a2658;
assign na2640 = ~a2640;
assign na2670 = ~a2670;
assign na2652 = ~a2652;
assign na2664 = ~a2664;
assign na2484 = ~a2484;
assign na2472 = ~a2472;
assign na2460 = ~a2460;
assign na2448 = ~a2448;
assign na2436 = ~a2436;
assign na2028 = ~a2028;
assign na2010 = ~a2010;
assign na2688 = ~a2688;
assign na1998 = ~a1998;
assign na2710 = ~a2710;
assign na2682 = ~a2682;
assign na2704 = ~a2704;
assign na2760 = ~a2760;
assign na2790 = ~a2790;
assign na2816 = ~a2816;
assign na2836 = ~a2836;
assign na1982 = ~a1982;
assign na2830 = ~a2830;
assign na2848 = ~a2848;
assign na2810 = ~a2810;
assign na2842 = ~a2842;
assign na2784 = ~a2784;
assign na2754 = ~a2754;
assign na1942 = ~a1942;
assign na1906 = ~a1906;
assign na1888 = ~a1888;
assign na1876 = ~a1876;
assign na1860 = ~a1860;
assign na1842 = ~a1842;
assign na1824 = ~a1824;
assign na1806 = ~a1806;
assign na1788 = ~a1788;
assign na2898 = ~a2898;
assign na2924 = ~a2924;
assign na2950 = ~a2950;
assign na2972 = ~a2972;
assign na2990 = ~a2990;
assign na3012 = ~a3012;
assign na3034 = ~a3034;
assign na3056 = ~a3056;
assign na3078 = ~a3078;
assign na1770 = ~a1770;
assign na3072 = ~a3072;
assign na3050 = ~a3050;
assign na3028 = ~a3028;
assign na3006 = ~a3006;
assign na2984 = ~a2984;
assign na2966 = ~a2966;
assign na2944 = ~a2944;
assign na2918 = ~a2918;
assign na2892 = ~a2892;
assign na1748 = ~a1748;
assign na1714 = ~a1714;
assign na1700 = ~a1700;
assign na1648 = ~a1648;
assign na1624 = ~a1624;
assign na1612 = ~a1612;
assign na1600 = ~a1600;
assign na1568 = ~a1568;
assign na1550 = ~a1550;
assign na1532 = ~a1532;
assign na1514 = ~a1514;
assign na1496 = ~a1496;
assign na1478 = ~a1478;
assign na1460 = ~a1460;
assign na1442 = ~a1442;
assign na1414 = ~a1414;
assign na972 = ~a972;
assign na3096 = ~a3096;
assign na3114 = ~a3114;
assign na3132 = ~a3132;
assign na3150 = ~a3150;
assign na848 = ~a848;
assign na3144 = ~a3144;
assign na3126 = ~a3126;
assign na3108 = ~a3108;
assign a3090 = ~a3088 & ~a3080;
assign na3156 = ~a3156;
assign na3530 = ~a3530;
assign na3546 = ~a3546;
assign na3550 = ~a3550;
assign na3540 = ~a3540;
assign na3562 = ~a3562;
assign na3580 = ~a3580;
assign na3598 = ~a3598;
assign na3616 = ~a3616;
assign na3634 = ~a3634;
assign na3652 = ~a3652;
assign na3670 = ~a3670;
assign na3688 = ~a3688;
assign na3706 = ~a3706;
assign na3734 = ~a3734;
assign na3746 = ~a3746;
assign na3796 = ~a3796;
assign na3808 = ~a3808;
assign na3832 = ~a3832;
assign na3872 = ~a3872;
assign na3884 = ~a3884;
assign na3902 = ~a3902;
assign na3920 = ~a3920;
assign na3938 = ~a3938;
assign na3956 = ~a3956;
assign na3974 = ~a3974;
assign na3992 = ~a3992;
assign na4008 = ~a4008;
assign na4042 = ~a4042;
assign na4076 = ~a4076;
assign na4092 = ~a4092;
assign na4098 = ~a4098;
assign na4116 = ~a4116;
assign na4156 = ~a4156;
assign na4168 = ~a4168;
assign na4186 = ~a4186;
assign na4202 = ~a4202;
assign na4220 = ~a4220;
assign na4232 = ~a4232;
assign na4254 = ~a4254;
assign na4270 = ~a4270;
assign na4276 = ~a4276;
assign na4292 = ~a4292;
assign na4298 = ~a4298;
assign na4316 = ~a4316;
assign na4334 = ~a4334;
assign na4352 = ~a4352;
assign na3524 = ~a3524;
assign na4346 = ~a4346;
assign na4328 = ~a4328;
assign na4310 = ~a4310;
assign na4366 = ~a4366;
assign na4286 = ~a4286;
assign na4360 = ~a4360;
assign na4380 = ~a4380;
assign na4264 = ~a4264;
assign na4394 = ~a4394;
assign na4408 = ~a4408;
assign na4374 = ~a4374;
assign na4402 = ~a4402;
assign na4388 = ~a4388;
assign na4248 = ~a4248;
assign na4226 = ~a4226;
assign na4214 = ~a4214;
assign na4196 = ~a4196;
assign na4426 = ~a4426;
assign na4448 = ~a4448;
assign na4180 = ~a4180;
assign na4442 = ~a4442;
assign na4466 = ~a4466;
assign na4420 = ~a4420;
assign na4460 = ~a4460;
assign na4162 = ~a4162;
assign na4472 = ~a4472;
assign na4488 = ~a4488;
assign na4494 = ~a4494;
assign na4500 = ~a4500;
assign na4506 = ~a4506;
assign na4518 = ~a4518;
assign na4538 = ~a4538;
assign na4556 = ~a4556;
assign na4150 = ~a4150;
assign na4550 = ~a4550;
assign na4532 = ~a4532;
assign na4568 = ~a4568;
assign na4512 = ~a4512;
assign na4580 = ~a4580;
assign na4562 = ~a4562;
assign na4592 = ~a4592;
assign na4574 = ~a4574;
assign na4604 = ~a4604;
assign na4586 = ~a4586;
assign na4616 = ~a4616;
assign na4598 = ~a4598;
assign na4628 = ~a4628;
assign na4610 = ~a4610;
assign na4640 = ~a4640;
assign na4622 = ~a4622;
assign na4652 = ~a4652;
assign na4634 = ~a4634;
assign na4664 = ~a4664;
assign na4646 = ~a4646;
assign na4676 = ~a4676;
assign na4658 = ~a4658;
assign na4688 = ~a4688;
assign na4670 = ~a4670;
assign na4682 = ~a4682;
assign na4482 = ~a4482;
assign na4110 = ~a4110;
assign na4706 = ~a4706;
assign na4086 = ~a4086;
assign na4728 = ~a4728;
assign na4700 = ~a4700;
assign na4722 = ~a4722;
assign na4770 = ~a4770;
assign na4798 = ~a4798;
assign na4824 = ~a4824;
assign na4844 = ~a4844;
assign na4070 = ~a4070;
assign na4838 = ~a4838;
assign na4850 = ~a4850;
assign na4818 = ~a4818;
assign na4792 = ~a4792;
assign na4764 = ~a4764;
assign na4036 = ~a4036;
assign na4002 = ~a4002;
assign na3986 = ~a3986;
assign na3968 = ~a3968;
assign na3950 = ~a3950;
assign na3932 = ~a3932;
assign na3914 = ~a3914;
assign na4900 = ~a4900;
assign na4926 = ~a4926;
assign na4952 = ~a4952;
assign na4974 = ~a4974;
assign na4992 = ~a4992;
assign na5014 = ~a5014;
assign na5036 = ~a5036;
assign na5058 = ~a5058;
assign na5080 = ~a5080;
assign na3896 = ~a3896;
assign na5074 = ~a5074;
assign na5052 = ~a5052;
assign na5030 = ~a5030;
assign na5008 = ~a5008;
assign na4986 = ~a4986;
assign na4968 = ~a4968;
assign na4946 = ~a4946;
assign na4920 = ~a4920;
assign na4894 = ~a4894;
assign na3878 = ~a3878;
assign na3866 = ~a3866;
assign na3826 = ~a3826;
assign na3802 = ~a3802;
assign na3790 = ~a3790;
assign na3740 = ~a3740;
assign na3728 = ~a3728;
assign na3700 = ~a3700;
assign na3682 = ~a3682;
assign na3664 = ~a3664;
assign na3646 = ~a3646;
assign na3628 = ~a3628;
assign na3610 = ~a3610;
assign na3592 = ~a3592;
assign na3574 = ~a3574;
assign na3556 = ~a3556;
assign c1 = 1;
assign a822 = l80 & ~l78;
assign a824 = ~l80 & l78;
assign a826 = ~a824 & ~a822;
assign a828 = l470 & ~l84;
assign a830 = a828 & l86;
assign a832 = ~a830 & i2;
assign a834 = l476 & ~l474;
assign a836 = a834 & ~l472;
assign a838 = a836 & l84;
assign a840 = ~l84 & l78;
assign a842 = ~a840 & ~a838;
assign a844 = ~a842 & l86;
assign a846 = l478 & ~l86;
assign a848 = ~a846 & ~a844;
assign a850 = ~a848 & a832;
assign a852 = ~a832 & l78;
assign a854 = ~a852 & ~a850;
assign a856 = ~l84 & l82;
assign a858 = a856 & l86;
assign a860 = ~a858 & i2;
assign a862 = l90 & ~l88;
assign a864 = a862 & ~l92;
assign a866 = a864 & l84;
assign a868 = ~l84 & l80;
assign a870 = ~a868 & ~a866;
assign a872 = ~a870 & l86;
assign a874 = l94 & ~l86;
assign a876 = ~a874 & ~a872;
assign a878 = ~a876 & a860;
assign a880 = ~a860 & l80;
assign a882 = ~a880 & ~a878;
assign a884 = ~l104 & ~l86;
assign a886 = ~a856 & l106;
assign a888 = l110 & l108;
assign a890 = ~a888 & l86;
assign a892 = a890 & a886;
assign a896 = a894 & a860;
assign a898 = ~a860 & l82;
assign a900 = ~a898 & ~a896;
assign a902 = l86 & i12;
assign a904 = l102 & ~l86;
assign a906 = ~a904 & ~a902;
assign a908 = ~a906 & i2;
assign a910 = l84 & ~i2;
assign a912 = ~a910 & ~a908;
assign a914 = l86 & i4;
assign a916 = ~a914 & i2;
assign a918 = a856 & i10;
assign a920 = ~a856 & l88;
assign a922 = ~a920 & ~a918;
assign a924 = ~a922 & l86;
assign a926 = l100 & ~l86;
assign a928 = ~a926 & ~a924;
assign a930 = ~a928 & a916;
assign a932 = ~a916 & l88;
assign a934 = ~a932 & ~a930;
assign a936 = a856 & i8;
assign a938 = ~a856 & l90;
assign a940 = ~a938 & ~a936;
assign a942 = ~a940 & l86;
assign a944 = l98 & ~l86;
assign a946 = ~a944 & ~a942;
assign a948 = ~a946 & a916;
assign a950 = ~a916 & l90;
assign a952 = ~a950 & ~a948;
assign a954 = a856 & i6;
assign a956 = ~a856 & l92;
assign a958 = ~a956 & ~a954;
assign a960 = ~a958 & l86;
assign a962 = l96 & ~l86;
assign a964 = ~a962 & ~a960;
assign a966 = ~a964 & a916;
assign a968 = ~a916 & l92;
assign a970 = ~a968 & ~a966;
assign a972 = ~l468 & ~l86;
assign a974 = ~a972 & a860;
assign a976 = ~a860 & l106;
assign a978 = ~a976 & ~a974;
assign a980 = ~l128 & ~l126;
assign a982 = a980 & ~l124;
assign a984 = a982 & ~l122;
assign a986 = a984 & l120;
assign a988 = l130 & ~l120;
assign a990 = a988 & a984;
assign a992 = ~l130 & ~l120;
assign a994 = a992 & a982;
assign a996 = ~a994 & ~a990;
assign a998 = a996 & ~a986;
assign a1000 = ~l90 & l88;
assign a1002 = l132 & l92;
assign a1004 = ~a1002 & a1000;
assign a1006 = a1004 & ~a998;
assign a1008 = l90 & l88;
assign a1010 = l130 & l120;
assign a1012 = a1010 & l122;
assign a1014 = l128 & l124;
assign a1016 = a1014 & l126;
assign a1018 = a1016 & a1012;
assign a1020 = a1018 & ~a1008;
assign a1022 = a864 & l134;
assign a1024 = a1022 & ~l132;
assign a1026 = a1024 & a986;
assign a1028 = ~a1026 & ~a1020;
assign a1030 = a1028 & ~a1006;
assign a1032 = ~l150 & ~l148;
assign a1034 = a1032 & ~l146;
assign a1036 = ~a1034 & ~l144;
assign a1038 = ~l158 & l156;
assign a1040 = a1038 & ~l154;
assign a1042 = a1040 & ~l152;
assign a1044 = ~l158 & ~l156;
assign a1046 = l160 & l152;
assign a1048 = a1046 & ~l154;
assign a1050 = a1048 & a1044;
assign a1052 = ~a1050 & ~a1042;
assign a1054 = ~l128 & l126;
assign a1056 = a1054 & ~l124;
assign a1058 = a1056 & a992;
assign a1060 = a1058 & ~l122;
assign a1062 = a1060 & ~a1052;
assign a1064 = ~l160 & l152;
assign a1066 = a1044 & l154;
assign a1068 = ~a1066 & ~a1040;
assign a1070 = ~a1068 & a1064;
assign a1072 = a1070 & ~a998;
assign a1074 = ~a1072 & ~a1062;
assign a1076 = a1074 & a1036;
assign a1078 = ~a1060 & a998;
assign a1080 = ~a1078 & a1000;
assign a1082 = a1080 & a1076;
assign a1084 = a1082 & l142;
assign a1086 = ~a1024 & ~l88;
assign a1088 = ~a1086 & a1060;
assign a1090 = ~a1088 & a998;
assign a1092 = a1090 & l112;
assign a1094 = l140 & ~l108;
assign a1096 = l162 & i14;
assign a1098 = ~a1096 & ~a1094;
assign a1100 = a1098 & ~a1092;
assign a1102 = a1100 & ~a1084;
assign a1104 = a1102 & ~l140;
assign a1106 = ~a1018 & l112;
assign a1108 = l164 & ~l108;
assign a1110 = l166 & i16;
assign a1112 = ~a1110 & ~a1108;
assign a1114 = a1112 & ~a1106;
assign a1116 = a1114 & ~l164;
assign a1118 = ~a1116 & l150;
assign a1120 = a1118 & ~a1104;
assign a1122 = a1120 & l138;
assign a1124 = a1122 & l168;
assign a1126 = a1124 & l136;
assign a1128 = a1124 & l170;
assign a1130 = ~a1128 & ~a1126;
assign a1132 = ~a1130 & ~a1030;
assign a1134 = l118 & ~l108;
assign a1136 = a1134 & ~a1132;
assign a1138 = l174 & l172;
assign a1140 = ~l90 & ~l88;
assign a1142 = ~l134 & l92;
assign a1144 = a1142 & a1140;
assign a1146 = a1144 & l130;
assign a1148 = a1056 & l122;
assign a1150 = a1148 & l120;
assign a1152 = a1150 & ~a1146;
assign a1154 = a1014 & ~l126;
assign a1156 = a1154 & a1012;
assign a1158 = ~a1156 & ~a1058;
assign a1160 = a1158 & ~a1152;
assign a1162 = a1002 & a1000;
assign a1164 = ~a1162 & ~a1008;
assign a1166 = ~a1164 & a986;
assign a1168 = a1018 & a1008;
assign a1170 = a1010 & ~l122;
assign a1172 = a980 & l124;
assign a1174 = a1172 & a1170;
assign a1176 = ~a1174 & ~a1168;
assign a1178 = a1176 & ~a1166;
assign a1180 = a1178 & a1160;
assign a1182 = a1164 & ~a1022;
assign a1184 = ~a1182 & ~a996;
assign a1186 = a1148 & a1010;
assign a1188 = a1172 & l122;
assign a1190 = a1188 & ~a1010;
assign a1192 = ~a1190 & ~a1186;
assign a1194 = ~a1192 & a1144;
assign a1196 = a1154 & ~l120;
assign a1198 = ~l176 & ~l130;
assign a1200 = a1198 & l122;
assign a1202 = ~a1200 & a1196;
assign a1204 = ~a1202 & ~a1188;
assign a1206 = a1204 & ~a1194;
assign a1208 = a1206 & ~a1184;
assign a1210 = a1208 & a1180;
assign a1212 = a1210 & l112;
assign a1214 = ~a1212 & ~a1138;
assign a1216 = a1214 & ~a1136;
assign a1218 = a1216 & ~l118;
assign a1220 = l178 & l86;
assign a1222 = a1220 & a1120;
assign a1224 = a1222 & ~a1218;
assign a1226 = a1008 & ~l92;
assign a1228 = a1226 & ~l134;
assign a1230 = a990 & ~l182;
assign a1232 = a1230 & a1228;
assign a1234 = a1188 & ~a1144;
assign a1236 = ~a1234 & ~a1232;
assign a1238 = a1236 & a1160;
assign a1240 = l132 & l88;
assign a1242 = a1240 & ~a1238;
assign a1244 = ~a1018 & a998;
assign a1246 = a1000 & ~l92;
assign a1248 = a1246 & l134;
assign a1250 = a1248 & ~a1244;
assign a1252 = a1000 & l92;
assign a1254 = ~a1252 & ~a1226;
assign a1256 = ~a1254 & l134;
assign a1258 = a1256 & ~a998;
assign a1260 = a1258 & l132;
assign a1262 = ~a1260 & ~a1250;
assign a1264 = a1262 & ~a1242;
assign a1266 = ~a1264 & l136;
assign a1268 = ~a1248 & ~a1194;
assign a1270 = ~a1268 & ~l136;
assign a1272 = ~a1270 & ~a1266;
assign a1274 = a1272 & l160;
assign a1276 = ~a1274 & ~l152;
assign a1278 = a1038 & l154;
assign a1280 = a1278 & ~a1046;
assign a1282 = a1280 & ~a1276;
assign a1284 = a1036 & l184;
assign a1286 = a1284 & ~a1282;
assign a1288 = a1286 & ~a1272;
assign a1290 = ~a1126 & ~l108;
assign a1292 = a1290 & l180;
assign a1294 = l186 & i18;
assign a1296 = a1008 & l188;
assign a1298 = ~a1296 & ~a1000;
assign a1300 = ~a1298 & a1142;
assign a1302 = ~a1300 & ~a1228;
assign a1304 = a1302 & ~a1246;
assign a1306 = ~a1304 & ~a1204;
assign a1308 = ~a1306 & ~a1194;
assign a1310 = a1308 & l112;
assign a1312 = ~a1310 & ~a1294;
assign a1314 = a1312 & ~a1292;
assign a1316 = a1314 & ~a1288;
assign a1318 = a1316 & ~l180;
assign a1320 = a1084 & l192;
assign a1322 = l190 & ~l108;
assign a1324 = l196 & l194;
assign a1326 = ~a1324 & ~a1322;
assign a1328 = a1306 & ~a1248;
assign a1330 = ~a1328 & a1092;
assign a1332 = ~a1330 & a1326;
assign a1334 = a1332 & ~a1320;
assign a1336 = a1334 & ~l190;
assign a1338 = ~a1272 & a1242;
assign a1340 = ~a1338 & a1126;
assign a1342 = ~a1340 & ~a1128;
assign a1344 = l138 & ~l108;
assign a1346 = a1344 & a1342;
assign a1348 = l200 & l198;
assign a1350 = ~l206 & ~l204;
assign a1352 = a1350 & l202;
assign a1354 = ~a1352 & ~a1348;
assign a1356 = a1238 & ~a1202;
assign a1358 = a1356 & l112;
assign a1360 = ~a1358 & a1354;
assign a1362 = a1360 & ~a1346;
assign a1364 = a1362 & ~l138;
assign a1366 = ~a1364 & ~a1336;
assign a1368 = a1366 & ~a1318;
assign a1370 = a1368 & a1224;
assign a1372 = l208 & ~l86;
assign a1374 = ~a1372 & ~a1370;
assign a1376 = ~a1374 & a860;
assign a1378 = ~a860 & l108;
assign a1380 = ~a1378 & ~a1376;
assign a1382 = l110 & ~l108;
assign a1384 = ~a1382 & ~l112;
assign a1386 = ~a1384 & l86;
assign a1388 = l114 & ~l86;
assign a1390 = ~a1388 & ~a1386;
assign a1392 = ~a1390 & a860;
assign a1394 = ~a860 & l110;
assign a1396 = ~a1394 & ~a1392;
assign a1398 = l86 & l84;
assign a1400 = l116 & ~l86;
assign a1402 = ~a1400 & ~a1398;
assign a1404 = ~a1402 & a860;
assign a1406 = ~a860 & l112;
assign a1408 = ~a1406 & ~a1404;
assign a1410 = ~a1216 & l86;
assign a1412 = l466 & ~l86;
assign a1414 = ~a1412 & ~a1410;
assign a1416 = ~a1414 & a860;
assign a1418 = ~a860 & l118;
assign a1420 = ~a1418 & ~a1416;
assign a1422 = i74 & i70;
assign a1424 = i72 & i66;
assign a1426 = a1424 & i68;
assign a1428 = a1426 & a1422;
assign a1430 = ~a1428 & i76;
assign a1432 = a1430 & a856;
assign a1434 = ~a856 & l120;
assign a1436 = ~a1434 & ~a1432;
assign a1438 = ~a1436 & l86;
assign a1440 = l464 & ~l86;
assign a1442 = ~a1440 & ~a1438;
assign a1444 = ~a1442 & a916;
assign a1446 = ~a916 & l120;
assign a1448 = ~a1446 & ~a1444;
assign a1450 = a856 & i74;
assign a1452 = ~a856 & l122;
assign a1454 = ~a1452 & ~a1450;
assign a1456 = ~a1454 & l86;
assign a1458 = l462 & ~l86;
assign a1460 = ~a1458 & ~a1456;
assign a1462 = ~a1460 & a916;
assign a1464 = ~a916 & l122;
assign a1466 = ~a1464 & ~a1462;
assign a1468 = a856 & i72;
assign a1470 = ~a856 & l124;
assign a1472 = ~a1470 & ~a1468;
assign a1474 = ~a1472 & l86;
assign a1476 = l460 & ~l86;
assign a1478 = ~a1476 & ~a1474;
assign a1480 = ~a1478 & a916;
assign a1482 = ~a916 & l124;
assign a1484 = ~a1482 & ~a1480;
assign a1486 = a856 & i70;
assign a1488 = ~a856 & l126;
assign a1490 = ~a1488 & ~a1486;
assign a1492 = ~a1490 & l86;
assign a1494 = l458 & ~l86;
assign a1496 = ~a1494 & ~a1492;
assign a1498 = ~a1496 & a916;
assign a1500 = ~a916 & l126;
assign a1502 = ~a1500 & ~a1498;
assign a1504 = a856 & i68;
assign a1506 = ~a856 & l128;
assign a1508 = ~a1506 & ~a1504;
assign a1510 = ~a1508 & l86;
assign a1512 = l456 & ~l86;
assign a1514 = ~a1512 & ~a1510;
assign a1516 = ~a1514 & a916;
assign a1518 = ~a916 & l128;
assign a1520 = ~a1518 & ~a1516;
assign a1522 = a856 & i66;
assign a1524 = ~a856 & l130;
assign a1526 = ~a1524 & ~a1522;
assign a1528 = ~a1526 & l86;
assign a1530 = l454 & ~l86;
assign a1532 = ~a1530 & ~a1528;
assign a1534 = ~a1532 & a916;
assign a1536 = ~a916 & l130;
assign a1538 = ~a1536 & ~a1534;
assign a1540 = a856 & i64;
assign a1542 = ~a856 & l132;
assign a1544 = ~a1542 & ~a1540;
assign a1546 = ~a1544 & l86;
assign a1548 = l452 & ~l86;
assign a1550 = ~a1548 & ~a1546;
assign a1552 = ~a1550 & a916;
assign a1554 = ~a916 & l132;
assign a1556 = ~a1554 & ~a1552;
assign a1558 = a856 & i62;
assign a1560 = ~a856 & l134;
assign a1562 = ~a1560 & ~a1558;
assign a1564 = ~a1562 & l86;
assign a1566 = l450 & ~l86;
assign a1568 = ~a1566 & ~a1564;
assign a1570 = ~a1568 & a916;
assign a1572 = ~a916 & l134;
assign a1574 = ~a1572 & ~a1570;
assign a1576 = l362 & l358;
assign a1578 = ~l360 & ~l358;
assign a1580 = ~a1578 & ~l364;
assign a1582 = a1580 & ~a1576;
assign a1584 = a1582 & ~a1090;
assign a1586 = ~a1304 & a1018;
assign a1588 = ~a1586 & l276;
assign a1590 = a1588 & ~a1584;
assign a1592 = ~l276 & ~l136;
assign a1594 = ~a1592 & a890;
assign a1596 = a1594 & ~a1590;
assign a1598 = l448 & ~l86;
assign a1600 = ~a1598 & ~a1596;
assign a1602 = ~a1600 & a860;
assign a1604 = ~a860 & l136;
assign a1606 = ~a1604 & ~a1602;
assign a1608 = ~a1362 & l86;
assign a1610 = l446 & ~l86;
assign a1612 = ~a1610 & ~a1608;
assign a1614 = ~a1612 & a860;
assign a1616 = ~a860 & l138;
assign a1618 = ~a1616 & ~a1614;
assign a1620 = ~a1102 & l86;
assign a1622 = l444 & ~l86;
assign a1624 = ~a1622 & ~a1620;
assign a1626 = ~a1624 & a860;
assign a1628 = ~a860 & l140;
assign a1630 = ~a1628 & ~a1626;
assign a1632 = ~a1090 & l112;
assign a1634 = ~a1074 & a1036;
assign a1636 = ~a1634 & a1080;
assign a1638 = a1636 & l142;
assign a1640 = a1638 & ~a1082;
assign a1642 = ~a1640 & ~a1632;
assign a1644 = ~a1642 & l86;
assign a1646 = l442 & ~l86;
assign a1648 = ~a1646 & ~a1644;
assign a1650 = ~a1648 & a860;
assign a1652 = ~a860 & l142;
assign a1654 = ~a1652 & ~a1650;
assign a1656 = a1282 & a1036;
assign a1658 = a1656 & l184;
assign a1660 = a1658 & l146;
assign a1662 = ~l230 & ~l186;
assign a1664 = ~l256 & ~l248;
assign a1666 = a1664 & a1662;
assign a1668 = ~a1666 & ~l184;
assign a1670 = ~a1668 & l144;
assign a1672 = a1670 & i50;
assign a1674 = ~a1672 & l144;
assign a1676 = l122 & l90;
assign a1678 = ~a1676 & a1058;
assign a1680 = ~a1678 & ~a1152;
assign a1682 = ~a1680 & l88;
assign a1684 = ~a1682 & a998;
assign a1686 = a1684 & a1308;
assign a1688 = ~a1686 & l112;
assign a1690 = ~a1688 & ~a1674;
assign a1692 = a1690 & ~a1126;
assign a1694 = a1692 & ~a1660;
assign a1696 = ~a1694 & l86;
assign a1698 = l440 & ~l86;
assign a1700 = ~a1698 & ~a1696;
assign a1702 = ~a1700 & a860;
assign a1704 = ~a860 & l144;
assign a1706 = ~a1704 & ~a1702;
assign a1708 = l86 & i50;
assign a1710 = a1708 & a1670;
assign a1712 = l438 & ~l86;
assign a1714 = ~a1712 & ~a1710;
assign a1716 = ~a1714 & a860;
assign a1718 = ~a860 & l146;
assign a1720 = ~a1718 & ~a1716;
assign a1722 = ~a1658 & l146;
assign a1724 = ~l400 & ~l398;
assign a1726 = ~l404 & ~l402;
assign a1728 = a1726 & a1724;
assign a1730 = ~l408 & ~l406;
assign a1732 = ~l412 & ~l410;
assign a1734 = a1732 & ~l414;
assign a1736 = a1734 & a1730;
assign a1738 = a1736 & a1728;
assign a1740 = ~a1738 & l148;
assign a1742 = ~a1740 & ~a1722;
assign a1744 = ~a1742 & l86;
assign a1746 = l436 & ~l86;
assign a1748 = ~a1746 & ~a1744;
assign a1750 = ~a1748 & a860;
assign a1752 = ~a860 & l148;
assign a1754 = ~a1752 & ~a1750;
assign a1756 = a1290 & l150;
assign a1758 = a1738 & l148;
assign a1760 = a1686 & l112;
assign a1762 = ~a1760 & ~a1758;
assign a1764 = a1762 & ~a1756;
assign a1766 = ~a1764 & l86;
assign a1768 = l416 & ~l86;
assign a1770 = ~a1768 & ~a1766;
assign a1772 = ~a1770 & a860;
assign a1774 = ~a860 & l150;
assign a1776 = ~a1774 & ~a1772;
assign a1778 = a1672 & i60;
assign a1780 = ~a1672 & l152;
assign a1782 = ~a1780 & ~a1778;
assign a1784 = ~a1782 & l86;
assign a1786 = l396 & ~l86;
assign a1788 = ~a1786 & ~a1784;
assign a1790 = ~a1788 & a860;
assign a1792 = ~a860 & l152;
assign a1794 = ~a1792 & ~a1790;
assign a1796 = a1672 & i58;
assign a1798 = ~a1672 & l154;
assign a1800 = ~a1798 & ~a1796;
assign a1802 = ~a1800 & l86;
assign a1804 = l394 & ~l86;
assign a1806 = ~a1804 & ~a1802;
assign a1808 = ~a1806 & a860;
assign a1810 = ~a860 & l154;
assign a1812 = ~a1810 & ~a1808;
assign a1814 = a1672 & i56;
assign a1816 = ~a1672 & l156;
assign a1818 = ~a1816 & ~a1814;
assign a1820 = ~a1818 & l86;
assign a1822 = l392 & ~l86;
assign a1824 = ~a1822 & ~a1820;
assign a1826 = ~a1824 & a860;
assign a1828 = ~a860 & l156;
assign a1830 = ~a1828 & ~a1826;
assign a1832 = a1672 & i54;
assign a1834 = ~a1672 & l158;
assign a1836 = ~a1834 & ~a1832;
assign a1838 = ~a1836 & l86;
assign a1840 = l390 & ~l86;
assign a1842 = ~a1840 & ~a1838;
assign a1844 = ~a1842 & a860;
assign a1846 = ~a860 & l158;
assign a1848 = ~a1846 & ~a1844;
assign a1850 = a1672 & i52;
assign a1852 = ~a1672 & l160;
assign a1854 = ~a1852 & ~a1850;
assign a1856 = ~a1854 & l86;
assign a1858 = l388 & ~l86;
assign a1860 = ~a1858 & ~a1856;
assign a1862 = ~a1860 & a860;
assign a1864 = ~a860 & l160;
assign a1866 = ~a1864 & ~a1862;
assign a1868 = l162 & ~i14;
assign a1870 = ~a1868 & ~l232;
assign a1872 = ~a1870 & l86;
assign a1874 = l386 & ~l86;
assign a1876 = ~a1874 & ~a1872;
assign a1878 = ~a1876 & a860;
assign a1880 = ~a860 & l162;
assign a1882 = ~a1880 & ~a1878;
assign a1884 = ~a1114 & l86;
assign a1886 = l384 & ~l86;
assign a1888 = ~a1886 & ~a1884;
assign a1890 = ~a1888 & a860;
assign a1892 = ~a860 & l164;
assign a1894 = ~a1892 & ~a1890;
assign a1896 = a1018 & l112;
assign a1898 = l166 & ~i16;
assign a1900 = ~a1898 & ~a1896;
assign a1902 = ~a1900 & l86;
assign a1904 = l382 & ~l86;
assign a1906 = ~a1904 & ~a1902;
assign a1908 = ~a1906 & a860;
assign a1910 = ~a860 & l166;
assign a1912 = ~a1910 & ~a1908;
assign a1914 = ~a1308 & l270;
assign a1916 = ~l274 & ~l270;
assign a1918 = a1916 & ~l272;
assign a1920 = a1244 & ~a1088;
assign a1922 = ~a1920 & ~a1918;
assign a1924 = ~a1922 & ~a1914;
assign a1926 = l278 & l276;
assign a1928 = a1926 & ~a1924;
assign a1930 = ~l170 & ~l136;
assign a1932 = ~a1930 & l168;
assign a1934 = a1932 & ~a1122;
assign a1936 = ~a1934 & ~a1928;
assign a1938 = ~a1936 & l86;
assign a1940 = l380 & ~l86;
assign a1942 = ~a1940 & ~a1938;
assign a1944 = ~a1942 & a860;
assign a1946 = ~a860 & l168;
assign a1948 = ~a1946 & ~a1944;
assign a1950 = l364 & ~l362;
assign a1952 = a1950 & a1578;
assign a1954 = ~l364 & l360;
assign a1956 = a1954 & a1576;
assign a1958 = ~a1956 & ~a1952;
assign a1960 = ~a1958 & ~a1090;
assign a1962 = ~a1256 & ~a862;
assign a1964 = ~a1962 & a1018;
assign a1966 = a1022 & a986;
assign a1968 = ~a1966 & l276;
assign a1970 = a1968 & ~a1964;
assign a1972 = a1970 & ~a1960;
assign a1974 = ~l276 & ~l170;
assign a1976 = ~a1974 & a890;
assign a1978 = a1976 & ~a1972;
assign a1980 = l366 & ~l86;
assign a1982 = ~a1980 & ~a1978;
assign a1984 = ~a1982 & a860;
assign a1986 = ~a860 & l170;
assign a1988 = ~a1986 & ~a1984;
assign a1990 = ~l174 & l172;
assign a1992 = ~a1990 & ~l348;
assign a1994 = ~a1992 & l86;
assign a1996 = l350 & ~l86;
assign a1998 = ~a1996 & ~a1994;
assign a2000 = ~a1998 & a860;
assign a2002 = ~a860 & l172;
assign a2004 = ~a2002 & ~a2000;
assign a2006 = l86 & i46;
assign a2008 = l346 & ~l86;
assign a2010 = ~a2008 & ~a2006;
assign a2012 = ~a2010 & a860;
assign a2014 = ~a860 & l174;
assign a2016 = ~a2014 & ~a2012;
assign a2018 = a856 & i44;
assign a2020 = ~a856 & l176;
assign a2022 = ~a2020 & ~a2018;
assign a2024 = ~a2022 & l86;
assign a2026 = l344 & ~l86;
assign a2028 = ~a2026 & ~a2024;
assign a2030 = ~a2028 & a916;
assign a2032 = ~a916 & l176;
assign a2034 = ~a2032 & ~a2030;
assign a2036 = a1084 & l266;
assign a2038 = ~a1328 & a1090;
assign a2040 = a2038 & ~a1018;
assign a2042 = ~a2040 & l268;
assign a2044 = ~a2042 & l112;
assign a2046 = ~a2044 & ~a2036;
assign a2048 = a1926 & a1924;
assign a2050 = ~l186 & ~l180;
assign a2052 = ~a2050 & l138;
assign a2054 = a2052 & l280;
assign a2056 = l178 & ~l108;
assign a2058 = a1930 & l168;
assign a2060 = ~a2058 & ~a2056;
assign a2062 = a2060 & ~a2054;
assign a2064 = a2062 & ~a2048;
assign a2066 = a2064 & a2046;
assign a2068 = ~a2066 & l86;
assign a2070 = l282 & ~l86;
assign a2072 = ~a2070 & ~a2068;
assign a2074 = ~a2072 & a860;
assign a2076 = ~a860 & l178;
assign a2078 = ~a2076 & ~a2074;
assign a2080 = ~a1316 & l86;
assign a2082 = l264 & ~l86;
assign a2084 = ~a2082 & ~a2080;
assign a2086 = ~a2084 & a860;
assign a2088 = ~a860 & l180;
assign a2090 = ~a2088 & ~a2086;
assign a2092 = l84 & i34;
assign a2094 = l182 & ~l84;
assign a2096 = ~a2094 & ~a2092;
assign a2098 = ~a2096 & l86;
assign a2100 = l262 & ~l86;
assign a2102 = ~a2100 & ~a2098;
assign a2104 = ~a2102 & a860;
assign a2106 = ~a860 & l182;
assign a2108 = ~a2106 & ~a2104;
assign a2110 = ~l250 & l248;
assign a2112 = ~a1036 & l184;
assign a2114 = ~a2112 & ~a2110;
assign a2116 = ~a2114 & l86;
assign a2118 = l252 & ~l86;
assign a2120 = ~a2118 & ~a2116;
assign a2122 = ~a2120 & a860;
assign a2124 = ~a860 & l184;
assign a2126 = ~a2124 & ~a2122;
assign a2128 = l186 & ~i18;
assign a2130 = ~a2128 & ~l230;
assign a2132 = ~a2130 & l86;
assign a2134 = l246 & ~l86;
assign a2136 = ~a2134 & ~a2132;
assign a2138 = ~a2136 & a860;
assign a2140 = ~a860 & l186;
assign a2142 = ~a2140 & ~a2138;
assign a2144 = a856 & i28;
assign a2146 = ~a856 & l188;
assign a2148 = ~a2146 & ~a2144;
assign a2150 = ~a2148 & l86;
assign a2152 = l244 & ~l86;
assign a2154 = ~a2152 & ~a2150;
assign a2156 = ~a2154 & a916;
assign a2158 = ~a916 & l188;
assign a2160 = ~a2158 & ~a2156;
assign a2162 = ~a1334 & l86;
assign a2164 = l242 & ~l86;
assign a2166 = ~a2164 & ~a2162;
assign a2168 = ~a2166 & a860;
assign a2170 = ~a860 & l190;
assign a2172 = ~a2170 & ~a2168;
assign a2174 = ~a2038 & l84;
assign a2176 = ~l232 & ~l230;
assign a2178 = a2176 & l192;
assign a2180 = a2178 & ~a1084;
assign a2182 = ~a2180 & ~a2174;
assign a2184 = ~a2182 & l86;
assign a2186 = l240 & ~l86;
assign a2188 = ~a2186 & ~a2184;
assign a2190 = ~a2188 & a860;
assign a2192 = ~a860 & l192;
assign a2194 = ~a2192 & ~a2190;
assign a2196 = ~l196 & l194;
assign a2198 = ~a2196 & ~l226;
assign a2200 = ~a2198 & l86;
assign a2202 = l228 & ~l86;
assign a2204 = ~a2202 & ~a2200;
assign a2206 = ~a2204 & a860;
assign a2208 = ~a860 & l194;
assign a2210 = ~a2208 & ~a2206;
assign a2212 = l86 & i26;
assign a2214 = l224 & ~l86;
assign a2216 = ~a2214 & ~a2212;
assign a2218 = ~a2216 & a860;
assign a2220 = ~a860 & l196;
assign a2222 = ~a2220 & ~a2218;
assign a2224 = ~l200 & l198;
assign a2226 = ~a2224 & ~l218;
assign a2228 = ~a2226 & l86;
assign a2230 = l220 & ~l86;
assign a2232 = ~a2230 & ~a2228;
assign a2234 = ~a2232 & a860;
assign a2236 = ~a860 & l198;
assign a2238 = ~a2236 & ~a2234;
assign a2240 = l86 & i24;
assign a2242 = l216 & ~l86;
assign a2244 = ~a2242 & ~a2240;
assign a2246 = ~a2244 & a860;
assign a2248 = ~a860 & l200;
assign a2250 = ~a2248 & ~a2246;
assign a2252 = ~a1356 & l112;
assign a2254 = ~a1342 & l138;
assign a2256 = ~a2254 & ~a2252;
assign a2258 = ~a2256 & l86;
assign a2260 = l214 & ~l86;
assign a2262 = ~a2260 & ~a2258;
assign a2264 = ~a2262 & a860;
assign a2266 = ~a860 & l202;
assign a2268 = ~a2266 & ~a2264;
assign a2270 = a856 & i22;
assign a2272 = ~a856 & l204;
assign a2274 = ~a2272 & ~a2270;
assign a2276 = ~a2274 & l86;
assign a2278 = l212 & ~l86;
assign a2280 = ~a2278 & ~a2276;
assign a2282 = ~a2280 & a916;
assign a2284 = ~a916 & l204;
assign a2286 = ~a2284 & ~a2282;
assign a2288 = a856 & i20;
assign a2290 = ~a856 & l206;
assign a2292 = ~a2290 & ~a2288;
assign a2294 = ~a2292 & l86;
assign a2296 = l210 & ~l86;
assign a2298 = ~a2296 & ~a2294;
assign a2300 = ~a2298 & a916;
assign a2302 = ~a916 & l206;
assign a2304 = ~a2302 & ~a2300;
assign a2306 = l202 & l86;
assign a2308 = a2306 & ~a1350;
assign a2310 = l222 & ~l86;
assign a2312 = ~a2310 & ~a2308;
assign a2314 = ~a2312 & a860;
assign a2316 = ~a860 & l218;
assign a2318 = ~a2316 & ~a2314;
assign a2320 = l192 & l86;
assign a2322 = a2320 & ~a2176;
assign a2324 = l234 & ~l86;
assign a2326 = ~a2324 & ~a2322;
assign a2328 = ~a2326 & a860;
assign a2330 = ~a860 & l226;
assign a2332 = ~a2330 & ~a2328;
assign a2334 = a1272 & l86;
assign a2336 = a2334 & a1286;
assign a2338 = l238 & ~l86;
assign a2340 = ~a2338 & ~a2336;
assign a2342 = ~a2340 & a860;
assign a2344 = ~a860 & l230;
assign a2346 = ~a2344 & ~a2342;
assign a2348 = l142 & l86;
assign a2350 = a2348 & ~a1636;
assign a2352 = l236 & ~l86;
assign a2354 = ~a2352 & ~a2350;
assign a2356 = ~a2354 & a860;
assign a2358 = ~a860 & l232;
assign a2360 = ~a2358 & ~a2356;
assign a2362 = l250 & l248;
assign a2364 = ~a2362 & ~l256;
assign a2366 = a2364 & ~a1658;
assign a2368 = ~a2366 & l86;
assign a2370 = l258 & ~l86;
assign a2372 = ~a2370 & ~a2368;
assign a2374 = ~a2372 & a860;
assign a2376 = ~a860 & l248;
assign a2378 = ~a2376 & ~a2374;
assign a2380 = a1656 & i30;
assign a2382 = ~a2380 & ~l250;
assign a2384 = ~a1656 & i32;
assign a2386 = l86 & ~l82;
assign a2388 = a2386 & ~a2384;
assign a2390 = a2388 & ~a2382;
assign a2392 = l254 & ~l86;
assign a2394 = ~a2392 & ~a2390;
assign a2396 = ~a2394 & a860;
assign a2398 = ~a860 & l250;
assign a2400 = ~a2398 & ~a2396;
assign a2402 = a1126 & l180;
assign a2404 = ~a1308 & l112;
assign a2406 = ~a2404 & ~a2402;
assign a2408 = ~a2406 & l86;
assign a2410 = l260 & ~l86;
assign a2412 = ~a2410 & ~a2408;
assign a2414 = ~a2412 & a860;
assign a2416 = ~a860 & l256;
assign a2418 = ~a2416 & ~a2414;
assign a2420 = a2042 & l112;
assign a2422 = ~a1336 & ~a1084;
assign a2424 = ~a2422 & ~a1018;
assign a2426 = ~a1084 & l266;
assign a2428 = a2426 & a2424;
assign a2430 = ~a2428 & ~a2420;
assign a2432 = ~a2430 & l86;
assign a2434 = l342 & ~l86;
assign a2436 = ~a2434 & ~a2432;
assign a2438 = ~a2436 & a860;
assign a2440 = ~a860 & l266;
assign a2442 = ~a2440 & ~a2438;
assign a2444 = l86 & i42;
assign a2446 = l340 & ~l86;
assign a2448 = ~a2446 & ~a2444;
assign a2450 = ~a2448 & a860;
assign a2452 = ~a860 & l268;
assign a2454 = ~a2452 & ~a2450;
assign a2456 = l86 & i40;
assign a2458 = l338 & ~l86;
assign a2460 = ~a2458 & ~a2456;
assign a2462 = ~a2460 & a860;
assign a2464 = ~a860 & l270;
assign a2466 = ~a2464 & ~a2462;
assign a2468 = l86 & i38;
assign a2470 = l336 & ~l86;
assign a2472 = ~a2470 & ~a2468;
assign a2474 = ~a2472 & a860;
assign a2476 = ~a860 & l272;
assign a2478 = ~a2476 & ~a2474;
assign a2480 = l86 & i36;
assign a2482 = l334 & ~l86;
assign a2484 = ~a2482 & ~a2480;
assign a2486 = ~a2484 & a860;
assign a2488 = ~a860 & l274;
assign a2490 = ~a2488 & ~a2486;
assign a2492 = l288 & l86;
assign a2494 = l290 & ~l86;
assign a2496 = ~a2494 & ~a2492;
assign a2498 = ~a2496 & a860;
assign a2500 = ~a860 & l276;
assign a2502 = ~a2500 & ~a2498;
assign a2504 = ~a2424 & l266;
assign a2506 = l278 & ~l276;
assign a2508 = ~a2506 & ~a2504;
assign a2510 = ~a2508 & l86;
assign a2512 = l286 & ~l86;
assign a2514 = ~a2512 & ~a2510;
assign a2516 = ~a2514 & a860;
assign a2518 = ~a860 & l278;
assign a2520 = ~a2518 & ~a2516;
assign a2522 = ~a2052 & l280;
assign a2524 = ~a2522 & a1130;
assign a2526 = ~a2524 & l86;
assign a2528 = l284 & ~l86;
assign a2530 = ~a2528 & ~a2526;
assign a2532 = ~a2530 & a860;
assign a2534 = ~a860 & l280;
assign a2536 = ~a2534 & ~a2532;
assign a2538 = l292 & l86;
assign a2540 = l294 & ~l86;
assign a2542 = ~a2540 & ~a2538;
assign a2544 = ~a2542 & a860;
assign a2546 = ~a860 & l288;
assign a2548 = ~a2546 & ~a2544;
assign a2550 = l296 & l86;
assign a2552 = l298 & ~l86;
assign a2554 = ~a2552 & ~a2550;
assign a2556 = ~a2554 & a860;
assign a2558 = ~a860 & l292;
assign a2560 = ~a2558 & ~a2556;
assign a2562 = l300 & l86;
assign a2564 = l302 & ~l86;
assign a2566 = ~a2564 & ~a2562;
assign a2568 = ~a2566 & a860;
assign a2570 = ~a860 & l296;
assign a2572 = ~a2570 & ~a2568;
assign a2574 = l304 & l86;
assign a2576 = l306 & ~l86;
assign a2578 = ~a2576 & ~a2574;
assign a2580 = ~a2578 & a860;
assign a2582 = ~a860 & l300;
assign a2584 = ~a2582 & ~a2580;
assign a2586 = l308 & l86;
assign a2588 = l310 & ~l86;
assign a2590 = ~a2588 & ~a2586;
assign a2592 = ~a2590 & a860;
assign a2594 = ~a860 & l304;
assign a2596 = ~a2594 & ~a2592;
assign a2598 = l312 & l86;
assign a2600 = l314 & ~l86;
assign a2602 = ~a2600 & ~a2598;
assign a2604 = ~a2602 & a860;
assign a2606 = ~a860 & l308;
assign a2608 = ~a2606 & ~a2604;
assign a2610 = ~a1896 & ~l316;
assign a2612 = ~a2610 & l86;
assign a2614 = l318 & ~l86;
assign a2616 = ~a2614 & ~a2612;
assign a2618 = ~a2616 & a860;
assign a2620 = ~a860 & l312;
assign a2622 = ~a2620 & ~a2618;
assign a2624 = l320 & l86;
assign a2626 = l322 & ~l86;
assign a2628 = ~a2626 & ~a2624;
assign a2630 = ~a2628 & a860;
assign a2632 = ~a860 & l316;
assign a2634 = ~a2632 & ~a2630;
assign a2636 = l324 & l86;
assign a2638 = l326 & ~l86;
assign a2640 = ~a2638 & ~a2636;
assign a2642 = ~a2640 & a860;
assign a2644 = ~a860 & l320;
assign a2646 = ~a2644 & ~a2642;
assign a2648 = l328 & l86;
assign a2650 = l330 & ~l86;
assign a2652 = ~a2650 & ~a2648;
assign a2654 = ~a2652 & a860;
assign a2656 = ~a860 & l324;
assign a2658 = ~a2656 & ~a2654;
assign a2660 = a2504 & l86;
assign a2662 = l332 & ~l86;
assign a2664 = ~a2662 & ~a2660;
assign a2666 = ~a2664 & a860;
assign a2668 = ~a860 & l328;
assign a2670 = ~a2668 & ~a2666;
assign a2672 = ~l280 & ~l178;
assign a2674 = ~a2672 & a1366;
assign a2676 = l352 & l86;
assign a2678 = a2676 & a2674;
assign a2680 = l354 & ~l86;
assign a2682 = ~a2680 & ~a2678;
assign a2684 = ~a2682 & a860;
assign a2686 = ~a860 & l348;
assign a2688 = ~a2686 & ~a2684;
assign a2690 = ~a2674 & l352;
assign a2692 = a1132 & l118;
assign a2694 = ~a1210 & l112;
assign a2696 = ~a2694 & ~a2692;
assign a2698 = a2696 & ~a2690;
assign a2700 = ~a2698 & l86;
assign a2702 = l356 & ~l86;
assign a2704 = ~a2702 & ~a2700;
assign a2706 = ~a2704 & a860;
assign a2708 = ~a860 & l352;
assign a2710 = ~a2708 & ~a2706;
assign a2712 = ~a1928 & l112;
assign a2714 = a1256 & a1018;
assign a2716 = a1258 & ~l132;
assign a2718 = ~a2716 & ~a2714;
assign a2720 = a2718 & ~a1242;
assign a2722 = ~a1140 & ~l132;
assign a2724 = a2722 & ~a1238;
assign a2726 = ~a1302 & a1018;
assign a2728 = ~a1230 & a1228;
assign a2730 = ~a2728 & ~a1300;
assign a2732 = ~a2730 & ~a998;
assign a2734 = a2732 & ~l132;
assign a2736 = ~a2734 & ~a2726;
assign a2738 = a2736 & ~a2724;
assign a2740 = a2738 & a2720;
assign a2742 = ~a2740 & a2712;
assign a2744 = ~a1928 & ~l112;
assign a2746 = a2744 & l358;
assign a2748 = ~a2746 & ~a2742;
assign a2750 = ~a2748 & l86;
assign a2752 = l378 & ~l86;
assign a2754 = ~a2752 & ~a2750;
assign a2756 = ~a2754 & a860;
assign a2758 = ~a860 & l358;
assign a2760 = ~a2758 & ~a2756;
assign a2762 = a2718 & a1262;
assign a2764 = a1246 & ~l134;
assign a2766 = a2764 & ~a1244;
assign a2768 = ~a2732 & ~a2726;
assign a2770 = a2768 & ~a2766;
assign a2772 = a2770 & a2762;
assign a2774 = ~a2772 & a2712;
assign a2776 = a2744 & l360;
assign a2778 = ~a2776 & ~a2774;
assign a2780 = ~a2778 & l86;
assign a2782 = l376 & ~l86;
assign a2784 = ~a2782 & ~a2780;
assign a2786 = ~a2784 & a860;
assign a2788 = ~a860 & l360;
assign a2790 = ~a2788 & ~a2786;
assign a2792 = l370 & l270;
assign a2794 = a2792 & a1928;
assign a2796 = a2762 & ~a2724;
assign a2798 = ~a2796 & a2712;
assign a2800 = ~a2798 & ~a2794;
assign a2802 = a2744 & l362;
assign a2804 = ~a2802 & a2800;
assign a2806 = ~a2804 & l86;
assign a2808 = l372 & ~l86;
assign a2810 = ~a2808 & ~a2806;
assign a2812 = ~a2810 & a860;
assign a2814 = ~a860 & l362;
assign a2816 = ~a2814 & ~a2812;
assign a2818 = a1022 & ~a998;
assign a2820 = a2818 & a2712;
assign a2822 = a2744 & l364;
assign a2824 = ~a2822 & ~a2820;
assign a2826 = ~a2824 & l86;
assign a2828 = l368 & ~l86;
assign a2830 = ~a2828 & ~a2826;
assign a2832 = ~a2830 & a860;
assign a2834 = ~a860 & l364;
assign a2836 = ~a2834 & ~a2832;
assign a2838 = l86 & i48;
assign a2840 = l374 & ~l86;
assign a2842 = ~a2840 & ~a2838;
assign a2844 = ~a2842 & a860;
assign a2846 = ~a860 & l370;
assign a2848 = ~a2846 & ~a2844;
assign a2850 = ~a1722 & ~l148;
assign a2852 = a2850 & l398;
assign a2854 = l410 & ~l146;
assign a2856 = l404 & ~l146;
assign a2858 = l406 & ~l146;
assign a2860 = ~a2858 & ~a2856;
assign a2862 = a2860 & ~a2854;
assign a2864 = l408 & ~l146;
assign a2866 = ~a2864 & a2862;
assign a2868 = l412 & ~l146;
assign a2870 = ~a2868 & a2866;
assign a2872 = l414 & ~l146;
assign a2874 = ~a2872 & a2870;
assign a2876 = l398 & ~l146;
assign a2878 = ~a2876 & a2874;
assign a2880 = a2876 & ~a2874;
assign a2882 = ~a2880 & ~a2878;
assign a2884 = ~a2882 & ~a2850;
assign a2886 = ~a2884 & ~a2852;
assign a2888 = ~a2886 & l86;
assign a2890 = l434 & ~l86;
assign a2892 = ~a2890 & ~a2888;
assign a2894 = ~a2892 & a860;
assign a2896 = ~a860 & l398;
assign a2898 = ~a2896 & ~a2894;
assign a2900 = a2850 & l400;
assign a2902 = l400 & ~l146;
assign a2904 = ~a2902 & a2878;
assign a2906 = a2902 & ~a2878;
assign a2908 = ~a2906 & ~a2904;
assign a2910 = ~a2908 & ~a2850;
assign a2912 = ~a2910 & ~a2900;
assign a2914 = ~a2912 & l86;
assign a2916 = l432 & ~l86;
assign a2918 = ~a2916 & ~a2914;
assign a2920 = ~a2918 & a860;
assign a2922 = ~a860 & l400;
assign a2924 = ~a2922 & ~a2920;
assign a2926 = a2850 & l402;
assign a2928 = l402 & ~l146;
assign a2930 = a2928 & ~a2904;
assign a2932 = ~a2928 & a2904;
assign a2934 = ~a2932 & ~a2930;
assign a2936 = ~a2934 & ~a2850;
assign a2938 = ~a2936 & ~a2926;
assign a2940 = ~a2938 & l86;
assign a2942 = l430 & ~l86;
assign a2944 = ~a2942 & ~a2940;
assign a2946 = ~a2944 & a860;
assign a2948 = ~a860 & l402;
assign a2950 = ~a2948 & ~a2946;
assign a2952 = a2850 & l404;
assign a2954 = a2856 & l406;
assign a2956 = ~a2954 & ~a2860;
assign a2958 = ~a2956 & ~a2850;
assign a2960 = ~a2958 & ~a2952;
assign a2962 = ~a2960 & l86;
assign a2964 = l428 & ~l86;
assign a2966 = ~a2964 & ~a2962;
assign a2968 = ~a2966 & a860;
assign a2970 = ~a860 & l404;
assign a2972 = ~a2970 & ~a2968;
assign a2974 = a2850 & l406;
assign a2976 = ~a2858 & ~a2850;
assign a2978 = ~a2976 & ~a2974;
assign a2980 = ~a2978 & l86;
assign a2982 = l426 & ~l86;
assign a2984 = ~a2982 & ~a2980;
assign a2986 = ~a2984 & a860;
assign a2988 = ~a860 & l406;
assign a2990 = ~a2988 & ~a2986;
assign a2992 = a2850 & l408;
assign a2994 = a2864 & ~a2862;
assign a2996 = ~a2994 & ~a2866;
assign a2998 = ~a2996 & ~a2850;
assign a3000 = ~a2998 & ~a2992;
assign a3002 = ~a3000 & l86;
assign a3004 = l424 & ~l86;
assign a3006 = ~a3004 & ~a3002;
assign a3008 = ~a3006 & a860;
assign a3010 = ~a860 & l408;
assign a3012 = ~a3010 & ~a3008;
assign a3014 = a2850 & l410;
assign a3016 = ~a2860 & a2854;
assign a3018 = ~a3016 & ~a2862;
assign a3020 = ~a3018 & ~a2850;
assign a3022 = ~a3020 & ~a3014;
assign a3024 = ~a3022 & l86;
assign a3026 = l422 & ~l86;
assign a3028 = ~a3026 & ~a3024;
assign a3030 = ~a3028 & a860;
assign a3032 = ~a860 & l410;
assign a3034 = ~a3032 & ~a3030;
assign a3036 = a2850 & l412;
assign a3038 = a2868 & ~a2866;
assign a3040 = ~a3038 & ~a2870;
assign a3042 = ~a3040 & ~a2850;
assign a3044 = ~a3042 & ~a3036;
assign a3046 = ~a3044 & l86;
assign a3048 = l420 & ~l86;
assign a3050 = ~a3048 & ~a3046;
assign a3052 = ~a3050 & a860;
assign a3054 = ~a860 & l412;
assign a3056 = ~a3054 & ~a3052;
assign a3058 = a2850 & l414;
assign a3060 = a2872 & ~a2870;
assign a3062 = ~a3060 & ~a2874;
assign a3064 = ~a3062 & ~a2850;
assign a3066 = ~a3064 & ~a3058;
assign a3068 = ~a3066 & l86;
assign a3070 = l418 & ~l86;
assign a3072 = ~a3070 & ~a3068;
assign a3074 = ~a3072 & a860;
assign a3076 = ~a860 & l414;
assign a3078 = ~a3076 & ~a3074;
assign a3080 = ~l486 & ~l86;
assign a3082 = ~a828 & l488;
assign a3084 = l492 & l490;
assign a3086 = ~a3084 & l86;
assign a3088 = a3086 & a3082;
assign a3092 = a3090 & a832;
assign a3094 = ~a832 & l470;
assign a3096 = ~a3094 & ~a3092;
assign a3098 = a828 & i10;
assign a3100 = ~a828 & l472;
assign a3102 = ~a3100 & ~a3098;
assign a3104 = ~a3102 & l86;
assign a3106 = l484 & ~l86;
assign a3108 = ~a3106 & ~a3104;
assign a3110 = ~a3108 & a916;
assign a3112 = ~a916 & l472;
assign a3114 = ~a3112 & ~a3110;
assign a3116 = a828 & i6;
assign a3118 = ~a828 & l474;
assign a3120 = ~a3118 & ~a3116;
assign a3122 = ~a3120 & l86;
assign a3124 = l482 & ~l86;
assign a3126 = ~a3124 & ~a3122;
assign a3128 = ~a3126 & a916;
assign a3130 = ~a916 & l474;
assign a3132 = ~a3130 & ~a3128;
assign a3134 = a828 & i8;
assign a3136 = ~a828 & l476;
assign a3138 = ~a3136 & ~a3134;
assign a3140 = ~a3138 & l86;
assign a3142 = l480 & ~l86;
assign a3144 = ~a3142 & ~a3140;
assign a3146 = ~a3144 & a916;
assign a3148 = ~a916 & l476;
assign a3150 = ~a3148 & ~a3146;
assign a3152 = ~a972 & a832;
assign a3154 = ~a832 & l488;
assign a3156 = ~a3154 & ~a3152;
assign a3158 = ~l508 & ~l506;
assign a3160 = a3158 & ~l504;
assign a3162 = a3160 & ~l502;
assign a3164 = a3162 & l500;
assign a3166 = l510 & ~l500;
assign a3168 = a3166 & a3162;
assign a3170 = ~l510 & ~l500;
assign a3172 = a3170 & a3160;
assign a3174 = ~a3172 & ~a3168;
assign a3176 = a3174 & ~a3164;
assign a3178 = ~l476 & l472;
assign a3180 = l512 & l474;
assign a3182 = ~a3180 & a3178;
assign a3184 = a3182 & ~a3176;
assign a3186 = a836 & l514;
assign a3188 = a3186 & ~l512;
assign a3190 = a3188 & a3164;
assign a3192 = ~a3190 & ~a3184;
assign a3194 = ~l530 & ~l520;
assign a3196 = a3194 & ~l528;
assign a3198 = ~a3196 & ~l526;
assign a3200 = ~l538 & l536;
assign a3202 = a3200 & ~l534;
assign a3204 = a3202 & ~l532;
assign a3206 = ~l538 & ~l536;
assign a3208 = l540 & l532;
assign a3210 = a3208 & ~l534;
assign a3212 = a3210 & a3206;
assign a3214 = ~a3212 & ~a3204;
assign a3216 = ~l508 & l506;
assign a3218 = a3216 & ~l504;
assign a3220 = a3218 & a3170;
assign a3222 = a3220 & ~l502;
assign a3224 = a3222 & ~a3214;
assign a3226 = ~l540 & l532;
assign a3228 = a3206 & l534;
assign a3230 = ~a3228 & ~a3202;
assign a3232 = ~a3230 & a3226;
assign a3234 = a3232 & ~a3176;
assign a3236 = ~a3234 & ~a3224;
assign a3238 = a3236 & a3198;
assign a3240 = ~a3222 & a3176;
assign a3242 = ~a3240 & a3178;
assign a3244 = a3242 & a3238;
assign a3246 = a3244 & l524;
assign a3248 = l522 & ~l490;
assign a3250 = l542 & i14;
assign a3252 = ~a3250 & ~a3248;
assign a3254 = ~a3188 & ~l472;
assign a3256 = ~a3254 & a3222;
assign a3258 = ~a3256 & a3176;
assign a3260 = a3258 & l494;
assign a3262 = ~a3260 & a3252;
assign a3264 = a3262 & ~a3246;
assign a3266 = a3264 & ~l522;
assign a3268 = ~a3266 & l520;
assign a3270 = a3268 & l518;
assign a3272 = a3270 & l544;
assign a3274 = a3272 & l516;
assign a3276 = a3272 & l546;
assign a3278 = ~a3276 & ~a3274;
assign a3280 = ~a3278 & ~a3192;
assign a3282 = l498 & ~l490;
assign a3284 = a3282 & ~a3280;
assign a3286 = l550 & l548;
assign a3288 = l476 & l472;
assign a3290 = a3180 & a3178;
assign a3292 = ~a3290 & ~a3288;
assign a3294 = a3186 & ~a3174;
assign a3296 = ~a3294 & a3292;
assign a3298 = ~a3296 & ~a3176;
assign a3300 = l510 & l500;
assign a3302 = a3300 & ~l502;
assign a3304 = a3158 & l504;
assign a3306 = a3304 & a3302;
assign a3308 = a3304 & l502;
assign a3310 = l508 & l504;
assign a3312 = a3310 & ~l506;
assign a3314 = a3312 & ~l500;
assign a3316 = ~l552 & ~l510;
assign a3318 = a3316 & l502;
assign a3320 = ~a3318 & a3314;
assign a3322 = ~a3320 & ~a3308;
assign a3324 = a3322 & ~a3306;
assign a3326 = ~l476 & ~l472;
assign a3328 = ~l514 & l474;
assign a3330 = a3328 & a3326;
assign a3332 = a3218 & l502;
assign a3334 = a3332 & a3300;
assign a3336 = a3308 & ~a3300;
assign a3338 = ~a3336 & ~a3334;
assign a3340 = ~a3338 & a3330;
assign a3342 = a3330 & l510;
assign a3344 = a3332 & l500;
assign a3346 = a3344 & ~a3342;
assign a3348 = a3300 & l502;
assign a3350 = a3348 & a3312;
assign a3352 = ~a3350 & ~a3220;
assign a3354 = a3352 & ~a3346;
assign a3356 = a3354 & ~a3340;
assign a3358 = a3356 & a3324;
assign a3360 = a3358 & ~a3298;
assign a3362 = a3360 & l494;
assign a3364 = ~a3362 & ~a3286;
assign a3366 = a3364 & ~a3284;
assign a3368 = a3366 & ~l498;
assign a3370 = l554 & l86;
assign a3372 = a3370 & a3268;
assign a3374 = a3372 & ~a3368;
assign a3376 = a3288 & ~l474;
assign a3378 = a3376 & ~l514;
assign a3380 = a3168 & ~l182;
assign a3382 = a3380 & a3378;
assign a3384 = ~a3330 & a3308;
assign a3386 = ~a3384 & ~a3382;
assign a3388 = a3386 & a3354;
assign a3390 = l512 & l472;
assign a3392 = a3390 & ~a3388;
assign a3394 = a3178 & ~l474;
assign a3396 = a3394 & l514;
assign a3398 = a3396 & ~a3176;
assign a3400 = a3178 & l474;
assign a3402 = ~a3400 & ~a3376;
assign a3404 = ~a3176 & l514;
assign a3406 = a3404 & ~a3402;
assign a3408 = a3406 & l512;
assign a3410 = ~a3408 & ~a3398;
assign a3412 = a3410 & ~a3392;
assign a3414 = ~a3412 & l516;
assign a3416 = ~a3396 & ~a3340;
assign a3418 = ~a3416 & ~l516;
assign a3420 = ~a3418 & ~a3414;
assign a3422 = a3420 & l540;
assign a3424 = ~a3422 & ~l532;
assign a3426 = a3200 & l534;
assign a3428 = a3426 & ~a3208;
assign a3430 = a3428 & ~a3424;
assign a3432 = a3198 & l558;
assign a3434 = a3432 & ~a3430;
assign a3436 = a3434 & ~a3420;
assign a3438 = ~a3274 & ~l490;
assign a3440 = a3438 & l556;
assign a3442 = l560 & i18;
assign a3444 = a3288 & l562;
assign a3446 = ~a3444 & ~a3178;
assign a3448 = ~a3446 & a3328;
assign a3450 = ~a3394 & ~a3378;
assign a3452 = a3450 & ~a3448;
assign a3454 = ~a3452 & ~a3322;
assign a3456 = ~a3454 & ~a3340;
assign a3458 = a3456 & l494;
assign a3460 = ~a3458 & ~a3442;
assign a3462 = a3460 & ~a3440;
assign a3464 = a3462 & ~a3436;
assign a3466 = a3464 & ~l556;
assign a3468 = a3246 & l566;
assign a3470 = l564 & ~l490;
assign a3472 = l570 & l568;
assign a3474 = ~a3472 & ~a3470;
assign a3476 = a3454 & ~a3396;
assign a3478 = ~a3476 & a3258;
assign a3480 = a3478 & l494;
assign a3482 = ~a3480 & a3474;
assign a3484 = a3482 & ~a3468;
assign a3486 = a3484 & ~l564;
assign a3488 = ~a3420 & a3392;
assign a3490 = ~a3488 & a3274;
assign a3492 = ~a3490 & ~a3276;
assign a3494 = l518 & ~l490;
assign a3496 = a3494 & a3492;
assign a3498 = l574 & l572;
assign a3500 = ~l580 & ~l578;
assign a3502 = a3500 & l576;
assign a3504 = ~a3502 & ~a3498;
assign a3506 = a3388 & ~a3320;
assign a3508 = a3506 & l494;
assign a3510 = ~a3508 & a3504;
assign a3512 = a3510 & ~a3496;
assign a3514 = a3512 & ~l518;
assign a3516 = ~a3514 & ~a3486;
assign a3518 = a3516 & ~a3466;
assign a3520 = a3518 & a3374;
assign a3522 = l582 & ~l86;
assign a3524 = ~a3522 & ~a3520;
assign a3526 = ~a3524 & a832;
assign a3528 = ~a832 & l490;
assign a3530 = ~a3528 & ~a3526;
assign a3532 = l492 & ~l490;
assign a3534 = ~a3532 & ~l494;
assign a3536 = ~a3534 & l86;
assign a3538 = l496 & ~l86;
assign a3540 = ~a3538 & ~a3536;
assign a3542 = ~a3540 & a832;
assign a3544 = ~a832 & l492;
assign a3546 = ~a3544 & ~a3542;
assign a3548 = ~a832 & l494;
assign a3550 = ~a3548 & ~a1404;
assign a3552 = ~a3366 & l86;
assign a3554 = l818 & ~l86;
assign a3556 = ~a3554 & ~a3552;
assign a3558 = ~a3556 & a832;
assign a3560 = ~a832 & l498;
assign a3562 = ~a3560 & ~a3558;
assign a3564 = a1430 & a828;
assign a3566 = ~a828 & l500;
assign a3568 = ~a3566 & ~a3564;
assign a3570 = ~a3568 & l86;
assign a3572 = l816 & ~l86;
assign a3574 = ~a3572 & ~a3570;
assign a3576 = ~a3574 & a916;
assign a3578 = ~a916 & l500;
assign a3580 = ~a3578 & ~a3576;
assign a3582 = a828 & i74;
assign a3584 = ~a828 & l502;
assign a3586 = ~a3584 & ~a3582;
assign a3588 = ~a3586 & l86;
assign a3590 = l814 & ~l86;
assign a3592 = ~a3590 & ~a3588;
assign a3594 = ~a3592 & a916;
assign a3596 = ~a916 & l502;
assign a3598 = ~a3596 & ~a3594;
assign a3600 = a828 & i72;
assign a3602 = ~a828 & l504;
assign a3604 = ~a3602 & ~a3600;
assign a3606 = ~a3604 & l86;
assign a3608 = l812 & ~l86;
assign a3610 = ~a3608 & ~a3606;
assign a3612 = ~a3610 & a916;
assign a3614 = ~a916 & l504;
assign a3616 = ~a3614 & ~a3612;
assign a3618 = a828 & i70;
assign a3620 = ~a828 & l506;
assign a3622 = ~a3620 & ~a3618;
assign a3624 = ~a3622 & l86;
assign a3626 = l810 & ~l86;
assign a3628 = ~a3626 & ~a3624;
assign a3630 = ~a3628 & a916;
assign a3632 = ~a916 & l506;
assign a3634 = ~a3632 & ~a3630;
assign a3636 = a828 & i68;
assign a3638 = ~a828 & l508;
assign a3640 = ~a3638 & ~a3636;
assign a3642 = ~a3640 & l86;
assign a3644 = l808 & ~l86;
assign a3646 = ~a3644 & ~a3642;
assign a3648 = ~a3646 & a916;
assign a3650 = ~a916 & l508;
assign a3652 = ~a3650 & ~a3648;
assign a3654 = a828 & i66;
assign a3656 = ~a828 & l510;
assign a3658 = ~a3656 & ~a3654;
assign a3660 = ~a3658 & l86;
assign a3662 = l806 & ~l86;
assign a3664 = ~a3662 & ~a3660;
assign a3666 = ~a3664 & a916;
assign a3668 = ~a916 & l510;
assign a3670 = ~a3668 & ~a3666;
assign a3672 = a828 & i64;
assign a3674 = ~a828 & l512;
assign a3676 = ~a3674 & ~a3672;
assign a3678 = ~a3676 & l86;
assign a3680 = l804 & ~l86;
assign a3682 = ~a3680 & ~a3678;
assign a3684 = ~a3682 & a916;
assign a3686 = ~a916 & l512;
assign a3688 = ~a3686 & ~a3684;
assign a3690 = a828 & i62;
assign a3692 = ~a828 & l514;
assign a3694 = ~a3692 & ~a3690;
assign a3696 = ~a3694 & l86;
assign a3698 = l802 & ~l86;
assign a3700 = ~a3698 & ~a3696;
assign a3702 = ~a3700 & a916;
assign a3704 = ~a916 & l514;
assign a3706 = ~a3704 & ~a3702;
assign a3708 = l720 & l716;
assign a3710 = ~l718 & ~l716;
assign a3712 = ~a3710 & ~l722;
assign a3714 = a3712 & ~a3708;
assign a3716 = a3714 & ~a3258;
assign a3718 = ~a3716 & l644;
assign a3720 = ~l644 & ~l516;
assign a3722 = ~a3720 & a3086;
assign a3724 = a3722 & ~a3718;
assign a3726 = l800 & ~l86;
assign a3728 = ~a3726 & ~a3724;
assign a3730 = ~a3728 & a832;
assign a3732 = ~a832 & l516;
assign a3734 = ~a3732 & ~a3730;
assign a3736 = ~a3512 & l86;
assign a3738 = l798 & ~l86;
assign a3740 = ~a3738 & ~a3736;
assign a3742 = ~a3740 & a832;
assign a3744 = ~a832 & l518;
assign a3746 = ~a3744 & ~a3742;
assign a3748 = a3438 & l520;
assign a3750 = ~l752 & ~l750;
assign a3752 = ~l756 & ~l754;
assign a3754 = a3752 & a3750;
assign a3756 = ~l760 & ~l758;
assign a3758 = ~l764 & ~l762;
assign a3760 = a3758 & ~l766;
assign a3762 = a3760 & a3756;
assign a3764 = a3762 & a3754;
assign a3766 = a3764 & l530;
assign a3768 = l502 & l476;
assign a3770 = ~a3768 & a3220;
assign a3772 = ~a3770 & ~a3346;
assign a3774 = ~a3772 & l472;
assign a3776 = ~a3774 & a3176;
assign a3778 = a3776 & a3456;
assign a3780 = a3778 & l494;
assign a3782 = ~a3780 & ~a3766;
assign a3784 = a3782 & ~a3748;
assign a3786 = ~a3784 & l86;
assign a3788 = l796 & ~l86;
assign a3790 = ~a3788 & ~a3786;
assign a3792 = ~a3790 & a832;
assign a3794 = ~a832 & l520;
assign a3796 = ~a3794 & ~a3792;
assign a3798 = ~a3264 & l86;
assign a3800 = l794 & ~l86;
assign a3802 = ~a3800 & ~a3798;
assign a3804 = ~a3802 & a832;
assign a3806 = ~a832 & l522;
assign a3808 = ~a3806 & ~a3804;
assign a3810 = ~a3258 & l494;
assign a3812 = ~a3236 & a3198;
assign a3814 = ~a3812 & a3242;
assign a3816 = a3814 & l524;
assign a3818 = a3816 & ~a3244;
assign a3820 = ~a3818 & ~a3810;
assign a3822 = ~a3820 & l86;
assign a3824 = l792 & ~l86;
assign a3826 = ~a3824 & ~a3822;
assign a3828 = ~a3826 & a832;
assign a3830 = ~a832 & l524;
assign a3832 = ~a3830 & ~a3828;
assign a3834 = a3430 & a3198;
assign a3836 = a3834 & l558;
assign a3838 = a3836 & l528;
assign a3840 = ~l600 & ~l560;
assign a3842 = ~l626 & ~l618;
assign a3844 = a3842 & a3840;
assign a3846 = ~a3844 & ~l558;
assign a3848 = ~a3846 & l526;
assign a3850 = a3848 & i50;
assign a3852 = ~a3850 & l526;
assign a3854 = ~a3778 & l494;
assign a3856 = ~a3854 & ~a3852;
assign a3858 = a3856 & ~a3274;
assign a3860 = a3858 & ~a3838;
assign a3862 = ~a3860 & l86;
assign a3864 = l790 & ~l86;
assign a3866 = ~a3864 & ~a3862;
assign a3868 = ~a3866 & a832;
assign a3870 = ~a832 & l526;
assign a3872 = ~a3870 & ~a3868;
assign a3874 = a3848 & a1708;
assign a3876 = l788 & ~l86;
assign a3878 = ~a3876 & ~a3874;
assign a3880 = ~a3878 & a832;
assign a3882 = ~a832 & l528;
assign a3884 = ~a3882 & ~a3880;
assign a3886 = ~a3836 & l528;
assign a3888 = ~a3764 & l530;
assign a3890 = ~a3888 & ~a3886;
assign a3892 = ~a3890 & l86;
assign a3894 = l768 & ~l86;
assign a3896 = ~a3894 & ~a3892;
assign a3898 = ~a3896 & a832;
assign a3900 = ~a832 & l530;
assign a3902 = ~a3900 & ~a3898;
assign a3904 = a3850 & i60;
assign a3906 = ~a3850 & l532;
assign a3908 = ~a3906 & ~a3904;
assign a3910 = ~a3908 & l86;
assign a3912 = l748 & ~l86;
assign a3914 = ~a3912 & ~a3910;
assign a3916 = ~a3914 & a832;
assign a3918 = ~a832 & l532;
assign a3920 = ~a3918 & ~a3916;
assign a3922 = a3850 & i58;
assign a3924 = ~a3850 & l534;
assign a3926 = ~a3924 & ~a3922;
assign a3928 = ~a3926 & l86;
assign a3930 = l746 & ~l86;
assign a3932 = ~a3930 & ~a3928;
assign a3934 = ~a3932 & a832;
assign a3936 = ~a832 & l534;
assign a3938 = ~a3936 & ~a3934;
assign a3940 = a3850 & i56;
assign a3942 = ~a3850 & l536;
assign a3944 = ~a3942 & ~a3940;
assign a3946 = ~a3944 & l86;
assign a3948 = l744 & ~l86;
assign a3950 = ~a3948 & ~a3946;
assign a3952 = ~a3950 & a832;
assign a3954 = ~a832 & l536;
assign a3956 = ~a3954 & ~a3952;
assign a3958 = a3850 & i54;
assign a3960 = ~a3850 & l538;
assign a3962 = ~a3960 & ~a3958;
assign a3964 = ~a3962 & l86;
assign a3966 = l742 & ~l86;
assign a3968 = ~a3966 & ~a3964;
assign a3970 = ~a3968 & a832;
assign a3972 = ~a832 & l538;
assign a3974 = ~a3972 & ~a3970;
assign a3976 = a3850 & i52;
assign a3978 = ~a3850 & l540;
assign a3980 = ~a3978 & ~a3976;
assign a3982 = ~a3980 & l86;
assign a3984 = l740 & ~l86;
assign a3986 = ~a3984 & ~a3982;
assign a3988 = ~a3986 & a832;
assign a3990 = ~a832 & l540;
assign a3992 = ~a3990 & ~a3988;
assign a3994 = l542 & ~i14;
assign a3996 = ~a3994 & ~l602;
assign a3998 = ~a3996 & l86;
assign a4000 = l738 & ~l86;
assign a4002 = ~a4000 & ~a3998;
assign a4004 = ~a4002 & a832;
assign a4006 = ~a832 & l542;
assign a4008 = ~a4006 & ~a4004;
assign a4010 = ~a3456 & l638;
assign a4012 = ~l642 & ~l638;
assign a4014 = a4012 & ~l640;
assign a4016 = ~a4014 & ~a3258;
assign a4018 = ~a4016 & ~a4010;
assign a4020 = l646 & l644;
assign a4022 = a4020 & ~a4018;
assign a4024 = ~l546 & ~l516;
assign a4026 = ~a4024 & l544;
assign a4028 = a4026 & ~a3270;
assign a4030 = ~a4028 & ~a4022;
assign a4032 = ~a4030 & l86;
assign a4034 = l736 & ~l86;
assign a4036 = ~a4034 & ~a4032;
assign a4038 = ~a4036 & a832;
assign a4040 = ~a832 & l544;
assign a4042 = ~a4040 & ~a4038;
assign a4044 = l722 & ~l720;
assign a4046 = a4044 & a3710;
assign a4048 = ~l722 & l718;
assign a4050 = a4048 & a3708;
assign a4052 = ~a4050 & ~a4046;
assign a4054 = ~a4052 & ~a3258;
assign a4056 = a3186 & a3164;
assign a4058 = ~a4056 & l644;
assign a4060 = a4058 & ~a4054;
assign a4062 = ~l644 & ~l546;
assign a4064 = ~a4062 & a3086;
assign a4066 = a4064 & ~a4060;
assign a4068 = l724 & ~l86;
assign a4070 = ~a4068 & ~a4066;
assign a4072 = ~a4070 & a832;
assign a4074 = ~a832 & l546;
assign a4076 = ~a4074 & ~a4072;
assign a4078 = ~l550 & l548;
assign a4080 = ~a4078 & ~l706;
assign a4082 = ~a4080 & l86;
assign a4084 = l708 & ~l86;
assign a4086 = ~a4084 & ~a4082;
assign a4088 = ~a4086 & a832;
assign a4090 = ~a832 & l548;
assign a4092 = ~a4090 & ~a4088;
assign a4094 = ~a2010 & a832;
assign a4096 = ~a832 & l550;
assign a4098 = ~a4096 & ~a4094;
assign a4100 = a828 & i44;
assign a4102 = ~a828 & l552;
assign a4104 = ~a4102 & ~a4100;
assign a4106 = ~a4104 & l86;
assign a4108 = l704 & ~l86;
assign a4110 = ~a4108 & ~a4106;
assign a4112 = ~a4110 & a916;
assign a4114 = ~a916 & l552;
assign a4116 = ~a4114 & ~a4112;
assign a4118 = ~a3478 & l634;
assign a4120 = ~a4118 & l494;
assign a4122 = ~l560 & ~l556;
assign a4124 = ~a4122 & l518;
assign a4126 = a4124 & l636;
assign a4128 = l554 & ~l490;
assign a4130 = a4024 & l544;
assign a4132 = ~a4130 & ~a4128;
assign a4134 = a4132 & ~a4126;
assign a4136 = a4134 & ~a4120;
assign a4138 = a4020 & a4018;
assign a4140 = a3246 & l648;
assign a4142 = ~a4140 & ~a4138;
assign a4144 = a4142 & a4136;
assign a4146 = ~a4144 & l86;
assign a4148 = l650 & ~l86;
assign a4150 = ~a4148 & ~a4146;
assign a4152 = ~a4150 & a832;
assign a4154 = ~a832 & l554;
assign a4156 = ~a4154 & ~a4152;
assign a4158 = ~a3464 & l86;
assign a4160 = l632 & ~l86;
assign a4162 = ~a4160 & ~a4158;
assign a4164 = ~a4162 & a832;
assign a4166 = ~a832 & l556;
assign a4168 = ~a4166 & ~a4164;
assign a4170 = ~l620 & l618;
assign a4172 = ~a3198 & l558;
assign a4174 = ~a4172 & ~a4170;
assign a4176 = ~a4174 & l86;
assign a4178 = l622 & ~l86;
assign a4180 = ~a4178 & ~a4176;
assign a4182 = ~a4180 & a832;
assign a4184 = ~a832 & l558;
assign a4186 = ~a4184 & ~a4182;
assign a4188 = l560 & ~i18;
assign a4190 = ~a4188 & ~l600;
assign a4192 = ~a4190 & l86;
assign a4194 = l616 & ~l86;
assign a4196 = ~a4194 & ~a4192;
assign a4198 = ~a4196 & a832;
assign a4200 = ~a832 & l560;
assign a4202 = ~a4200 & ~a4198;
assign a4204 = a828 & i28;
assign a4206 = ~a828 & l562;
assign a4208 = ~a4206 & ~a4204;
assign a4210 = ~a4208 & l86;
assign a4212 = l614 & ~l86;
assign a4214 = ~a4212 & ~a4210;
assign a4216 = ~a4214 & a916;
assign a4218 = ~a916 & l562;
assign a4220 = ~a4218 & ~a4216;
assign a4222 = ~a3484 & l86;
assign a4224 = l612 & ~l86;
assign a4226 = ~a4224 & ~a4222;
assign a4228 = ~a4226 & a832;
assign a4230 = ~a832 & l564;
assign a4232 = ~a4230 & ~a4228;
assign a4234 = ~a3478 & l84;
assign a4236 = ~l602 & ~l600;
assign a4238 = a4236 & l566;
assign a4240 = a4238 & ~a3246;
assign a4242 = ~a4240 & ~a4234;
assign a4244 = ~a4242 & l86;
assign a4246 = l610 & ~l86;
assign a4248 = ~a4246 & ~a4244;
assign a4250 = ~a4248 & a832;
assign a4252 = ~a832 & l566;
assign a4254 = ~a4252 & ~a4250;
assign a4256 = ~l570 & l568;
assign a4258 = ~a4256 & ~l596;
assign a4260 = ~a4258 & l86;
assign a4262 = l598 & ~l86;
assign a4264 = ~a4262 & ~a4260;
assign a4266 = ~a4264 & a832;
assign a4268 = ~a832 & l568;
assign a4270 = ~a4268 & ~a4266;
assign a4272 = ~a2216 & a832;
assign a4274 = ~a832 & l570;
assign a4276 = ~a4274 & ~a4272;
assign a4278 = ~l574 & l572;
assign a4280 = ~a4278 & ~l590;
assign a4282 = ~a4280 & l86;
assign a4284 = l592 & ~l86;
assign a4286 = ~a4284 & ~a4282;
assign a4288 = ~a4286 & a832;
assign a4290 = ~a832 & l572;
assign a4292 = ~a4290 & ~a4288;
assign a4294 = ~a2244 & a832;
assign a4296 = ~a832 & l574;
assign a4298 = ~a4296 & ~a4294;
assign a4300 = ~a3506 & l494;
assign a4302 = ~a3492 & l518;
assign a4304 = ~a4302 & ~a4300;
assign a4306 = ~a4304 & l86;
assign a4308 = l588 & ~l86;
assign a4310 = ~a4308 & ~a4306;
assign a4312 = ~a4310 & a832;
assign a4314 = ~a832 & l576;
assign a4316 = ~a4314 & ~a4312;
assign a4318 = a828 & i22;
assign a4320 = ~a828 & l578;
assign a4322 = ~a4320 & ~a4318;
assign a4324 = ~a4322 & l86;
assign a4326 = l586 & ~l86;
assign a4328 = ~a4326 & ~a4324;
assign a4330 = ~a4328 & a916;
assign a4332 = ~a916 & l578;
assign a4334 = ~a4332 & ~a4330;
assign a4336 = a828 & i20;
assign a4338 = ~a828 & l580;
assign a4340 = ~a4338 & ~a4336;
assign a4342 = ~a4340 & l86;
assign a4344 = l584 & ~l86;
assign a4346 = ~a4344 & ~a4342;
assign a4348 = ~a4346 & a916;
assign a4350 = ~a916 & l580;
assign a4352 = ~a4350 & ~a4348;
assign a4354 = l576 & l86;
assign a4356 = a4354 & ~a3500;
assign a4358 = l594 & ~l86;
assign a4360 = ~a4358 & ~a4356;
assign a4362 = ~a4360 & a832;
assign a4364 = ~a832 & l590;
assign a4366 = ~a4364 & ~a4362;
assign a4368 = l566 & l86;
assign a4370 = a4368 & ~a4236;
assign a4372 = l604 & ~l86;
assign a4374 = ~a4372 & ~a4370;
assign a4376 = ~a4374 & a832;
assign a4378 = ~a832 & l596;
assign a4380 = ~a4378 & ~a4376;
assign a4382 = a3420 & l86;
assign a4384 = a4382 & a3434;
assign a4386 = l608 & ~l86;
assign a4388 = ~a4386 & ~a4384;
assign a4390 = ~a4388 & a832;
assign a4392 = ~a832 & l600;
assign a4394 = ~a4392 & ~a4390;
assign a4396 = l524 & l86;
assign a4398 = a4396 & ~a3814;
assign a4400 = l606 & ~l86;
assign a4402 = ~a4400 & ~a4398;
assign a4404 = ~a4402 & a832;
assign a4406 = ~a832 & l602;
assign a4408 = ~a4406 & ~a4404;
assign a4410 = l620 & l618;
assign a4412 = ~a4410 & ~l626;
assign a4414 = a4412 & ~a3836;
assign a4416 = ~a4414 & l86;
assign a4418 = l628 & ~l86;
assign a4420 = ~a4418 & ~a4416;
assign a4422 = ~a4420 & a832;
assign a4424 = ~a832 & l618;
assign a4426 = ~a4424 & ~a4422;
assign a4428 = a3834 & i30;
assign a4430 = ~a4428 & ~l620;
assign a4432 = ~a3834 & i32;
assign a4434 = ~l470 & l86;
assign a4436 = a4434 & ~a4432;
assign a4438 = a4436 & ~a4430;
assign a4440 = l624 & ~l86;
assign a4442 = ~a4440 & ~a4438;
assign a4444 = ~a4442 & a832;
assign a4446 = ~a832 & l620;
assign a4448 = ~a4446 & ~a4444;
assign a4450 = a3274 & l556;
assign a4452 = ~a3456 & l494;
assign a4454 = ~a4452 & ~a4450;
assign a4456 = ~a4454 & l86;
assign a4458 = l630 & ~l86;
assign a4460 = ~a4458 & ~a4456;
assign a4462 = ~a4460 & a832;
assign a4464 = ~a832 & l626;
assign a4466 = ~a4464 & ~a4462;
assign a4468 = ~a2448 & a832;
assign a4470 = ~a832 & l634;
assign a4472 = ~a4470 & ~a4468;
assign a4474 = ~a4124 & l636;
assign a4476 = ~a4474 & a3278;
assign a4478 = ~a4476 & l86;
assign a4480 = l702 & ~l86;
assign a4482 = ~a4480 & ~a4478;
assign a4484 = ~a4482 & a832;
assign a4486 = ~a832 & l636;
assign a4488 = ~a4486 & ~a4484;
assign a4490 = ~a2460 & a832;
assign a4492 = ~a832 & l638;
assign a4494 = ~a4492 & ~a4490;
assign a4496 = ~a2472 & a832;
assign a4498 = ~a832 & l640;
assign a4500 = ~a4498 & ~a4496;
assign a4502 = ~a2484 & a832;
assign a4504 = ~a832 & l642;
assign a4506 = ~a4504 & ~a4502;
assign a4508 = l656 & l86;
assign a4510 = l658 & ~l86;
assign a4512 = ~a4510 & ~a4508;
assign a4514 = ~a4512 & a832;
assign a4516 = ~a832 & l644;
assign a4518 = ~a4516 & ~a4514;
assign a4520 = ~a3246 & l648;
assign a4522 = a4520 & ~a3486;
assign a4524 = l646 & ~l644;
assign a4526 = ~a4524 & ~a4522;
assign a4528 = ~a4526 & l86;
assign a4530 = l654 & ~l86;
assign a4532 = ~a4530 & ~a4528;
assign a4534 = ~a4532 & a832;
assign a4536 = ~a832 & l646;
assign a4538 = ~a4536 & ~a4534;
assign a4540 = a4118 & l494;
assign a4542 = a4520 & a3486;
assign a4544 = ~a4542 & ~a4540;
assign a4546 = ~a4544 & l86;
assign a4548 = l652 & ~l86;
assign a4550 = ~a4548 & ~a4546;
assign a4552 = ~a4550 & a832;
assign a4554 = ~a832 & l648;
assign a4556 = ~a4554 & ~a4552;
assign a4558 = l660 & l86;
assign a4560 = l662 & ~l86;
assign a4562 = ~a4560 & ~a4558;
assign a4564 = ~a4562 & a832;
assign a4566 = ~a832 & l656;
assign a4568 = ~a4566 & ~a4564;
assign a4570 = l664 & l86;
assign a4572 = l666 & ~l86;
assign a4574 = ~a4572 & ~a4570;
assign a4576 = ~a4574 & a832;
assign a4578 = ~a832 & l660;
assign a4580 = ~a4578 & ~a4576;
assign a4582 = l668 & l86;
assign a4584 = l670 & ~l86;
assign a4586 = ~a4584 & ~a4582;
assign a4588 = ~a4586 & a832;
assign a4590 = ~a832 & l664;
assign a4592 = ~a4590 & ~a4588;
assign a4594 = l672 & l86;
assign a4596 = l674 & ~l86;
assign a4598 = ~a4596 & ~a4594;
assign a4600 = ~a4598 & a832;
assign a4602 = ~a832 & l668;
assign a4604 = ~a4602 & ~a4600;
assign a4606 = l676 & l86;
assign a4608 = l678 & ~l86;
assign a4610 = ~a4608 & ~a4606;
assign a4612 = ~a4610 & a832;
assign a4614 = ~a832 & l672;
assign a4616 = ~a4614 & ~a4612;
assign a4618 = l680 & l86;
assign a4620 = l682 & ~l86;
assign a4622 = ~a4620 & ~a4618;
assign a4624 = ~a4622 & a832;
assign a4626 = ~a832 & l676;
assign a4628 = ~a4626 & ~a4624;
assign a4630 = l684 & l86;
assign a4632 = l686 & ~l86;
assign a4634 = ~a4632 & ~a4630;
assign a4636 = ~a4634 & a832;
assign a4638 = ~a832 & l680;
assign a4640 = ~a4638 & ~a4636;
assign a4642 = l688 & l86;
assign a4644 = l690 & ~l86;
assign a4646 = ~a4644 & ~a4642;
assign a4648 = ~a4646 & a832;
assign a4650 = ~a832 & l684;
assign a4652 = ~a4650 & ~a4648;
assign a4654 = l692 & l86;
assign a4656 = l694 & ~l86;
assign a4658 = ~a4656 & ~a4654;
assign a4660 = ~a4658 & a832;
assign a4662 = ~a832 & l688;
assign a4664 = ~a4662 & ~a4660;
assign a4666 = l696 & l86;
assign a4668 = l698 & ~l86;
assign a4670 = ~a4668 & ~a4666;
assign a4672 = ~a4670 & a832;
assign a4674 = ~a832 & l692;
assign a4676 = ~a4674 & ~a4672;
assign a4678 = a4522 & l86;
assign a4680 = l700 & ~l86;
assign a4682 = ~a4680 & ~a4678;
assign a4684 = ~a4682 & a832;
assign a4686 = ~a832 & l696;
assign a4688 = ~a4686 & ~a4684;
assign a4690 = ~l636 & ~l554;
assign a4692 = ~a4690 & a3516;
assign a4694 = l710 & l86;
assign a4696 = a4694 & a4692;
assign a4698 = l712 & ~l86;
assign a4700 = ~a4698 & ~a4696;
assign a4702 = ~a4700 & a832;
assign a4704 = ~a832 & l706;
assign a4706 = ~a4704 & ~a4702;
assign a4708 = ~a4692 & l710;
assign a4710 = a3280 & l498;
assign a4712 = ~a3360 & l494;
assign a4714 = ~a4712 & ~a4710;
assign a4716 = a4714 & ~a4708;
assign a4718 = ~a4716 & l86;
assign a4720 = l714 & ~l86;
assign a4722 = ~a4720 & ~a4718;
assign a4724 = ~a4722 & a832;
assign a4726 = ~a832 & l710;
assign a4728 = ~a4726 & ~a4724;
assign a4730 = ~a4022 & l494;
assign a4732 = ~a3380 & a3378;
assign a4734 = ~a4732 & ~a3448;
assign a4736 = ~a4734 & ~a3176;
assign a4738 = a4736 & ~l512;
assign a4740 = ~a4738 & ~a3392;
assign a4742 = ~a3326 & ~l512;
assign a4744 = a4742 & ~a3388;
assign a4746 = a3406 & ~l512;
assign a4748 = ~a4746 & ~a4744;
assign a4750 = a4748 & a4740;
assign a4752 = ~a4750 & a4730;
assign a4754 = ~a4022 & ~l494;
assign a4756 = a4754 & l716;
assign a4758 = ~a4756 & ~a4752;
assign a4760 = ~a4758 & l86;
assign a4762 = l734 & ~l86;
assign a4764 = ~a4762 & ~a4760;
assign a4766 = ~a4764 & a832;
assign a4768 = ~a832 & l716;
assign a4770 = ~a4768 & ~a4766;
assign a4772 = ~a4746 & a3410;
assign a4774 = a3394 & ~l514;
assign a4776 = a4774 & ~a3176;
assign a4778 = ~a4776 & ~a4736;
assign a4780 = a4778 & a4772;
assign a4782 = ~a4780 & a4730;
assign a4784 = a4754 & l718;
assign a4786 = ~a4784 & ~a4782;
assign a4788 = ~a4786 & l86;
assign a4790 = l732 & ~l86;
assign a4792 = ~a4790 & ~a4788;
assign a4794 = ~a4792 & a832;
assign a4796 = ~a832 & l718;
assign a4798 = ~a4796 & ~a4794;
assign a4800 = l728 & l638;
assign a4802 = a4800 & a4022;
assign a4804 = a4772 & ~a4744;
assign a4806 = ~a4804 & a4730;
assign a4808 = ~a4806 & ~a4802;
assign a4810 = a4754 & l720;
assign a4812 = ~a4810 & a4808;
assign a4814 = ~a4812 & l86;
assign a4816 = l730 & ~l86;
assign a4818 = ~a4816 & ~a4814;
assign a4820 = ~a4818 & a832;
assign a4822 = ~a832 & l720;
assign a4824 = ~a4822 & ~a4820;
assign a4826 = a3404 & a836;
assign a4828 = a4826 & a4730;
assign a4830 = a4754 & l722;
assign a4832 = ~a4830 & ~a4828;
assign a4834 = ~a4832 & l86;
assign a4836 = l726 & ~l86;
assign a4838 = ~a4836 & ~a4834;
assign a4840 = ~a4838 & a832;
assign a4842 = ~a832 & l722;
assign a4844 = ~a4842 & ~a4840;
assign a4846 = ~a2842 & a832;
assign a4848 = ~a832 & l728;
assign a4850 = ~a4848 & ~a4846;
assign a4852 = ~a3886 & ~l530;
assign a4854 = a4852 & l750;
assign a4856 = l762 & ~l528;
assign a4858 = l756 & ~l528;
assign a4860 = l758 & ~l528;
assign a4862 = ~a4860 & ~a4858;
assign a4864 = a4862 & ~a4856;
assign a4866 = l760 & ~l528;
assign a4868 = ~a4866 & a4864;
assign a4870 = l764 & ~l528;
assign a4872 = ~a4870 & a4868;
assign a4874 = l766 & ~l528;
assign a4876 = ~a4874 & a4872;
assign a4878 = l750 & ~l528;
assign a4880 = ~a4878 & a4876;
assign a4882 = a4878 & ~a4876;
assign a4884 = ~a4882 & ~a4880;
assign a4886 = ~a4884 & ~a4852;
assign a4888 = ~a4886 & ~a4854;
assign a4890 = ~a4888 & l86;
assign a4892 = l786 & ~l86;
assign a4894 = ~a4892 & ~a4890;
assign a4896 = ~a4894 & a832;
assign a4898 = ~a832 & l750;
assign a4900 = ~a4898 & ~a4896;
assign a4902 = a4852 & l752;
assign a4904 = l752 & ~l528;
assign a4906 = ~a4904 & a4880;
assign a4908 = a4904 & ~a4880;
assign a4910 = ~a4908 & ~a4906;
assign a4912 = ~a4910 & ~a4852;
assign a4914 = ~a4912 & ~a4902;
assign a4916 = ~a4914 & l86;
assign a4918 = l784 & ~l86;
assign a4920 = ~a4918 & ~a4916;
assign a4922 = ~a4920 & a832;
assign a4924 = ~a832 & l752;
assign a4926 = ~a4924 & ~a4922;
assign a4928 = a4852 & l754;
assign a4930 = l754 & ~l528;
assign a4932 = a4930 & ~a4906;
assign a4934 = ~a4930 & a4906;
assign a4936 = ~a4934 & ~a4932;
assign a4938 = ~a4936 & ~a4852;
assign a4940 = ~a4938 & ~a4928;
assign a4942 = ~a4940 & l86;
assign a4944 = l782 & ~l86;
assign a4946 = ~a4944 & ~a4942;
assign a4948 = ~a4946 & a832;
assign a4950 = ~a832 & l754;
assign a4952 = ~a4950 & ~a4948;
assign a4954 = a4852 & l756;
assign a4956 = a4858 & l758;
assign a4958 = ~a4956 & ~a4862;
assign a4960 = ~a4958 & ~a4852;
assign a4962 = ~a4960 & ~a4954;
assign a4964 = ~a4962 & l86;
assign a4966 = l780 & ~l86;
assign a4968 = ~a4966 & ~a4964;
assign a4970 = ~a4968 & a832;
assign a4972 = ~a832 & l756;
assign a4974 = ~a4972 & ~a4970;
assign a4976 = a4852 & l758;
assign a4978 = ~a4860 & ~a4852;
assign a4980 = ~a4978 & ~a4976;
assign a4982 = ~a4980 & l86;
assign a4984 = l778 & ~l86;
assign a4986 = ~a4984 & ~a4982;
assign a4988 = ~a4986 & a832;
assign a4990 = ~a832 & l758;
assign a4992 = ~a4990 & ~a4988;
assign a4994 = a4852 & l760;
assign a4996 = a4866 & ~a4864;
assign a4998 = ~a4996 & ~a4868;
assign a5000 = ~a4998 & ~a4852;
assign a5002 = ~a5000 & ~a4994;
assign a5004 = ~a5002 & l86;
assign a5006 = l776 & ~l86;
assign a5008 = ~a5006 & ~a5004;
assign a5010 = ~a5008 & a832;
assign a5012 = ~a832 & l760;
assign a5014 = ~a5012 & ~a5010;
assign a5016 = a4852 & l762;
assign a5018 = ~a4862 & a4856;
assign a5020 = ~a5018 & ~a4864;
assign a5022 = ~a5020 & ~a4852;
assign a5024 = ~a5022 & ~a5016;
assign a5026 = ~a5024 & l86;
assign a5028 = l774 & ~l86;
assign a5030 = ~a5028 & ~a5026;
assign a5032 = ~a5030 & a832;
assign a5034 = ~a832 & l762;
assign a5036 = ~a5034 & ~a5032;
assign a5038 = a4852 & l764;
assign a5040 = a4870 & ~a4868;
assign a5042 = ~a5040 & ~a4872;
assign a5044 = ~a5042 & ~a4852;
assign a5046 = ~a5044 & ~a5038;
assign a5048 = ~a5046 & l86;
assign a5050 = l772 & ~l86;
assign a5052 = ~a5050 & ~a5048;
assign a5054 = ~a5052 & a832;
assign a5056 = ~a832 & l764;
assign a5058 = ~a5056 & ~a5054;
assign a5060 = a4852 & l766;
assign a5062 = a4874 & ~a4872;
assign a5064 = ~a5062 & ~a4876;
assign a5066 = ~a5064 & ~a4852;
assign a5068 = ~a5066 & ~a5060;
assign a5070 = ~a5068 & l86;
assign a5072 = l770 & ~l86;
assign a5074 = ~a5072 & ~a5070;
assign a5076 = ~a5074 & a832;
assign a5078 = ~a832 & l766;
assign a5080 = ~a5078 & ~a5076;
assign p0 = ~a826;

assert property (~p0);

endmodule
