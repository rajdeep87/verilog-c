module m6s13 (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474,i476,i478,i480,
i482,i484,i486,i488,i490,i492,i494,i496,i498,i500,i502,i504,i506,i508,i510,
i512,i514,i516,i518,i520,i522,i524,i526,i528,i530,i532,i534,i536,i538,i540,
i542,i544,i546,i548,i550,i552,i554,i556,i558,i560,i562,i564,i566,i568,i570,
i572,i574,i576,i578,i580,i582,i584,i586,i588,i590,i592,i594,i596,i598,i600,
i602,i604,i606,i608,i610,i612,i614,i616,i618,i620,i622,i624,i626,i628,i630,
i632,i634,i636,i638,i640,i642,i644,i646,i648,i650,i652,i654,i656,i658,i660,
i662,i664,i666,i668,i670,i672,i674,i676,i678,i680,i682,i684,i686,i688,i690,
i692,i694,i696,i698,i700,i702,i704,i706,i708,i710,i712,i714,i716,i718,i720,
i722,i724,i726,i728,i730,i732,i734,i736,i738,i740,i742,i744,i746,i748,i750,
i752,i754,i756,i758,i760,i762,i764,i766,i768,i770,i772,i774,i776,i778,i780,
i782,i784,i786,i788,i790,i792,i794,i796,i798,i800,i802,i804,i806,i808,i810,
i812,i814,i816,i818,i820,i822,i824,i826,i828,i830,i832,i834,i836,i838,i840,
i842,i844,i846,i848,i850,i852,i854,i856,i858,i860,i862,i864,i866,i868,i870,
i872,i874,i876,i878,p0);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,i246,i248,i250,i252,i254,i256,i258,i260,i262,i264,i266,i268,i270,
i272,i274,i276,i278,i280,i282,i284,i286,i288,i290,i292,i294,i296,i298,i300,
i302,i304,i306,i308,i310,i312,i314,i316,i318,i320,i322,i324,i326,i328,i330,
i332,i334,i336,i338,i340,i342,i344,i346,i348,i350,i352,i354,i356,i358,i360,
i362,i364,i366,i368,i370,i372,i374,i376,i378,i380,i382,i384,i386,i388,i390,
i392,i394,i396,i398,i400,i402,i404,i406,i408,i410,i412,i414,i416,i418,i420,
i422,i424,i426,i428,i430,i432,i434,i436,i438,i440,i442,i444,i446,i448,i450,
i452,i454,i456,i458,i460,i462,i464,i466,i468,i470,i472,i474,i476,i478,i480,
i482,i484,i486,i488,i490,i492,i494,i496,i498,i500,i502,i504,i506,i508,i510,
i512,i514,i516,i518,i520,i522,i524,i526,i528,i530,i532,i534,i536,i538,i540,
i542,i544,i546,i548,i550,i552,i554,i556,i558,i560,i562,i564,i566,i568,i570,
i572,i574,i576,i578,i580,i582,i584,i586,i588,i590,i592,i594,i596,i598,i600,
i602,i604,i606,i608,i610,i612,i614,i616,i618,i620,i622,i624,i626,i628,i630,
i632,i634,i636,i638,i640,i642,i644,i646,i648,i650,i652,i654,i656,i658,i660,
i662,i664,i666,i668,i670,i672,i674,i676,i678,i680,i682,i684,i686,i688,i690,
i692,i694,i696,i698,i700,i702,i704,i706,i708,i710,i712,i714,i716,i718,i720,
i722,i724,i726,i728,i730,i732,i734,i736,i738,i740,i742,i744,i746,i748,i750,
i752,i754,i756,i758,i760,i762,i764,i766,i768,i770,i772,i774,i776,i778,i780,
i782,i784,i786,i788,i790,i792,i794,i796,i798,i800,i802,i804,i806,i808,i810,
i812,i814,i816,i818,i820,i822,i824,i826,i828,i830,i832,i834,i836,i838,i840,
i842,i844,i846,i848,i850,i852,i854,i856,i858,i860,i862,i864,i866,i868,i870,
i872,i874,i876,i878;

output p0;

wire na2504,na2780,a5360,a17682,c1,a5374,a16196,a18514,na18518,a18520,a18542,a18556,a18562,a19756,a19892,
na8812,a19894,a19900,a16186,a21664,a23736,a23742,z0,a8150,a24056,a24188,a24322,a24450,a24582,a24714,
a24846,a24974,a25106,a25236,na25240,a25242,na25818,na19408,a5352,z1,a25838,a25846,a25850,a25852,na26072,
na20174,na26078,na26106,na26594,na2536,na2752,na2516,na26612,a28188,a28194,a28236,a20078,a18850,a28448,a16250,
na28452,na25504,na25804,a25534,na28462,a25578,a28706,a18924,a28944,a19004,a29210,a19086,a29462,a19168,a29508,
na19250,a29548,na19332,na29552,a25628,na29562,na29572,a25672,na29582,na25716,na29592,na25760,na29602,a29642,na16278,
na29646,na29650,na29654,na29658,na29662,a16608,a29722,a20054,z2,a29728,a16712,a29788,a20028,a29794,a16816,
a29854,a20002,a29860,a16920,a29920,a19976,a29926,na17016,a29986,na19950,na29992,na17112,na30052,na19922,na30058,
na8954,na30072,a31018,a31020,a31040,na31048,a8946,na8986,na31060,na31072,na31086,na8924,na8870,a31088,na31092,
z3,na31152,na18526,a31160,na17784,z4,na31102,na31176,a31182,a8970,na31110,na31202,a31208,a9006,na31118,
na31222,na31228,na8906,a32370,a32380,na12366,na32396,a32386,na32402,na12312,na32408,na32414,na12250,na32420,na32426,
na12190,na32432,na32438,na16376,na17092,na18282,a16996,na18208,a16892,na18134,a16788,na18060,a16684,na17986,a16580,
na17912,a16514,na17844,na32454,a32470,a32486,na22814,na22822,na22834,na22842,na22854,na22862,na22878,na22886,na22898,
na22906,na21710,na21720,na21740,na21752,na21766,na21776,a21800,a21810,a21828,na21840,na21886,na21894,na21906,na21914,
na21926,na21934,a21950,a21958,a21970,na21978,na22020,na22028,na22040,na22048,na22060,na22068,a22084,a22092,a22104,
na22112,na22154,na22162,na22174,na22182,na22194,na22202,a22218,a22226,a22238,na22246,na22288,na22296,na22308,na22316,
na22328,na22336,a22352,a22360,a22372,na22380,na22422,na22430,na22442,na22450,na22462,na22470,a22486,a22494,a22506,
na22514,na22556,na22564,na22576,na22584,na22596,na22604,a22620,a22628,na22640,na22648,na26200,na26238,na26282,na26326,
na26370,na26414,a32504,a32508,a32538,a16440,na33374,na33380,na33402,na33408,a33430,na33436,a33458,na33464,a32966,
na33468,a32978,na33506,na33526,a31042,na24030,na33570,na33624,na33636,na33642,na33652,a34176,a32998,z5,na23774,
na24826,na34252,na34268,na34290,na34308,na34326,na25216,a34338,na24954,na34350,a34362,na24694,na24562,na24430,na24302,
na24168,na24036,na25086,a33014,a33032,a33046,a33066,a33078,a33094,a33106,na34374,na34380,na34386,na34392,na34398,
na34404,na34410,na34416,na34422,na34428,na34440,na34446,na34452,na34458,na34464,na34470,na34476,na34482,a34488,a34494,
na34506,na34512,na34518,na34524,na34530,na34536,na34542,na34548,a34554,a34560,na34572,na34578,na34584,na34590,na34596,
na34602,na34608,na34614,a34620,a34626,na34638,na34644,na34650,na34656,na34662,na34668,na34674,na34680,a34686,a34692,
na34704,na34710,na34716,na34722,na34728,na34734,na34740,na34746,a34752,a34758,na34770,na34776,na34782,na34788,na34794,
na34800,na34806,na34812,a34818,na34824,na34836,na34842,na34848,na34854,na34860,na34866,na34872,na34878,na34884,na34890,
a34894,z6,z7,z8,na17454,a34896,a34898,a34900,a34902,na17592,a34904,a34910,a21670,na34920,na34928,
na34936,na34946,na34954,na34962,na34970,na34976,a34988,a21880,na34994,a35000,na35006,na35012,na35018,na35024,na35030,
na35036,na35042,a35054,a22014,na35060,a35066,na35072,na35078,na35084,na35090,na35096,na35102,na35108,a35120,a22148,
na35126,a35132,na35138,na35144,na35150,na35156,na35162,na35168,na35174,a35186,a22282,na35192,a35198,na35204,na35210,
na35216,na35222,na35228,na35234,na35240,a35252,a22416,na35258,a35264,na35270,na35276,na35282,na35288,na35294,na35300,
na35306,na35318,a22550,na35324,a35330,na35336,na35342,na35348,na35354,na35360,na35366,na35372,na35386,a22808,na35392,
na35398,na35404,na35410,na35416,na35422,na35428,na35434,na35440,a35472,na8846,na8836,na8860,na8826,a35514,a35554,
a35588,a35636,a35664,a35700,a35720,a35748,na35754,na35760,na35766,na35772,na35778,na35784,na35790,na35796,na35802,
a32592,a32634,a32680,a32722,a32772,a32814,a32860,a32908,a33156,a33198,na35828,z9,z10,z11,z12,
na35836,na35856,na35862,na35880,na35886,na35896,na35902,na35912,na35922,na18744,a35930,z13,a35946,a35960,a35968,
na36056,na37126,na37160,na37184,na37206,na37222,na37246,na37266,na37386,na37400,na37448,na37476,na37482,a41638,a41644,
na41660,a41670,a41672,na41678,a41736,na41742,na41800,na41806,na41846,a44408,a44428,a41654,a44442,a44450,a44462,
a44472,a44482,a44490,a44498,a44506,a44514,a44520,a44526,a44532,a44538,a44544,a44550,a44556,a44562,a44568,
a44574,a44580,a44586,a44592,a44598,a44604,a44610,a44616,a44622,a44628,a44634,a44640,a44646,a44652,a44658,
a44664,a44670,a44676,a44682,a44688,a44694,a44700,a44706,a44712,a44718,a44724,a44730,a44736,a44742,a44748,
a44754,a44760,a44766,a44772,a44778,a44784,a44790,a44796,a44802,a44808,a44814,a44834,a45596,na8818,z14,
a8814,z15,z16,z17,na40992,na45602,a45608,a40642,z18,a45622,a46176,a48022,a48034,a48048,na48062,
a48584,a48590,a48596,a48602,a48608,a48614,a48620,a48626,a48632,a48638,a48644,a48650,a48656,a48662,a48668,
a48674,a48680,a48686,a48692,a48698,a48704,a48728,a48792,a48808,a49932,na49946,na49958,a49740,a49996,a49758,
a50024,a49784,a50066,a50084,a49802,a50114,a49824,a49842,a50136,a49862,a50164,a49880,a50176,z19,z20,
z21,z22,na50182,na50188,na50194,na50200,na50248,na50254,na50260,na50266,na50272,na50278,na50284,a50346,a50420,
na50426,a50620,a50646,a50672,a50698,a50724,a50750,a50776,a50802,a50828,a50854,na50954,na50958,na50962,na50970,
a50972,na18534,a50986,a50990,na50996,a51000,a5624,z23,z24,z25,z26,z27,a2502,a2504,a2506,
a2508,a2510,a2512,a2514,a2516,a2518,a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,
a2538,a2540,a2542,a2544,a2546,a2548,a2550,a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,
a2568,a2570,a2572,a2574,a2576,a2578,a2580,a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,
a2598,a2600,a2602,a2604,a2606,a2608,a2610,a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,
a2628,a2630,a2632,a2634,a2636,a2638,a2640,a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,
a2658,a2660,a2662,a2664,a2666,a2668,a2670,a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,
a2688,a2690,a2692,a2694,a2696,a2698,a2700,a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,
a2718,a2720,a2722,a2724,a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,
a2748,a2750,a2752,a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,
a2778,a2780,a2782,a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,
a2808,a2810,a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,
a2838,a2840,a2842,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,
a2868,a2870,a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,
a2898,a2900,a2902,a2904,a2906,a2908,a2910,a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,
a2928,a2930,a2932,a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,
a2958,a2960,a2962,a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,
a2988,a2990,a2992,a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,
a3018,a3020,a3022,a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,
a3048,a3050,a3052,a3054,a3056,a3058,a3060,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,
a3078,a3080,a3082,a3084,a3086,a3088,a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,
a3108,a3110,a3112,a3114,a3116,a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,
a3138,a3140,a3142,a3144,a3146,a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,
a3168,a3170,a3172,a3174,a3176,a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,
a3198,a3200,a3202,a3204,a3206,a3208,a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,
a3228,a3230,a3232,a3234,a3236,a3238,a3240,a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,
a3258,a3260,a3262,a3264,a3266,a3268,a3270,a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,
a3288,a3290,a3292,a3294,a3296,a3298,a3300,a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,
a3318,a3320,a3322,a3324,a3326,a3328,a3330,a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,
a3348,a3350,a3352,a3354,a3356,a3358,a3360,a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,
a3378,a3380,a3382,a3384,a3386,a3388,a3390,a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,
a3408,a3410,a3412,a3414,a3416,a3418,a3420,a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,
a3438,a3440,a3442,a3444,a3446,a3448,a3450,a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,
a3468,a3470,a3472,a3474,a3476,a3478,a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,
a3498,a3500,a3502,a3504,a3506,a3508,a3510,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,
a3528,a3530,a3532,a3534,a3536,a3538,a3540,a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,
a3558,a3560,a3562,a3564,a3566,a3568,a3570,a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,
a3588,a3590,a3592,a3594,a3596,a3598,a3600,a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,
a3618,a3620,a3622,a3624,a3626,a3628,a3630,a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,
a3648,a3650,a3652,a3654,a3656,a3658,a3660,a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,
a3678,a3680,a3682,a3684,a3686,a3688,a3690,a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,
a3708,a3710,a3712,a3714,a3716,a3718,a3720,a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,
a3738,a3740,a3742,a3744,a3746,a3748,a3750,a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,
a3768,a3770,a3772,a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,
a3798,a3800,a3802,a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,
a3828,a3830,a3832,a3834,a3836,a3838,a3840,a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,
a3858,a3860,a3862,a3864,a3866,a3868,a3870,a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,
a3888,a3890,a3892,a3894,a3896,a3898,a3900,a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,
a3918,a3920,a3922,a3924,a3926,a3928,a3930,a3932,a3934,a3936,a3938,a3940,a3942,a3944,a3946,
a3948,a3950,a3952,a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,
a3978,a3980,a3982,a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,
a4008,a4010,a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,
a4038,a4040,a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,
a4068,a4070,a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,a4096,
a4098,a4100,a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4124,a4126,
a4128,a4130,a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,a4152,a4154,a4156,
a4158,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,a4184,a4186,
a4188,a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,a4214,a4216,
a4218,a4220,a4222,a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,a4244,a4246,
a4248,a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,a4274,a4276,
a4278,a4280,a4282,a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,a4306,
a4308,a4310,a4312,a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4330,a4332,a4334,a4336,
a4338,a4340,a4342,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,
a4368,a4370,a4372,a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4390,a4392,a4394,a4396,
a4398,a4400,a4402,a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,
a4428,a4430,a4432,a4434,a4436,a4438,a4440,a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,
a4458,a4460,a4462,a4464,a4466,a4468,a4470,a4472,a4474,a4476,a4478,a4480,a4482,a4484,a4486,
a4488,a4490,a4492,a4494,a4496,a4498,a4500,a4502,a4504,a4506,a4508,a4510,a4512,a4514,a4516,
a4518,a4520,a4522,a4524,a4526,a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,
a4548,a4550,a4552,a4554,a4556,a4558,a4560,a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,
a4578,a4580,a4582,a4584,a4586,a4588,a4590,a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,
a4608,a4610,a4612,a4614,a4616,a4618,a4620,a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,
a4638,a4640,a4642,a4644,a4646,a4648,a4650,a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,
a4668,a4670,a4672,a4674,a4676,a4678,a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,a4696,
a4698,a4700,a4702,a4704,a4706,a4708,a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,a4726,
a4728,a4730,a4732,a4734,a4736,a4738,a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,a4756,
a4758,a4760,a4762,a4764,a4766,a4768,a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4784,a4786,
a4788,a4790,a4792,a4794,a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,
a4818,a4820,a4822,a4824,a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,a4844,a4846,
a4848,a4850,a4852,a4854,a4856,a4858,a4860,a4862,a4864,a4866,a4868,a4870,a4872,a4874,a4876,
a4878,a4880,a4882,a4884,a4886,a4888,a4890,a4892,a4894,a4896,a4898,a4900,a4902,a4904,a4906,
a4908,a4910,a4912,a4914,a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,
a4938,a4940,a4942,a4944,a4946,a4948,a4950,a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,
a4968,a4970,a4972,a4974,a4976,a4978,a4980,a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,
a4998,a5000,a5002,a5004,a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,
a5028,a5030,a5032,a5034,a5036,a5038,a5040,a5042,a5044,a5046,a5048,a5050,a5052,a5054,a5056,
a5058,a5060,a5062,a5064,a5066,a5068,a5070,a5072,a5074,a5076,a5078,a5080,a5082,a5084,a5086,
a5088,a5090,a5092,a5094,a5096,a5098,a5100,a5102,a5104,a5106,a5108,a5110,a5112,a5114,a5116,
a5118,a5120,a5122,a5124,a5126,a5128,a5130,a5132,a5134,a5136,a5138,a5140,a5142,a5144,a5146,
a5148,a5150,a5152,a5154,a5156,a5158,a5160,a5162,a5164,a5166,a5168,a5170,a5172,a5174,a5176,
a5178,a5180,a5182,a5184,a5186,a5188,a5190,a5192,a5194,a5196,a5198,a5200,a5202,a5204,a5206,
a5208,a5210,a5212,a5214,a5216,a5218,a5220,a5222,a5224,a5226,a5228,a5230,a5232,a5234,a5236,
a5238,a5240,a5242,a5244,a5246,a5248,a5250,a5252,a5254,a5256,a5258,a5260,a5262,a5264,a5266,
a5268,a5270,a5272,a5274,a5276,a5278,a5280,a5282,a5284,a5286,a5288,a5290,a5292,a5294,a5296,
a5298,a5300,a5302,a5304,a5306,a5308,a5310,a5312,a5314,a5316,a5318,a5320,a5322,a5324,a5326,
a5328,a5330,a5332,a5334,a5336,a5338,a5340,a5342,a5344,a5346,a5348,a5350,a5354,a5356,a5358,
a5362,a5364,a5366,a5368,a5370,a5372,a5376,a5378,a5380,a5382,a5384,a5386,a5388,a5390,a5392,
a5394,a5396,a5398,a5400,a5402,a5404,a5406,a5408,a5410,a5412,a5414,a5416,a5418,a5420,a5422,
a5424,a5426,a5428,a5430,a5432,a5434,a5436,a5438,a5440,a5442,a5444,a5446,a5448,a5450,a5452,
a5454,a5456,a5458,a5460,a5462,a5464,a5466,a5468,a5470,a5472,a5474,a5476,a5478,a5480,a5482,
a5484,a5486,a5488,a5490,a5492,a5494,a5496,a5498,a5500,a5502,a5504,a5506,a5508,a5510,a5512,
a5514,a5516,a5518,a5520,a5522,a5524,a5526,a5528,a5530,a5532,a5534,a5536,a5538,a5540,a5542,
a5544,a5546,a5548,a5550,a5552,a5554,a5556,a5558,a5560,a5562,a5564,a5566,a5568,a5570,a5572,
a5574,a5576,a5578,a5580,a5582,a5584,a5586,a5588,a5590,a5592,a5594,a5596,a5598,a5600,a5602,
a5604,a5606,a5608,a5610,a5612,a5614,a5616,a5618,a5620,a5622,a5626,a5628,a5630,a5632,a5634,
a5636,a5638,a5640,a5642,a5644,a5646,a5648,a5650,a5652,a5654,a5656,a5658,a5660,a5662,a5664,
a5666,a5668,a5670,a5672,a5674,a5676,a5678,a5680,a5682,a5684,a5686,a5688,a5690,a5692,a5694,
a5696,a5698,a5700,a5702,a5704,a5706,a5708,a5710,a5712,a5714,a5716,a5718,a5720,a5722,a5724,
a5726,a5728,a5730,a5732,a5734,a5736,a5738,a5740,a5742,a5744,a5746,a5748,a5750,a5752,a5754,
a5756,a5758,a5760,a5762,a5764,a5766,a5768,a5770,a5772,a5774,a5776,a5778,a5780,a5782,a5784,
a5786,a5788,a5790,a5792,a5794,a5796,a5798,a5800,a5802,a5804,a5806,a5808,a5810,a5812,a5814,
a5816,a5818,a5820,a5822,a5824,a5826,a5828,a5830,a5832,a5834,a5836,a5838,a5840,a5842,a5844,
a5846,a5848,a5850,a5852,a5854,a5856,a5858,a5860,a5862,a5864,a5866,a5868,a5870,a5872,a5874,
a5876,a5878,a5880,a5882,a5884,a5886,a5888,a5890,a5892,a5894,a5896,a5898,a5900,a5902,a5904,
a5906,a5908,a5910,a5912,a5914,a5916,a5918,a5920,a5922,a5924,a5926,a5928,a5930,a5932,a5934,
a5936,a5938,a5940,a5942,a5944,a5946,a5948,a5950,a5952,a5954,a5956,a5958,a5960,a5962,a5964,
a5966,a5968,a5970,a5972,a5974,a5976,a5978,a5980,a5982,a5984,a5986,a5988,a5990,a5992,a5994,
a5996,a5998,a6000,a6002,a6004,a6006,a6008,a6010,a6012,a6014,a6016,a6018,a6020,a6022,a6024,
a6026,a6028,a6030,a6032,a6034,a6036,a6038,a6040,a6042,a6044,a6046,a6048,a6050,a6052,a6054,
a6056,a6058,a6060,a6062,a6064,a6066,a6068,a6070,a6072,a6074,a6076,a6078,a6080,a6082,a6084,
a6086,a6088,a6090,a6092,a6094,a6096,a6098,a6100,a6102,a6104,a6106,a6108,a6110,a6112,a6114,
a6116,a6118,a6120,a6122,a6124,a6126,a6128,a6130,a6132,a6134,a6136,a6138,a6140,a6142,a6144,
a6146,a6148,a6150,a6152,a6154,a6156,a6158,a6160,a6162,a6164,a6166,a6168,a6170,a6172,a6174,
a6176,a6178,a6180,a6182,a6184,a6186,a6188,a6190,a6192,a6194,a6196,a6198,a6200,a6202,a6204,
a6206,a6208,a6210,a6212,a6214,a6216,a6218,a6220,a6222,a6224,a6226,a6228,a6230,a6232,a6234,
a6236,a6238,a6240,a6242,a6244,a6246,a6248,a6250,a6252,a6254,a6256,a6258,a6260,a6262,a6264,
a6266,a6268,a6270,a6272,a6274,a6276,a6278,a6280,a6282,a6284,a6286,a6288,a6290,a6292,a6294,
a6296,a6298,a6300,a6302,a6304,a6306,a6308,a6310,a6312,a6314,a6316,a6318,a6320,a6322,a6324,
a6326,a6328,a6330,a6332,a6334,a6336,a6338,a6340,a6342,a6344,a6346,a6348,a6350,a6352,a6354,
a6356,a6358,a6360,a6362,a6364,a6366,a6368,a6370,a6372,a6374,a6376,a6378,a6380,a6382,a6384,
a6386,a6388,a6390,a6392,a6394,a6396,a6398,a6400,a6402,a6404,a6406,a6408,a6410,a6412,a6414,
a6416,a6418,a6420,a6422,a6424,a6426,a6428,a6430,a6432,a6434,a6436,a6438,a6440,a6442,a6444,
a6446,a6448,a6450,a6452,a6454,a6456,a6458,a6460,a6462,a6464,a6466,a6468,a6470,a6472,a6474,
a6476,a6478,a6480,a6482,a6484,a6486,a6488,a6490,a6492,a6494,a6496,a6498,a6500,a6502,a6504,
a6506,a6508,a6510,a6512,a6514,a6516,a6518,a6520,a6522,a6524,a6526,a6528,a6530,a6532,a6534,
a6536,a6538,a6540,a6542,a6544,a6546,a6548,a6550,a6552,a6554,a6556,a6558,a6560,a6562,a6564,
a6566,a6568,a6570,a6572,a6574,a6576,a6578,a6580,a6582,a6584,a6586,a6588,a6590,a6592,a6594,
a6596,a6598,a6600,a6602,a6604,a6606,a6608,a6610,a6612,a6614,a6616,a6618,a6620,a6622,a6624,
a6626,a6628,a6630,a6632,a6634,a6636,a6638,a6640,a6642,a6644,a6646,a6648,a6650,a6652,a6654,
a6656,a6658,a6660,a6662,a6664,a6666,a6668,a6670,a6672,a6674,a6676,a6678,a6680,a6682,a6684,
a6686,a6688,a6690,a6692,a6694,a6696,a6698,a6700,a6702,a6704,a6706,a6708,a6710,a6712,a6714,
a6716,a6718,a6720,a6722,a6724,a6726,a6728,a6730,a6732,a6734,a6736,a6738,a6740,a6742,a6744,
a6746,a6748,a6750,a6752,a6754,a6756,a6758,a6760,a6762,a6764,a6766,a6768,a6770,a6772,a6774,
a6776,a6778,a6780,a6782,a6784,a6786,a6788,a6790,a6792,a6794,a6796,a6798,a6800,a6802,a6804,
a6806,a6808,a6810,a6812,a6814,a6816,a6818,a6820,a6822,a6824,a6826,a6828,a6830,a6832,a6834,
a6836,a6838,a6840,a6842,a6844,a6846,a6848,a6850,a6852,a6854,a6856,a6858,a6860,a6862,a6864,
a6866,a6868,a6870,a6872,a6874,a6876,a6878,a6880,a6882,a6884,a6886,a6888,a6890,a6892,a6894,
a6896,a6898,a6900,a6902,a6904,a6906,a6908,a6910,a6912,a6914,a6916,a6918,a6920,a6922,a6924,
a6926,a6928,a6930,a6932,a6934,a6936,a6938,a6940,a6942,a6944,a6946,a6948,a6950,a6952,a6954,
a6956,a6958,a6960,a6962,a6964,a6966,a6968,a6970,a6972,a6974,a6976,a6978,a6980,a6982,a6984,
a6986,a6988,a6990,a6992,a6994,a6996,a6998,a7000,a7002,a7004,a7006,a7008,a7010,a7012,a7014,
a7016,a7018,a7020,a7022,a7024,a7026,a7028,a7030,a7032,a7034,a7036,a7038,a7040,a7042,a7044,
a7046,a7048,a7050,a7052,a7054,a7056,a7058,a7060,a7062,a7064,a7066,a7068,a7070,a7072,a7074,
a7076,a7078,a7080,a7082,a7084,a7086,a7088,a7090,a7092,a7094,a7096,a7098,a7100,a7102,a7104,
a7106,a7108,a7110,a7112,a7114,a7116,a7118,a7120,a7122,a7124,a7126,a7128,a7130,a7132,a7134,
a7136,a7138,a7140,a7142,a7144,a7146,a7148,a7150,a7152,a7154,a7156,a7158,a7160,a7162,a7164,
a7166,a7168,a7170,a7172,a7174,a7176,a7178,a7180,a7182,a7184,a7186,a7188,a7190,a7192,a7194,
a7196,a7198,a7200,a7202,a7204,a7206,a7208,a7210,a7212,a7214,a7216,a7218,a7220,a7222,a7224,
a7226,a7228,a7230,a7232,a7234,a7236,a7238,a7240,a7242,a7244,a7246,a7248,a7250,a7252,a7254,
a7256,a7258,a7260,a7262,a7264,a7266,a7268,a7270,a7272,a7274,a7276,a7278,a7280,a7282,a7284,
a7286,a7288,a7290,a7292,a7294,a7296,a7298,a7300,a7302,a7304,a7306,a7308,a7310,a7312,a7314,
a7316,a7318,a7320,a7322,a7324,a7326,a7328,a7330,a7332,a7334,a7336,a7338,a7340,a7342,a7344,
a7346,a7348,a7350,a7352,a7354,a7356,a7358,a7360,a7362,a7364,a7366,a7368,a7370,a7372,a7374,
a7376,a7378,a7380,a7382,a7384,a7386,a7388,a7390,a7392,a7394,a7396,a7398,a7400,a7402,a7404,
a7406,a7408,a7410,a7412,a7414,a7416,a7418,a7420,a7422,a7424,a7426,a7428,a7430,a7432,a7434,
a7436,a7438,a7440,a7442,a7444,a7446,a7448,a7450,a7452,a7454,a7456,a7458,a7460,a7462,a7464,
a7466,a7468,a7470,a7472,a7474,a7476,a7478,a7480,a7482,a7484,a7486,a7488,a7490,a7492,a7494,
a7496,a7498,a7500,a7502,a7504,a7506,a7508,a7510,a7512,a7514,a7516,a7518,a7520,a7522,a7524,
a7526,a7528,a7530,a7532,a7534,a7536,a7538,a7540,a7542,a7544,a7546,a7548,a7550,a7552,a7554,
a7556,a7558,a7560,a7562,a7564,a7566,a7568,a7570,a7572,a7574,a7576,a7578,a7580,a7582,a7584,
a7586,a7588,a7590,a7592,a7594,a7596,a7598,a7600,a7602,a7604,a7606,a7608,a7610,a7612,a7614,
a7616,a7618,a7620,a7622,a7624,a7626,a7628,a7630,a7632,a7634,a7636,a7638,a7640,a7642,a7644,
a7646,a7648,a7650,a7652,a7654,a7656,a7658,a7660,a7662,a7664,a7666,a7668,a7670,a7672,a7674,
a7676,a7678,a7680,a7682,a7684,a7686,a7688,a7690,a7692,a7694,a7696,a7698,a7700,a7702,a7704,
a7706,a7708,a7710,a7712,a7714,a7716,a7718,a7720,a7722,a7724,a7726,a7728,a7730,a7732,a7734,
a7736,a7738,a7740,a7742,a7744,a7746,a7748,a7750,a7752,a7754,a7756,a7758,a7760,a7762,a7764,
a7766,a7768,a7770,a7772,a7774,a7776,a7778,a7780,a7782,a7784,a7786,a7788,a7790,a7792,a7794,
a7796,a7798,a7800,a7802,a7804,a7806,a7808,a7810,a7812,a7814,a7816,a7818,a7820,a7822,a7824,
a7826,a7828,a7830,a7832,a7834,a7836,a7838,a7840,a7842,a7844,a7846,a7848,a7850,a7852,a7854,
a7856,a7858,a7860,a7862,a7864,a7866,a7868,a7870,a7872,a7874,a7876,a7878,a7880,a7882,a7884,
a7886,a7888,a7890,a7892,a7894,a7896,a7898,a7900,a7902,a7904,a7906,a7908,a7910,a7912,a7914,
a7916,a7918,a7920,a7922,a7924,a7926,a7928,a7930,a7932,a7934,a7936,a7938,a7940,a7942,a7944,
a7946,a7948,a7950,a7952,a7954,a7956,a7958,a7960,a7962,a7964,a7966,a7968,a7970,a7972,a7974,
a7976,a7978,a7980,a7982,a7984,a7986,a7988,a7990,a7992,a7994,a7996,a7998,a8000,a8002,a8004,
a8006,a8008,a8010,a8012,a8014,a8016,a8018,a8020,a8022,a8024,a8026,a8028,a8030,a8032,a8034,
a8036,a8038,a8040,a8042,a8044,a8046,a8048,a8050,a8052,a8054,a8056,a8058,a8060,a8062,a8064,
a8066,a8068,a8070,a8072,a8074,a8076,a8078,a8080,a8082,a8084,a8086,a8088,a8090,a8092,a8094,
a8096,a8098,a8100,a8102,a8104,a8106,a8108,a8110,a8112,a8114,a8116,a8118,a8120,a8122,a8124,
a8126,a8128,a8130,a8132,a8134,a8136,a8138,a8140,a8142,a8144,a8146,a8148,a8152,a8154,a8156,
a8158,a8160,a8162,a8164,a8166,a8168,a8170,a8172,a8174,a8176,a8178,a8180,a8182,a8184,a8186,
a8188,a8190,a8192,a8194,a8196,a8198,a8200,a8202,a8204,a8206,a8208,a8210,a8212,a8214,a8216,
a8218,a8220,a8222,a8224,a8226,a8228,a8230,a8232,a8234,a8236,a8238,a8240,a8242,a8244,a8246,
a8248,a8250,a8252,a8254,a8256,a8258,a8260,a8262,a8264,a8266,a8268,a8270,a8272,a8274,a8276,
a8278,a8280,a8282,a8284,a8286,a8288,a8290,a8292,a8294,a8296,a8298,a8300,a8302,a8304,a8306,
a8308,a8310,a8312,a8314,a8316,a8318,a8320,a8322,a8324,a8326,a8328,a8330,a8332,a8334,a8336,
a8338,a8340,a8342,a8344,a8346,a8348,a8350,a8352,a8354,a8356,a8358,a8360,a8362,a8364,a8366,
a8368,a8370,a8372,a8374,a8376,a8378,a8380,a8382,a8384,a8386,a8388,a8390,a8392,a8394,a8396,
a8398,a8400,a8402,a8404,a8406,a8408,a8410,a8412,a8414,a8416,a8418,a8420,a8422,a8424,a8426,
a8428,a8430,a8432,a8434,a8436,a8438,a8440,a8442,a8444,a8446,a8448,a8450,a8452,a8454,a8456,
a8458,a8460,a8462,a8464,a8466,a8468,a8470,a8472,a8474,a8476,a8478,a8480,a8482,a8484,a8486,
a8488,a8490,a8492,a8494,a8496,a8498,a8500,a8502,a8504,a8506,a8508,a8510,a8512,a8514,a8516,
a8518,a8520,a8522,a8524,a8526,a8528,a8530,a8532,a8534,a8536,a8538,a8540,a8542,a8544,a8546,
a8548,a8550,a8552,a8554,a8556,a8558,a8560,a8562,a8564,a8566,a8568,a8570,a8572,a8574,a8576,
a8578,a8580,a8582,a8584,a8586,a8588,a8590,a8592,a8594,a8596,a8598,a8600,a8602,a8604,a8606,
a8608,a8610,a8612,a8614,a8616,a8618,a8620,a8622,a8624,a8626,a8628,a8630,a8632,a8634,a8636,
a8638,a8640,a8642,a8644,a8646,a8648,a8650,a8652,a8654,a8656,a8658,a8660,a8662,a8664,a8666,
a8668,a8670,a8672,a8674,a8676,a8678,a8680,a8682,a8684,a8686,a8688,a8690,a8692,a8694,a8696,
a8698,a8700,a8702,a8704,a8706,a8708,a8710,a8712,a8714,a8716,a8718,a8720,a8722,a8724,a8726,
a8728,a8730,a8732,a8734,a8736,a8738,a8740,a8742,a8744,a8746,a8748,a8750,a8752,a8754,a8756,
a8758,a8760,a8762,a8764,a8766,a8768,a8770,a8772,a8774,a8776,a8778,a8780,a8782,a8784,a8786,
a8788,a8790,a8792,a8794,a8796,a8798,a8800,a8802,a8804,a8806,a8808,a8810,a8812,a8816,a8818,
a8820,a8822,a8824,a8826,a8828,a8830,a8832,a8834,a8836,a8838,a8840,a8842,a8844,a8846,a8848,
a8850,a8852,a8854,a8856,a8858,a8860,a8862,a8864,a8866,a8868,a8870,a8872,a8874,a8876,a8878,
a8880,a8882,a8884,a8886,a8888,a8890,a8892,a8894,a8896,a8898,a8900,a8902,a8904,a8906,a8908,
a8910,a8912,a8914,a8916,a8918,a8920,a8922,a8924,a8926,a8928,a8930,a8932,a8934,a8936,a8938,
a8940,a8942,a8944,a8948,a8950,a8952,a8954,a8956,a8958,a8960,a8962,a8964,a8966,a8968,a8972,
a8974,a8976,a8978,a8980,a8982,a8984,a8986,a8988,a8990,a8992,a8994,a8996,a8998,a9000,a9002,
a9004,a9008,a9010,a9012,a9014,a9016,a9018,a9020,a9022,a9024,a9026,a9028,a9030,a9032,a9034,
a9036,a9038,a9040,a9042,a9044,a9046,a9048,a9050,a9052,a9054,a9056,a9058,a9060,a9062,a9064,
a9066,a9068,a9070,a9072,a9074,a9076,a9078,a9080,a9082,a9084,a9086,a9088,a9090,a9092,a9094,
a9096,a9098,a9100,a9102,a9104,a9106,a9108,a9110,a9112,a9114,a9116,a9118,a9120,a9122,a9124,
a9126,a9128,a9130,a9132,a9134,a9136,a9138,a9140,a9142,a9144,a9146,a9148,a9150,a9152,a9154,
a9156,a9158,a9160,a9162,a9164,a9166,a9168,a9170,a9172,a9174,a9176,a9178,a9180,a9182,a9184,
a9186,a9188,a9190,a9192,a9194,a9196,a9198,a9200,a9202,a9204,a9206,a9208,a9210,a9212,a9214,
a9216,a9218,a9220,a9222,a9224,a9226,a9228,a9230,a9232,a9234,a9236,a9238,a9240,a9242,a9244,
a9246,a9248,a9250,a9252,a9254,a9256,a9258,a9260,a9262,a9264,a9266,a9268,a9270,a9272,a9274,
a9276,a9278,a9280,a9282,a9284,a9286,a9288,a9290,a9292,a9294,a9296,a9298,a9300,a9302,a9304,
a9306,a9308,a9310,a9312,a9314,a9316,a9318,a9320,a9322,a9324,a9326,a9328,a9330,a9332,a9334,
a9336,a9338,a9340,a9342,a9344,a9346,a9348,a9350,a9352,a9354,a9356,a9358,a9360,a9362,a9364,
a9366,a9368,a9370,a9372,a9374,a9376,a9378,a9380,a9382,a9384,a9386,a9388,a9390,a9392,a9394,
a9396,a9398,a9400,a9402,a9404,a9406,a9408,a9410,a9412,a9414,a9416,a9418,a9420,a9422,a9424,
a9426,a9428,a9430,a9432,a9434,a9436,a9438,a9440,a9442,a9444,a9446,a9448,a9450,a9452,a9454,
a9456,a9458,a9460,a9462,a9464,a9466,a9468,a9470,a9472,a9474,a9476,a9478,a9480,a9482,a9484,
a9486,a9488,a9490,a9492,a9494,a9496,a9498,a9500,a9502,a9504,a9506,a9508,a9510,a9512,a9514,
a9516,a9518,a9520,a9522,a9524,a9526,a9528,a9530,a9532,a9534,a9536,a9538,a9540,a9542,a9544,
a9546,a9548,a9550,a9552,a9554,a9556,a9558,a9560,a9562,a9564,a9566,a9568,a9570,a9572,a9574,
a9576,a9578,a9580,a9582,a9584,a9586,a9588,a9590,a9592,a9594,a9596,a9598,a9600,a9602,a9604,
a9606,a9608,a9610,a9612,a9614,a9616,a9618,a9620,a9622,a9624,a9626,a9628,a9630,a9632,a9634,
a9636,a9638,a9640,a9642,a9644,a9646,a9648,a9650,a9652,a9654,a9656,a9658,a9660,a9662,a9664,
a9666,a9668,a9670,a9672,a9674,a9676,a9678,a9680,a9682,a9684,a9686,a9688,a9690,a9692,a9694,
a9696,a9698,a9700,a9702,a9704,a9706,a9708,a9710,a9712,a9714,a9716,a9718,a9720,a9722,a9724,
a9726,a9728,a9730,a9732,a9734,a9736,a9738,a9740,a9742,a9744,a9746,a9748,a9750,a9752,a9754,
a9756,a9758,a9760,a9762,a9764,a9766,a9768,a9770,a9772,a9774,a9776,a9778,a9780,a9782,a9784,
a9786,a9788,a9790,a9792,a9794,a9796,a9798,a9800,a9802,a9804,a9806,a9808,a9810,a9812,a9814,
a9816,a9818,a9820,a9822,a9824,a9826,a9828,a9830,a9832,a9834,a9836,a9838,a9840,a9842,a9844,
a9846,a9848,a9850,a9852,a9854,a9856,a9858,a9860,a9862,a9864,a9866,a9868,a9870,a9872,a9874,
a9876,a9878,a9880,a9882,a9884,a9886,a9888,a9890,a9892,a9894,a9896,a9898,a9900,a9902,a9904,
a9906,a9908,a9910,a9912,a9914,a9916,a9918,a9920,a9922,a9924,a9926,a9928,a9930,a9932,a9934,
a9936,a9938,a9940,a9942,a9944,a9946,a9948,a9950,a9952,a9954,a9956,a9958,a9960,a9962,a9964,
a9966,a9968,a9970,a9972,a9974,a9976,a9978,a9980,a9982,a9984,a9986,a9988,a9990,a9992,a9994,
a9996,a9998,a10000,a10002,a10004,a10006,a10008,a10010,a10012,a10014,a10016,a10018,a10020,a10022,a10024,
a10026,a10028,a10030,a10032,a10034,a10036,a10038,a10040,a10042,a10044,a10046,a10048,a10050,a10052,a10054,
a10056,a10058,a10060,a10062,a10064,a10066,a10068,a10070,a10072,a10074,a10076,a10078,a10080,a10082,a10084,
a10086,a10088,a10090,a10092,a10094,a10096,a10098,a10100,a10102,a10104,a10106,a10108,a10110,a10112,a10114,
a10116,a10118,a10120,a10122,a10124,a10126,a10128,a10130,a10132,a10134,a10136,a10138,a10140,a10142,a10144,
a10146,a10148,a10150,a10152,a10154,a10156,a10158,a10160,a10162,a10164,a10166,a10168,a10170,a10172,a10174,
a10176,a10178,a10180,a10182,a10184,a10186,a10188,a10190,a10192,a10194,a10196,a10198,a10200,a10202,a10204,
a10206,a10208,a10210,a10212,a10214,a10216,a10218,a10220,a10222,a10224,a10226,a10228,a10230,a10232,a10234,
a10236,a10238,a10240,a10242,a10244,a10246,a10248,a10250,a10252,a10254,a10256,a10258,a10260,a10262,a10264,
a10266,a10268,a10270,a10272,a10274,a10276,a10278,a10280,a10282,a10284,a10286,a10288,a10290,a10292,a10294,
a10296,a10298,a10300,a10302,a10304,a10306,a10308,a10310,a10312,a10314,a10316,a10318,a10320,a10322,a10324,
a10326,a10328,a10330,a10332,a10334,a10336,a10338,a10340,a10342,a10344,a10346,a10348,a10350,a10352,a10354,
a10356,a10358,a10360,a10362,a10364,a10366,a10368,a10370,a10372,a10374,a10376,a10378,a10380,a10382,a10384,
a10386,a10388,a10390,a10392,a10394,a10396,a10398,a10400,a10402,a10404,a10406,a10408,a10410,a10412,a10414,
a10416,a10418,a10420,a10422,a10424,a10426,a10428,a10430,a10432,a10434,a10436,a10438,a10440,a10442,a10444,
a10446,a10448,a10450,a10452,a10454,a10456,a10458,a10460,a10462,a10464,a10466,a10468,a10470,a10472,a10474,
a10476,a10478,a10480,a10482,a10484,a10486,a10488,a10490,a10492,a10494,a10496,a10498,a10500,a10502,a10504,
a10506,a10508,a10510,a10512,a10514,a10516,a10518,a10520,a10522,a10524,a10526,a10528,a10530,a10532,a10534,
a10536,a10538,a10540,a10542,a10544,a10546,a10548,a10550,a10552,a10554,a10556,a10558,a10560,a10562,a10564,
a10566,a10568,a10570,a10572,a10574,a10576,a10578,a10580,a10582,a10584,a10586,a10588,a10590,a10592,a10594,
a10596,a10598,a10600,a10602,a10604,a10606,a10608,a10610,a10612,a10614,a10616,a10618,a10620,a10622,a10624,
a10626,a10628,a10630,a10632,a10634,a10636,a10638,a10640,a10642,a10644,a10646,a10648,a10650,a10652,a10654,
a10656,a10658,a10660,a10662,a10664,a10666,a10668,a10670,a10672,a10674,a10676,a10678,a10680,a10682,a10684,
a10686,a10688,a10690,a10692,a10694,a10696,a10698,a10700,a10702,a10704,a10706,a10708,a10710,a10712,a10714,
a10716,a10718,a10720,a10722,a10724,a10726,a10728,a10730,a10732,a10734,a10736,a10738,a10740,a10742,a10744,
a10746,a10748,a10750,a10752,a10754,a10756,a10758,a10760,a10762,a10764,a10766,a10768,a10770,a10772,a10774,
a10776,a10778,a10780,a10782,a10784,a10786,a10788,a10790,a10792,a10794,a10796,a10798,a10800,a10802,a10804,
a10806,a10808,a10810,a10812,a10814,a10816,a10818,a10820,a10822,a10824,a10826,a10828,a10830,a10832,a10834,
a10836,a10838,a10840,a10842,a10844,a10846,a10848,a10850,a10852,a10854,a10856,a10858,a10860,a10862,a10864,
a10866,a10868,a10870,a10872,a10874,a10876,a10878,a10880,a10882,a10884,a10886,a10888,a10890,a10892,a10894,
a10896,a10898,a10900,a10902,a10904,a10906,a10908,a10910,a10912,a10914,a10916,a10918,a10920,a10922,a10924,
a10926,a10928,a10930,a10932,a10934,a10936,a10938,a10940,a10942,a10944,a10946,a10948,a10950,a10952,a10954,
a10956,a10958,a10960,a10962,a10964,a10966,a10968,a10970,a10972,a10974,a10976,a10978,a10980,a10982,a10984,
a10986,a10988,a10990,a10992,a10994,a10996,a10998,a11000,a11002,a11004,a11006,a11008,a11010,a11012,a11014,
a11016,a11018,a11020,a11022,a11024,a11026,a11028,a11030,a11032,a11034,a11036,a11038,a11040,a11042,a11044,
a11046,a11048,a11050,a11052,a11054,a11056,a11058,a11060,a11062,a11064,a11066,a11068,a11070,a11072,a11074,
a11076,a11078,a11080,a11082,a11084,a11086,a11088,a11090,a11092,a11094,a11096,a11098,a11100,a11102,a11104,
a11106,a11108,a11110,a11112,a11114,a11116,a11118,a11120,a11122,a11124,a11126,a11128,a11130,a11132,a11134,
a11136,a11138,a11140,a11142,a11144,a11146,a11148,a11150,a11152,a11154,a11156,a11158,a11160,a11162,a11164,
a11166,a11168,a11170,a11172,a11174,a11176,a11178,a11180,a11182,a11184,a11186,a11188,a11190,a11192,a11194,
a11196,a11198,a11200,a11202,a11204,a11206,a11208,a11210,a11212,a11214,a11216,a11218,a11220,a11222,a11224,
a11226,a11228,a11230,a11232,a11234,a11236,a11238,a11240,a11242,a11244,a11246,a11248,a11250,a11252,a11254,
a11256,a11258,a11260,a11262,a11264,a11266,a11268,a11270,a11272,a11274,a11276,a11278,a11280,a11282,a11284,
a11286,a11288,a11290,a11292,a11294,a11296,a11298,a11300,a11302,a11304,a11306,a11308,a11310,a11312,a11314,
a11316,a11318,a11320,a11322,a11324,a11326,a11328,a11330,a11332,a11334,a11336,a11338,a11340,a11342,a11344,
a11346,a11348,a11350,a11352,a11354,a11356,a11358,a11360,a11362,a11364,a11366,a11368,a11370,a11372,a11374,
a11376,a11378,a11380,a11382,a11384,a11386,a11388,a11390,a11392,a11394,a11396,a11398,a11400,a11402,a11404,
a11406,a11408,a11410,a11412,a11414,a11416,a11418,a11420,a11422,a11424,a11426,a11428,a11430,a11432,a11434,
a11436,a11438,a11440,a11442,a11444,a11446,a11448,a11450,a11452,a11454,a11456,a11458,a11460,a11462,a11464,
a11466,a11468,a11470,a11472,a11474,a11476,a11478,a11480,a11482,a11484,a11486,a11488,a11490,a11492,a11494,
a11496,a11498,a11500,a11502,a11504,a11506,a11508,a11510,a11512,a11514,a11516,a11518,a11520,a11522,a11524,
a11526,a11528,a11530,a11532,a11534,a11536,a11538,a11540,a11542,a11544,a11546,a11548,a11550,a11552,a11554,
a11556,a11558,a11560,a11562,a11564,a11566,a11568,a11570,a11572,a11574,a11576,a11578,a11580,a11582,a11584,
a11586,a11588,a11590,a11592,a11594,a11596,a11598,a11600,a11602,a11604,a11606,a11608,a11610,a11612,a11614,
a11616,a11618,a11620,a11622,a11624,a11626,a11628,a11630,a11632,a11634,a11636,a11638,a11640,a11642,a11644,
a11646,a11648,a11650,a11652,a11654,a11656,a11658,a11660,a11662,a11664,a11666,a11668,a11670,a11672,a11674,
a11676,a11678,a11680,a11682,a11684,a11686,a11688,a11690,a11692,a11694,a11696,a11698,a11700,a11702,a11704,
a11706,a11708,a11710,a11712,a11714,a11716,a11718,a11720,a11722,a11724,a11726,a11728,a11730,a11732,a11734,
a11736,a11738,a11740,a11742,a11744,a11746,a11748,a11750,a11752,a11754,a11756,a11758,a11760,a11762,a11764,
a11766,a11768,a11770,a11772,a11774,a11776,a11778,a11780,a11782,a11784,a11786,a11788,a11790,a11792,a11794,
a11796,a11798,a11800,a11802,a11804,a11806,a11808,a11810,a11812,a11814,a11816,a11818,a11820,a11822,a11824,
a11826,a11828,a11830,a11832,a11834,a11836,a11838,a11840,a11842,a11844,a11846,a11848,a11850,a11852,a11854,
a11856,a11858,a11860,a11862,a11864,a11866,a11868,a11870,a11872,a11874,a11876,a11878,a11880,a11882,a11884,
a11886,a11888,a11890,a11892,a11894,a11896,a11898,a11900,a11902,a11904,a11906,a11908,a11910,a11912,a11914,
a11916,a11918,a11920,a11922,a11924,a11926,a11928,a11930,a11932,a11934,a11936,a11938,a11940,a11942,a11944,
a11946,a11948,a11950,a11952,a11954,a11956,a11958,a11960,a11962,a11964,a11966,a11968,a11970,a11972,a11974,
a11976,a11978,a11980,a11982,a11984,a11986,a11988,a11990,a11992,a11994,a11996,a11998,a12000,a12002,a12004,
a12006,a12008,a12010,a12012,a12014,a12016,a12018,a12020,a12022,a12024,a12026,a12028,a12030,a12032,a12034,
a12036,a12038,a12040,a12042,a12044,a12046,a12048,a12050,a12052,a12054,a12056,a12058,a12060,a12062,a12064,
a12066,a12068,a12070,a12072,a12074,a12076,a12078,a12080,a12082,a12084,a12086,a12088,a12090,a12092,a12094,
a12096,a12098,a12100,a12102,a12104,a12106,a12108,a12110,a12112,a12114,a12116,a12118,a12120,a12122,a12124,
a12126,a12128,a12130,a12132,a12134,a12136,a12138,a12140,a12142,a12144,a12146,a12148,a12150,a12152,a12154,
a12156,a12158,a12160,a12162,a12164,a12166,a12168,a12170,a12172,a12174,a12176,a12178,a12180,a12182,a12184,
a12186,a12188,a12190,a12192,a12194,a12196,a12198,a12200,a12202,a12204,a12206,a12208,a12210,a12212,a12214,
a12216,a12218,a12220,a12222,a12224,a12226,a12228,a12230,a12232,a12234,a12236,a12238,a12240,a12242,a12244,
a12246,a12248,a12250,a12252,a12254,a12256,a12258,a12260,a12262,a12264,a12266,a12268,a12270,a12272,a12274,
a12276,a12278,a12280,a12282,a12284,a12286,a12288,a12290,a12292,a12294,a12296,a12298,a12300,a12302,a12304,
a12306,a12308,a12310,a12312,a12314,a12316,a12318,a12320,a12322,a12324,a12326,a12328,a12330,a12332,a12334,
a12336,a12338,a12340,a12342,a12344,a12346,a12348,a12350,a12352,a12354,a12356,a12358,a12360,a12362,a12364,
a12366,a12368,a12370,a12372,a12374,a12376,a12378,a12380,a12382,a12384,a12386,a12388,a12390,a12392,a12394,
a12396,a12398,a12400,a12402,a12404,a12406,a12408,a12410,a12412,a12414,a12416,a12418,a12420,a12422,a12424,
a12426,a12428,a12430,a12432,a12434,a12436,a12438,a12440,a12442,a12444,a12446,a12448,a12450,a12452,a12454,
a12456,a12458,a12460,a12462,a12464,a12466,a12468,a12470,a12472,a12474,a12476,a12478,a12480,a12482,a12484,
a12486,a12488,a12490,a12492,a12494,a12496,a12498,a12500,a12502,a12504,a12506,a12508,a12510,a12512,a12514,
a12516,a12518,a12520,a12522,a12524,a12526,a12528,a12530,a12532,a12534,a12536,a12538,a12540,a12542,a12544,
a12546,a12548,a12550,a12552,a12554,a12556,a12558,a12560,a12562,a12564,a12566,a12568,a12570,a12572,a12574,
a12576,a12578,a12580,a12582,a12584,a12586,a12588,a12590,a12592,a12594,a12596,a12598,a12600,a12602,a12604,
a12606,a12608,a12610,a12612,a12614,a12616,a12618,a12620,a12622,a12624,a12626,a12628,a12630,a12632,a12634,
a12636,a12638,a12640,a12642,a12644,a12646,a12648,a12650,a12652,a12654,a12656,a12658,a12660,a12662,a12664,
a12666,a12668,a12670,a12672,a12674,a12676,a12678,a12680,a12682,a12684,a12686,a12688,a12690,a12692,a12694,
a12696,a12698,a12700,a12702,a12704,a12706,a12708,a12710,a12712,a12714,a12716,a12718,a12720,a12722,a12724,
a12726,a12728,a12730,a12732,a12734,a12736,a12738,a12740,a12742,a12744,a12746,a12748,a12750,a12752,a12754,
a12756,a12758,a12760,a12762,a12764,a12766,a12768,a12770,a12772,a12774,a12776,a12778,a12780,a12782,a12784,
a12786,a12788,a12790,a12792,a12794,a12796,a12798,a12800,a12802,a12804,a12806,a12808,a12810,a12812,a12814,
a12816,a12818,a12820,a12822,a12824,a12826,a12828,a12830,a12832,a12834,a12836,a12838,a12840,a12842,a12844,
a12846,a12848,a12850,a12852,a12854,a12856,a12858,a12860,a12862,a12864,a12866,a12868,a12870,a12872,a12874,
a12876,a12878,a12880,a12882,a12884,a12886,a12888,a12890,a12892,a12894,a12896,a12898,a12900,a12902,a12904,
a12906,a12908,a12910,a12912,a12914,a12916,a12918,a12920,a12922,a12924,a12926,a12928,a12930,a12932,a12934,
a12936,a12938,a12940,a12942,a12944,a12946,a12948,a12950,a12952,a12954,a12956,a12958,a12960,a12962,a12964,
a12966,a12968,a12970,a12972,a12974,a12976,a12978,a12980,a12982,a12984,a12986,a12988,a12990,a12992,a12994,
a12996,a12998,a13000,a13002,a13004,a13006,a13008,a13010,a13012,a13014,a13016,a13018,a13020,a13022,a13024,
a13026,a13028,a13030,a13032,a13034,a13036,a13038,a13040,a13042,a13044,a13046,a13048,a13050,a13052,a13054,
a13056,a13058,a13060,a13062,a13064,a13066,a13068,a13070,a13072,a13074,a13076,a13078,a13080,a13082,a13084,
a13086,a13088,a13090,a13092,a13094,a13096,a13098,a13100,a13102,a13104,a13106,a13108,a13110,a13112,a13114,
a13116,a13118,a13120,a13122,a13124,a13126,a13128,a13130,a13132,a13134,a13136,a13138,a13140,a13142,a13144,
a13146,a13148,a13150,a13152,a13154,a13156,a13158,a13160,a13162,a13164,a13166,a13168,a13170,a13172,a13174,
a13176,a13178,a13180,a13182,a13184,a13186,a13188,a13190,a13192,a13194,a13196,a13198,a13200,a13202,a13204,
a13206,a13208,a13210,a13212,a13214,a13216,a13218,a13220,a13222,a13224,a13226,a13228,a13230,a13232,a13234,
a13236,a13238,a13240,a13242,a13244,a13246,a13248,a13250,a13252,a13254,a13256,a13258,a13260,a13262,a13264,
a13266,a13268,a13270,a13272,a13274,a13276,a13278,a13280,a13282,a13284,a13286,a13288,a13290,a13292,a13294,
a13296,a13298,a13300,a13302,a13304,a13306,a13308,a13310,a13312,a13314,a13316,a13318,a13320,a13322,a13324,
a13326,a13328,a13330,a13332,a13334,a13336,a13338,a13340,a13342,a13344,a13346,a13348,a13350,a13352,a13354,
a13356,a13358,a13360,a13362,a13364,a13366,a13368,a13370,a13372,a13374,a13376,a13378,a13380,a13382,a13384,
a13386,a13388,a13390,a13392,a13394,a13396,a13398,a13400,a13402,a13404,a13406,a13408,a13410,a13412,a13414,
a13416,a13418,a13420,a13422,a13424,a13426,a13428,a13430,a13432,a13434,a13436,a13438,a13440,a13442,a13444,
a13446,a13448,a13450,a13452,a13454,a13456,a13458,a13460,a13462,a13464,a13466,a13468,a13470,a13472,a13474,
a13476,a13478,a13480,a13482,a13484,a13486,a13488,a13490,a13492,a13494,a13496,a13498,a13500,a13502,a13504,
a13506,a13508,a13510,a13512,a13514,a13516,a13518,a13520,a13522,a13524,a13526,a13528,a13530,a13532,a13534,
a13536,a13538,a13540,a13542,a13544,a13546,a13548,a13550,a13552,a13554,a13556,a13558,a13560,a13562,a13564,
a13566,a13568,a13570,a13572,a13574,a13576,a13578,a13580,a13582,a13584,a13586,a13588,a13590,a13592,a13594,
a13596,a13598,a13600,a13602,a13604,a13606,a13608,a13610,a13612,a13614,a13616,a13618,a13620,a13622,a13624,
a13626,a13628,a13630,a13632,a13634,a13636,a13638,a13640,a13642,a13644,a13646,a13648,a13650,a13652,a13654,
a13656,a13658,a13660,a13662,a13664,a13666,a13668,a13670,a13672,a13674,a13676,a13678,a13680,a13682,a13684,
a13686,a13688,a13690,a13692,a13694,a13696,a13698,a13700,a13702,a13704,a13706,a13708,a13710,a13712,a13714,
a13716,a13718,a13720,a13722,a13724,a13726,a13728,a13730,a13732,a13734,a13736,a13738,a13740,a13742,a13744,
a13746,a13748,a13750,a13752,a13754,a13756,a13758,a13760,a13762,a13764,a13766,a13768,a13770,a13772,a13774,
a13776,a13778,a13780,a13782,a13784,a13786,a13788,a13790,a13792,a13794,a13796,a13798,a13800,a13802,a13804,
a13806,a13808,a13810,a13812,a13814,a13816,a13818,a13820,a13822,a13824,a13826,a13828,a13830,a13832,a13834,
a13836,a13838,a13840,a13842,a13844,a13846,a13848,a13850,a13852,a13854,a13856,a13858,a13860,a13862,a13864,
a13866,a13868,a13870,a13872,a13874,a13876,a13878,a13880,a13882,a13884,a13886,a13888,a13890,a13892,a13894,
a13896,a13898,a13900,a13902,a13904,a13906,a13908,a13910,a13912,a13914,a13916,a13918,a13920,a13922,a13924,
a13926,a13928,a13930,a13932,a13934,a13936,a13938,a13940,a13942,a13944,a13946,a13948,a13950,a13952,a13954,
a13956,a13958,a13960,a13962,a13964,a13966,a13968,a13970,a13972,a13974,a13976,a13978,a13980,a13982,a13984,
a13986,a13988,a13990,a13992,a13994,a13996,a13998,a14000,a14002,a14004,a14006,a14008,a14010,a14012,a14014,
a14016,a14018,a14020,a14022,a14024,a14026,a14028,a14030,a14032,a14034,a14036,a14038,a14040,a14042,a14044,
a14046,a14048,a14050,a14052,a14054,a14056,a14058,a14060,a14062,a14064,a14066,a14068,a14070,a14072,a14074,
a14076,a14078,a14080,a14082,a14084,a14086,a14088,a14090,a14092,a14094,a14096,a14098,a14100,a14102,a14104,
a14106,a14108,a14110,a14112,a14114,a14116,a14118,a14120,a14122,a14124,a14126,a14128,a14130,a14132,a14134,
a14136,a14138,a14140,a14142,a14144,a14146,a14148,a14150,a14152,a14154,a14156,a14158,a14160,a14162,a14164,
a14166,a14168,a14170,a14172,a14174,a14176,a14178,a14180,a14182,a14184,a14186,a14188,a14190,a14192,a14194,
a14196,a14198,a14200,a14202,a14204,a14206,a14208,a14210,a14212,a14214,a14216,a14218,a14220,a14222,a14224,
a14226,a14228,a14230,a14232,a14234,a14236,a14238,a14240,a14242,a14244,a14246,a14248,a14250,a14252,a14254,
a14256,a14258,a14260,a14262,a14264,a14266,a14268,a14270,a14272,a14274,a14276,a14278,a14280,a14282,a14284,
a14286,a14288,a14290,a14292,a14294,a14296,a14298,a14300,a14302,a14304,a14306,a14308,a14310,a14312,a14314,
a14316,a14318,a14320,a14322,a14324,a14326,a14328,a14330,a14332,a14334,a14336,a14338,a14340,a14342,a14344,
a14346,a14348,a14350,a14352,a14354,a14356,a14358,a14360,a14362,a14364,a14366,a14368,a14370,a14372,a14374,
a14376,a14378,a14380,a14382,a14384,a14386,a14388,a14390,a14392,a14394,a14396,a14398,a14400,a14402,a14404,
a14406,a14408,a14410,a14412,a14414,a14416,a14418,a14420,a14422,a14424,a14426,a14428,a14430,a14432,a14434,
a14436,a14438,a14440,a14442,a14444,a14446,a14448,a14450,a14452,a14454,a14456,a14458,a14460,a14462,a14464,
a14466,a14468,a14470,a14472,a14474,a14476,a14478,a14480,a14482,a14484,a14486,a14488,a14490,a14492,a14494,
a14496,a14498,a14500,a14502,a14504,a14506,a14508,a14510,a14512,a14514,a14516,a14518,a14520,a14522,a14524,
a14526,a14528,a14530,a14532,a14534,a14536,a14538,a14540,a14542,a14544,a14546,a14548,a14550,a14552,a14554,
a14556,a14558,a14560,a14562,a14564,a14566,a14568,a14570,a14572,a14574,a14576,a14578,a14580,a14582,a14584,
a14586,a14588,a14590,a14592,a14594,a14596,a14598,a14600,a14602,a14604,a14606,a14608,a14610,a14612,a14614,
a14616,a14618,a14620,a14622,a14624,a14626,a14628,a14630,a14632,a14634,a14636,a14638,a14640,a14642,a14644,
a14646,a14648,a14650,a14652,a14654,a14656,a14658,a14660,a14662,a14664,a14666,a14668,a14670,a14672,a14674,
a14676,a14678,a14680,a14682,a14684,a14686,a14688,a14690,a14692,a14694,a14696,a14698,a14700,a14702,a14704,
a14706,a14708,a14710,a14712,a14714,a14716,a14718,a14720,a14722,a14724,a14726,a14728,a14730,a14732,a14734,
a14736,a14738,a14740,a14742,a14744,a14746,a14748,a14750,a14752,a14754,a14756,a14758,a14760,a14762,a14764,
a14766,a14768,a14770,a14772,a14774,a14776,a14778,a14780,a14782,a14784,a14786,a14788,a14790,a14792,a14794,
a14796,a14798,a14800,a14802,a14804,a14806,a14808,a14810,a14812,a14814,a14816,a14818,a14820,a14822,a14824,
a14826,a14828,a14830,a14832,a14834,a14836,a14838,a14840,a14842,a14844,a14846,a14848,a14850,a14852,a14854,
a14856,a14858,a14860,a14862,a14864,a14866,a14868,a14870,a14872,a14874,a14876,a14878,a14880,a14882,a14884,
a14886,a14888,a14890,a14892,a14894,a14896,a14898,a14900,a14902,a14904,a14906,a14908,a14910,a14912,a14914,
a14916,a14918,a14920,a14922,a14924,a14926,a14928,a14930,a14932,a14934,a14936,a14938,a14940,a14942,a14944,
a14946,a14948,a14950,a14952,a14954,a14956,a14958,a14960,a14962,a14964,a14966,a14968,a14970,a14972,a14974,
a14976,a14978,a14980,a14982,a14984,a14986,a14988,a14990,a14992,a14994,a14996,a14998,a15000,a15002,a15004,
a15006,a15008,a15010,a15012,a15014,a15016,a15018,a15020,a15022,a15024,a15026,a15028,a15030,a15032,a15034,
a15036,a15038,a15040,a15042,a15044,a15046,a15048,a15050,a15052,a15054,a15056,a15058,a15060,a15062,a15064,
a15066,a15068,a15070,a15072,a15074,a15076,a15078,a15080,a15082,a15084,a15086,a15088,a15090,a15092,a15094,
a15096,a15098,a15100,a15102,a15104,a15106,a15108,a15110,a15112,a15114,a15116,a15118,a15120,a15122,a15124,
a15126,a15128,a15130,a15132,a15134,a15136,a15138,a15140,a15142,a15144,a15146,a15148,a15150,a15152,a15154,
a15156,a15158,a15160,a15162,a15164,a15166,a15168,a15170,a15172,a15174,a15176,a15178,a15180,a15182,a15184,
a15186,a15188,a15190,a15192,a15194,a15196,a15198,a15200,a15202,a15204,a15206,a15208,a15210,a15212,a15214,
a15216,a15218,a15220,a15222,a15224,a15226,a15228,a15230,a15232,a15234,a15236,a15238,a15240,a15242,a15244,
a15246,a15248,a15250,a15252,a15254,a15256,a15258,a15260,a15262,a15264,a15266,a15268,a15270,a15272,a15274,
a15276,a15278,a15280,a15282,a15284,a15286,a15288,a15290,a15292,a15294,a15296,a15298,a15300,a15302,a15304,
a15306,a15308,a15310,a15312,a15314,a15316,a15318,a15320,a15322,a15324,a15326,a15328,a15330,a15332,a15334,
a15336,a15338,a15340,a15342,a15344,a15346,a15348,a15350,a15352,a15354,a15356,a15358,a15360,a15362,a15364,
a15366,a15368,a15370,a15372,a15374,a15376,a15378,a15380,a15382,a15384,a15386,a15388,a15390,a15392,a15394,
a15396,a15398,a15400,a15402,a15404,a15406,a15408,a15410,a15412,a15414,a15416,a15418,a15420,a15422,a15424,
a15426,a15428,a15430,a15432,a15434,a15436,a15438,a15440,a15442,a15444,a15446,a15448,a15450,a15452,a15454,
a15456,a15458,a15460,a15462,a15464,a15466,a15468,a15470,a15472,a15474,a15476,a15478,a15480,a15482,a15484,
a15486,a15488,a15490,a15492,a15494,a15496,a15498,a15500,a15502,a15504,a15506,a15508,a15510,a15512,a15514,
a15516,a15518,a15520,a15522,a15524,a15526,a15528,a15530,a15532,a15534,a15536,a15538,a15540,a15542,a15544,
a15546,a15548,a15550,a15552,a15554,a15556,a15558,a15560,a15562,a15564,a15566,a15568,a15570,a15572,a15574,
a15576,a15578,a15580,a15582,a15584,a15586,a15588,a15590,a15592,a15594,a15596,a15598,a15600,a15602,a15604,
a15606,a15608,a15610,a15612,a15614,a15616,a15618,a15620,a15622,a15624,a15626,a15628,a15630,a15632,a15634,
a15636,a15638,a15640,a15642,a15644,a15646,a15648,a15650,a15652,a15654,a15656,a15658,a15660,a15662,a15664,
a15666,a15668,a15670,a15672,a15674,a15676,a15678,a15680,a15682,a15684,a15686,a15688,a15690,a15692,a15694,
a15696,a15698,a15700,a15702,a15704,a15706,a15708,a15710,a15712,a15714,a15716,a15718,a15720,a15722,a15724,
a15726,a15728,a15730,a15732,a15734,a15736,a15738,a15740,a15742,a15744,a15746,a15748,a15750,a15752,a15754,
a15756,a15758,a15760,a15762,a15764,a15766,a15768,a15770,a15772,a15774,a15776,a15778,a15780,a15782,a15784,
a15786,a15788,a15790,a15792,a15794,a15796,a15798,a15800,a15802,a15804,a15806,a15808,a15810,a15812,a15814,
a15816,a15818,a15820,a15822,a15824,a15826,a15828,a15830,a15832,a15834,a15836,a15838,a15840,a15842,a15844,
a15846,a15848,a15850,a15852,a15854,a15856,a15858,a15860,a15862,a15864,a15866,a15868,a15870,a15872,a15874,
a15876,a15878,a15880,a15882,a15884,a15886,a15888,a15890,a15892,a15894,a15896,a15898,a15900,a15902,a15904,
a15906,a15908,a15910,a15912,a15914,a15916,a15918,a15920,a15922,a15924,a15926,a15928,a15930,a15932,a15934,
a15936,a15938,a15940,a15942,a15944,a15946,a15948,a15950,a15952,a15954,a15956,a15958,a15960,a15962,a15964,
a15966,a15968,a15970,a15972,a15974,a15976,a15978,a15980,a15982,a15984,a15986,a15988,a15990,a15992,a15994,
a15996,a15998,a16000,a16002,a16004,a16006,a16008,a16010,a16012,a16014,a16016,a16018,a16020,a16022,a16024,
a16026,a16028,a16030,a16032,a16034,a16036,a16038,a16040,a16042,a16044,a16046,a16048,a16050,a16052,a16054,
a16056,a16058,a16060,a16062,a16064,a16066,a16068,a16070,a16072,a16074,a16076,a16078,a16080,a16082,a16084,
a16086,a16088,a16090,a16092,a16094,a16096,a16098,a16100,a16102,a16104,a16106,a16108,a16110,a16112,a16114,
a16116,a16118,a16120,a16122,a16124,a16126,a16128,a16130,a16132,a16134,a16136,a16138,a16140,a16142,a16144,
a16146,a16148,a16150,a16152,a16154,a16156,a16158,a16160,a16162,a16164,a16166,a16168,a16170,a16172,a16174,
a16176,a16178,a16180,a16182,a16184,a16188,a16190,a16192,a16194,a16198,a16200,a16202,a16204,a16206,a16208,
a16210,a16212,a16214,a16216,a16218,a16220,a16222,a16224,a16226,a16228,a16230,a16232,a16234,a16236,a16238,
a16240,a16242,a16244,a16246,a16248,a16252,a16254,a16256,a16258,a16260,a16262,a16264,a16266,a16268,a16270,
a16272,a16274,a16276,a16278,a16280,a16282,a16284,a16286,a16288,a16290,a16292,a16294,a16296,a16298,a16300,
a16302,a16304,a16306,a16308,a16310,a16312,a16314,a16316,a16318,a16320,a16322,a16324,a16326,a16328,a16330,
a16332,a16334,a16336,a16338,a16340,a16342,a16344,a16346,a16348,a16350,a16352,a16354,a16356,a16358,a16360,
a16362,a16364,a16366,a16368,a16370,a16372,a16374,a16376,a16378,a16380,a16382,a16384,a16386,a16388,a16390,
a16392,a16394,a16396,a16398,a16400,a16402,a16404,a16406,a16408,a16410,a16412,a16414,a16416,a16418,a16420,
a16422,a16424,a16426,a16428,a16430,a16432,a16434,a16436,a16438,a16442,a16444,a16446,a16448,a16450,a16452,
a16454,a16456,a16458,a16460,a16462,a16464,a16466,a16468,a16470,a16472,a16474,a16476,a16478,a16480,a16482,
a16484,a16486,a16488,a16490,a16492,a16494,a16496,a16498,a16500,a16502,a16504,a16506,a16508,a16510,a16512,
a16516,a16518,a16520,a16522,a16524,a16526,a16528,a16530,a16532,a16534,a16536,a16538,a16540,a16542,a16544,
a16546,a16548,a16550,a16552,a16554,a16556,a16558,a16560,a16562,a16564,a16566,a16568,a16570,a16572,a16574,
a16576,a16578,a16582,a16584,a16586,a16588,a16590,a16592,a16594,a16596,a16598,a16600,a16602,a16604,a16606,
a16610,a16612,a16614,a16616,a16618,a16620,a16622,a16624,a16626,a16628,a16630,a16632,a16634,a16636,a16638,
a16640,a16642,a16644,a16646,a16648,a16650,a16652,a16654,a16656,a16658,a16660,a16662,a16664,a16666,a16668,
a16670,a16672,a16674,a16676,a16678,a16680,a16682,a16686,a16688,a16690,a16692,a16694,a16696,a16698,a16700,
a16702,a16704,a16706,a16708,a16710,a16714,a16716,a16718,a16720,a16722,a16724,a16726,a16728,a16730,a16732,
a16734,a16736,a16738,a16740,a16742,a16744,a16746,a16748,a16750,a16752,a16754,a16756,a16758,a16760,a16762,
a16764,a16766,a16768,a16770,a16772,a16774,a16776,a16778,a16780,a16782,a16784,a16786,a16790,a16792,a16794,
a16796,a16798,a16800,a16802,a16804,a16806,a16808,a16810,a16812,a16814,a16818,a16820,a16822,a16824,a16826,
a16828,a16830,a16832,a16834,a16836,a16838,a16840,a16842,a16844,a16846,a16848,a16850,a16852,a16854,a16856,
a16858,a16860,a16862,a16864,a16866,a16868,a16870,a16872,a16874,a16876,a16878,a16880,a16882,a16884,a16886,
a16888,a16890,a16894,a16896,a16898,a16900,a16902,a16904,a16906,a16908,a16910,a16912,a16914,a16916,a16918,
a16922,a16924,a16926,a16928,a16930,a16932,a16934,a16936,a16938,a16940,a16942,a16944,a16946,a16948,a16950,
a16952,a16954,a16956,a16958,a16960,a16962,a16964,a16966,a16968,a16970,a16972,a16974,a16976,a16978,a16980,
a16982,a16984,a16986,a16988,a16990,a16992,a16994,a16998,a17000,a17002,a17004,a17006,a17008,a17010,a17012,
a17014,a17016,a17018,a17020,a17022,a17024,a17026,a17028,a17030,a17032,a17034,a17036,a17038,a17040,a17042,
a17044,a17046,a17048,a17050,a17052,a17054,a17056,a17058,a17060,a17062,a17064,a17066,a17068,a17070,a17072,
a17074,a17076,a17078,a17080,a17082,a17084,a17086,a17088,a17090,a17092,a17094,a17096,a17098,a17100,a17102,
a17104,a17106,a17108,a17110,a17112,a17114,a17116,a17118,a17120,a17122,a17124,a17126,a17128,a17130,a17132,
a17134,a17136,a17138,a17140,a17142,a17144,a17146,a17148,a17150,a17152,a17154,a17156,a17158,a17160,a17162,
a17164,a17166,a17168,a17170,a17172,a17174,a17176,a17178,a17180,a17182,a17184,a17186,a17188,a17190,a17192,
a17194,a17196,a17198,a17200,a17202,a17204,a17206,a17208,a17210,a17212,a17214,a17216,a17218,a17220,a17222,
a17224,a17226,a17228,a17230,a17232,a17234,a17236,a17238,a17240,a17242,a17244,a17246,a17248,a17250,a17252,
a17254,a17256,a17258,a17260,a17262,a17264,a17266,a17268,a17270,a17272,a17274,a17276,a17278,a17280,a17282,
a17284,a17286,a17288,a17290,a17292,a17294,a17296,a17298,a17300,a17302,a17304,a17306,a17308,a17310,a17312,
a17314,a17316,a17318,a17320,a17322,a17324,a17326,a17328,a17330,a17332,a17334,a17336,a17338,a17340,a17342,
a17344,a17346,a17348,a17350,a17352,a17354,a17356,a17358,a17360,a17362,a17364,a17366,a17368,a17370,a17372,
a17374,a17376,a17378,a17380,a17382,a17384,a17386,a17388,a17390,a17392,a17394,a17396,a17398,a17400,a17402,
a17404,a17406,a17408,a17410,a17412,a17414,a17416,a17418,a17420,a17422,a17424,a17426,a17428,a17430,a17432,
a17434,a17436,a17438,a17440,a17442,a17444,a17446,a17448,a17450,a17452,a17454,a17456,a17458,a17460,a17462,
a17464,a17466,a17468,a17470,a17472,a17474,a17476,a17478,a17480,a17482,a17484,a17486,a17488,a17490,a17492,
a17494,a17496,a17498,a17500,a17502,a17504,a17506,a17508,a17510,a17512,a17514,a17516,a17518,a17520,a17522,
a17524,a17526,a17528,a17530,a17532,a17534,a17536,a17538,a17540,a17542,a17544,a17546,a17548,a17550,a17552,
a17554,a17556,a17558,a17560,a17562,a17564,a17566,a17568,a17570,a17572,a17574,a17576,a17578,a17580,a17582,
a17584,a17586,a17588,a17590,a17592,a17594,a17596,a17598,a17600,a17602,a17604,a17606,a17608,a17610,a17612,
a17614,a17616,a17618,a17620,a17622,a17624,a17626,a17628,a17630,a17632,a17634,a17636,a17638,a17640,a17642,
a17644,a17646,a17648,a17650,a17652,a17654,a17656,a17658,a17660,a17662,a17664,a17666,a17668,a17670,a17672,
a17674,a17676,a17678,a17680,a17684,a17686,a17688,a17690,a17692,a17694,a17696,a17698,a17700,a17702,a17704,
a17706,a17708,a17710,a17712,a17714,a17716,a17718,a17720,a17722,a17724,a17726,a17728,a17730,a17732,a17734,
a17736,a17738,a17740,a17742,a17744,a17746,a17748,a17750,a17752,a17754,a17756,a17758,a17760,a17762,a17764,
a17766,a17768,a17770,a17772,a17774,a17776,a17778,a17780,a17782,a17784,a17786,a17788,a17790,a17792,a17794,
a17796,a17798,a17800,a17802,a17804,a17806,a17808,a17810,a17812,a17814,a17816,a17818,a17820,a17822,a17824,
a17826,a17828,a17830,a17832,a17834,a17836,a17838,a17840,a17842,a17844,a17846,a17848,a17850,a17852,a17854,
a17856,a17858,a17860,a17862,a17864,a17866,a17868,a17870,a17872,a17874,a17876,a17878,a17880,a17882,a17884,
a17886,a17888,a17890,a17892,a17894,a17896,a17898,a17900,a17902,a17904,a17906,a17908,a17910,a17912,a17914,
a17916,a17918,a17920,a17922,a17924,a17926,a17928,a17930,a17932,a17934,a17936,a17938,a17940,a17942,a17944,
a17946,a17948,a17950,a17952,a17954,a17956,a17958,a17960,a17962,a17964,a17966,a17968,a17970,a17972,a17974,
a17976,a17978,a17980,a17982,a17984,a17986,a17988,a17990,a17992,a17994,a17996,a17998,a18000,a18002,a18004,
a18006,a18008,a18010,a18012,a18014,a18016,a18018,a18020,a18022,a18024,a18026,a18028,a18030,a18032,a18034,
a18036,a18038,a18040,a18042,a18044,a18046,a18048,a18050,a18052,a18054,a18056,a18058,a18060,a18062,a18064,
a18066,a18068,a18070,a18072,a18074,a18076,a18078,a18080,a18082,a18084,a18086,a18088,a18090,a18092,a18094,
a18096,a18098,a18100,a18102,a18104,a18106,a18108,a18110,a18112,a18114,a18116,a18118,a18120,a18122,a18124,
a18126,a18128,a18130,a18132,a18134,a18136,a18138,a18140,a18142,a18144,a18146,a18148,a18150,a18152,a18154,
a18156,a18158,a18160,a18162,a18164,a18166,a18168,a18170,a18172,a18174,a18176,a18178,a18180,a18182,a18184,
a18186,a18188,a18190,a18192,a18194,a18196,a18198,a18200,a18202,a18204,a18206,a18208,a18210,a18212,a18214,
a18216,a18218,a18220,a18222,a18224,a18226,a18228,a18230,a18232,a18234,a18236,a18238,a18240,a18242,a18244,
a18246,a18248,a18250,a18252,a18254,a18256,a18258,a18260,a18262,a18264,a18266,a18268,a18270,a18272,a18274,
a18276,a18278,a18280,a18282,a18284,a18286,a18288,a18290,a18292,a18294,a18296,a18298,a18300,a18302,a18304,
a18306,a18308,a18310,a18312,a18314,a18316,a18318,a18320,a18322,a18324,a18326,a18328,a18330,a18332,a18334,
a18336,a18338,a18340,a18342,a18344,a18346,a18348,a18350,a18352,a18354,a18356,a18358,a18360,a18362,a18364,
a18366,a18368,a18370,a18372,a18374,a18376,a18378,a18380,a18382,a18384,a18386,a18388,a18390,a18392,a18394,
a18396,a18398,a18400,a18402,a18404,a18406,a18408,a18410,a18412,a18414,a18416,a18418,a18420,a18422,a18424,
a18426,a18428,a18430,a18432,a18434,a18436,a18438,a18440,a18442,a18444,a18446,a18448,a18450,a18452,a18454,
a18456,a18458,a18460,a18462,a18464,a18466,a18468,a18470,a18472,a18474,a18476,a18478,a18480,a18482,a18484,
a18486,a18488,a18490,a18492,a18494,a18496,a18498,a18500,a18502,a18504,a18506,a18508,a18510,a18512,a18516,
a18518,a18522,a18524,a18526,a18528,a18530,a18532,a18534,a18536,a18538,a18540,a18544,a18546,a18548,a18550,
a18552,a18554,a18558,a18560,a18564,a18566,a18568,a18570,a18572,a18574,a18576,a18578,a18580,a18582,a18584,
a18586,a18588,a18590,a18592,a18594,a18596,a18598,a18600,a18602,a18604,a18606,a18608,a18610,a18612,a18614,
a18616,a18618,a18620,a18622,a18624,a18626,a18628,a18630,a18632,a18634,a18636,a18638,a18640,a18642,a18644,
a18646,a18648,a18650,a18652,a18654,a18656,a18658,a18660,a18662,a18664,a18666,a18668,a18670,a18672,a18674,
a18676,a18678,a18680,a18682,a18684,a18686,a18688,a18690,a18692,a18694,a18696,a18698,a18700,a18702,a18704,
a18706,a18708,a18710,a18712,a18714,a18716,a18718,a18720,a18722,a18724,a18726,a18728,a18730,a18732,a18734,
a18736,a18738,a18740,a18742,a18744,a18746,a18748,a18750,a18752,a18754,a18756,a18758,a18760,a18762,a18764,
a18766,a18768,a18770,a18772,a18774,a18776,a18778,a18780,a18782,a18784,a18786,a18788,a18790,a18792,a18794,
a18796,a18798,a18800,a18802,a18804,a18806,a18808,a18810,a18812,a18814,a18816,a18818,a18820,a18822,a18824,
a18826,a18828,a18830,a18832,a18834,a18836,a18838,a18840,a18842,a18844,a18846,a18848,a18852,a18854,a18856,
a18858,a18860,a18862,a18864,a18866,a18868,a18870,a18872,a18874,a18876,a18878,a18880,a18882,a18884,a18886,
a18888,a18890,a18892,a18894,a18896,a18898,a18900,a18902,a18904,a18906,a18908,a18910,a18912,a18914,a18916,
a18918,a18920,a18922,a18926,a18928,a18930,a18932,a18934,a18936,a18938,a18940,a18942,a18944,a18946,a18948,
a18950,a18952,a18954,a18956,a18958,a18960,a18962,a18964,a18966,a18968,a18970,a18972,a18974,a18976,a18978,
a18980,a18982,a18984,a18986,a18988,a18990,a18992,a18994,a18996,a18998,a19000,a19002,a19006,a19008,a19010,
a19012,a19014,a19016,a19018,a19020,a19022,a19024,a19026,a19028,a19030,a19032,a19034,a19036,a19038,a19040,
a19042,a19044,a19046,a19048,a19050,a19052,a19054,a19056,a19058,a19060,a19062,a19064,a19066,a19068,a19070,
a19072,a19074,a19076,a19078,a19080,a19082,a19084,a19088,a19090,a19092,a19094,a19096,a19098,a19100,a19102,
a19104,a19106,a19108,a19110,a19112,a19114,a19116,a19118,a19120,a19122,a19124,a19126,a19128,a19130,a19132,
a19134,a19136,a19138,a19140,a19142,a19144,a19146,a19148,a19150,a19152,a19154,a19156,a19158,a19160,a19162,
a19164,a19166,a19170,a19172,a19174,a19176,a19178,a19180,a19182,a19184,a19186,a19188,a19190,a19192,a19194,
a19196,a19198,a19200,a19202,a19204,a19206,a19208,a19210,a19212,a19214,a19216,a19218,a19220,a19222,a19224,
a19226,a19228,a19230,a19232,a19234,a19236,a19238,a19240,a19242,a19244,a19246,a19248,a19250,a19252,a19254,
a19256,a19258,a19260,a19262,a19264,a19266,a19268,a19270,a19272,a19274,a19276,a19278,a19280,a19282,a19284,
a19286,a19288,a19290,a19292,a19294,a19296,a19298,a19300,a19302,a19304,a19306,a19308,a19310,a19312,a19314,
a19316,a19318,a19320,a19322,a19324,a19326,a19328,a19330,a19332,a19334,a19336,a19338,a19340,a19342,a19344,
a19346,a19348,a19350,a19352,a19354,a19356,a19358,a19360,a19362,a19364,a19366,a19368,a19370,a19372,a19374,
a19376,a19378,a19380,a19382,a19384,a19386,a19388,a19390,a19392,a19394,a19396,a19398,a19400,a19402,a19404,
a19406,a19408,a19410,a19412,a19414,a19416,a19418,a19420,a19422,a19424,a19426,a19428,a19430,a19432,a19434,
a19436,a19438,a19440,a19442,a19444,a19446,a19448,a19450,a19452,a19454,a19456,a19458,a19460,a19462,a19464,
a19466,a19468,a19470,a19472,a19474,a19476,a19478,a19480,a19482,a19484,a19486,a19488,a19490,a19492,a19494,
a19496,a19498,a19500,a19502,a19504,a19506,a19508,a19510,a19512,a19514,a19516,a19518,a19520,a19522,a19524,
a19526,a19528,a19530,a19532,a19534,a19536,a19538,a19540,a19542,a19544,a19546,a19548,a19550,a19552,a19554,
a19556,a19558,a19560,a19562,a19564,a19566,a19568,a19570,a19572,a19574,a19576,a19578,a19580,a19582,a19584,
a19586,a19588,a19590,a19592,a19594,a19596,a19598,a19600,a19602,a19604,a19606,a19608,a19610,a19612,a19614,
a19616,a19618,a19620,a19622,a19624,a19626,a19628,a19630,a19632,a19634,a19636,a19638,a19640,a19642,a19644,
a19646,a19648,a19650,a19652,a19654,a19656,a19658,a19660,a19662,a19664,a19666,a19668,a19670,a19672,a19674,
a19676,a19678,a19680,a19682,a19684,a19686,a19688,a19690,a19692,a19694,a19696,a19698,a19700,a19702,a19704,
a19706,a19708,a19710,a19712,a19714,a19716,a19718,a19720,a19722,a19724,a19726,a19728,a19730,a19732,a19734,
a19736,a19738,a19740,a19742,a19744,a19746,a19748,a19750,a19752,a19754,a19758,a19760,a19762,a19764,a19766,
a19768,a19770,a19772,a19774,a19776,a19778,a19780,a19782,a19784,a19786,a19788,a19790,a19792,a19794,a19796,
a19798,a19800,a19802,a19804,a19806,a19808,a19810,a19812,a19814,a19816,a19818,a19820,a19822,a19824,a19826,
a19828,a19830,a19832,a19834,a19836,a19838,a19840,a19842,a19844,a19846,a19848,a19850,a19852,a19854,a19856,
a19858,a19860,a19862,a19864,a19866,a19868,a19870,a19872,a19874,a19876,a19878,a19880,a19882,a19884,a19886,
a19888,a19890,a19896,a19898,a19902,a19904,a19906,a19908,a19910,a19912,a19914,a19916,a19918,a19920,a19922,
a19924,a19926,a19928,a19930,a19932,a19934,a19936,a19938,a19940,a19942,a19944,a19946,a19948,a19950,a19952,
a19954,a19956,a19958,a19960,a19962,a19964,a19966,a19968,a19970,a19972,a19974,a19978,a19980,a19982,a19984,
a19986,a19988,a19990,a19992,a19994,a19996,a19998,a20000,a20004,a20006,a20008,a20010,a20012,a20014,a20016,
a20018,a20020,a20022,a20024,a20026,a20030,a20032,a20034,a20036,a20038,a20040,a20042,a20044,a20046,a20048,
a20050,a20052,a20056,a20058,a20060,a20062,a20064,a20066,a20068,a20070,a20072,a20074,a20076,a20080,a20082,
a20084,a20086,a20088,a20090,a20092,a20094,a20096,a20098,a20100,a20102,a20104,a20106,a20108,a20110,a20112,
a20114,a20116,a20118,a20120,a20122,a20124,a20126,a20128,a20130,a20132,a20134,a20136,a20138,a20140,a20142,
a20144,a20146,a20148,a20150,a20152,a20154,a20156,a20158,a20160,a20162,a20164,a20166,a20168,a20170,a20172,
a20174,a20176,a20178,a20180,a20182,a20184,a20186,a20188,a20190,a20192,a20194,a20196,a20198,a20200,a20202,
a20204,a20206,a20208,a20210,a20212,a20214,a20216,a20218,a20220,a20222,a20224,a20226,a20228,a20230,a20232,
a20234,a20236,a20238,a20240,a20242,a20244,a20246,a20248,a20250,a20252,a20254,a20256,a20258,a20260,a20262,
a20264,a20266,a20268,a20270,a20272,a20274,a20276,a20278,a20280,a20282,a20284,a20286,a20288,a20290,a20292,
a20294,a20296,a20298,a20300,a20302,a20304,a20306,a20308,a20310,a20312,a20314,a20316,a20318,a20320,a20322,
a20324,a20326,a20328,a20330,a20332,a20334,a20336,a20338,a20340,a20342,a20344,a20346,a20348,a20350,a20352,
a20354,a20356,a20358,a20360,a20362,a20364,a20366,a20368,a20370,a20372,a20374,a20376,a20378,a20380,a20382,
a20384,a20386,a20388,a20390,a20392,a20394,a20396,a20398,a20400,a20402,a20404,a20406,a20408,a20410,a20412,
a20414,a20416,a20418,a20420,a20422,a20424,a20426,a20428,a20430,a20432,a20434,a20436,a20438,a20440,a20442,
a20444,a20446,a20448,a20450,a20452,a20454,a20456,a20458,a20460,a20462,a20464,a20466,a20468,a20470,a20472,
a20474,a20476,a20478,a20480,a20482,a20484,a20486,a20488,a20490,a20492,a20494,a20496,a20498,a20500,a20502,
a20504,a20506,a20508,a20510,a20512,a20514,a20516,a20518,a20520,a20522,a20524,a20526,a20528,a20530,a20532,
a20534,a20536,a20538,a20540,a20542,a20544,a20546,a20548,a20550,a20552,a20554,a20556,a20558,a20560,a20562,
a20564,a20566,a20568,a20570,a20572,a20574,a20576,a20578,a20580,a20582,a20584,a20586,a20588,a20590,a20592,
a20594,a20596,a20598,a20600,a20602,a20604,a20606,a20608,a20610,a20612,a20614,a20616,a20618,a20620,a20622,
a20624,a20626,a20628,a20630,a20632,a20634,a20636,a20638,a20640,a20642,a20644,a20646,a20648,a20650,a20652,
a20654,a20656,a20658,a20660,a20662,a20664,a20666,a20668,a20670,a20672,a20674,a20676,a20678,a20680,a20682,
a20684,a20686,a20688,a20690,a20692,a20694,a20696,a20698,a20700,a20702,a20704,a20706,a20708,a20710,a20712,
a20714,a20716,a20718,a20720,a20722,a20724,a20726,a20728,a20730,a20732,a20734,a20736,a20738,a20740,a20742,
a20744,a20746,a20748,a20750,a20752,a20754,a20756,a20758,a20760,a20762,a20764,a20766,a20768,a20770,a20772,
a20774,a20776,a20778,a20780,a20782,a20784,a20786,a20788,a20790,a20792,a20794,a20796,a20798,a20800,a20802,
a20804,a20806,a20808,a20810,a20812,a20814,a20816,a20818,a20820,a20822,a20824,a20826,a20828,a20830,a20832,
a20834,a20836,a20838,a20840,a20842,a20844,a20846,a20848,a20850,a20852,a20854,a20856,a20858,a20860,a20862,
a20864,a20866,a20868,a20870,a20872,a20874,a20876,a20878,a20880,a20882,a20884,a20886,a20888,a20890,a20892,
a20894,a20896,a20898,a20900,a20902,a20904,a20906,a20908,a20910,a20912,a20914,a20916,a20918,a20920,a20922,
a20924,a20926,a20928,a20930,a20932,a20934,a20936,a20938,a20940,a20942,a20944,a20946,a20948,a20950,a20952,
a20954,a20956,a20958,a20960,a20962,a20964,a20966,a20968,a20970,a20972,a20974,a20976,a20978,a20980,a20982,
a20984,a20986,a20988,a20990,a20992,a20994,a20996,a20998,a21000,a21002,a21004,a21006,a21008,a21010,a21012,
a21014,a21016,a21018,a21020,a21022,a21024,a21026,a21028,a21030,a21032,a21034,a21036,a21038,a21040,a21042,
a21044,a21046,a21048,a21050,a21052,a21054,a21056,a21058,a21060,a21062,a21064,a21066,a21068,a21070,a21072,
a21074,a21076,a21078,a21080,a21082,a21084,a21086,a21088,a21090,a21092,a21094,a21096,a21098,a21100,a21102,
a21104,a21106,a21108,a21110,a21112,a21114,a21116,a21118,a21120,a21122,a21124,a21126,a21128,a21130,a21132,
a21134,a21136,a21138,a21140,a21142,a21144,a21146,a21148,a21150,a21152,a21154,a21156,a21158,a21160,a21162,
a21164,a21166,a21168,a21170,a21172,a21174,a21176,a21178,a21180,a21182,a21184,a21186,a21188,a21190,a21192,
a21194,a21196,a21198,a21200,a21202,a21204,a21206,a21208,a21210,a21212,a21214,a21216,a21218,a21220,a21222,
a21224,a21226,a21228,a21230,a21232,a21234,a21236,a21238,a21240,a21242,a21244,a21246,a21248,a21250,a21252,
a21254,a21256,a21258,a21260,a21262,a21264,a21266,a21268,a21270,a21272,a21274,a21276,a21278,a21280,a21282,
a21284,a21286,a21288,a21290,a21292,a21294,a21296,a21298,a21300,a21302,a21304,a21306,a21308,a21310,a21312,
a21314,a21316,a21318,a21320,a21322,a21324,a21326,a21328,a21330,a21332,a21334,a21336,a21338,a21340,a21342,
a21344,a21346,a21348,a21350,a21352,a21354,a21356,a21358,a21360,a21362,a21364,a21366,a21368,a21370,a21372,
a21374,a21376,a21378,a21380,a21382,a21384,a21386,a21388,a21390,a21392,a21394,a21396,a21398,a21400,a21402,
a21404,a21406,a21408,a21410,a21412,a21414,a21416,a21418,a21420,a21422,a21424,a21426,a21428,a21430,a21432,
a21434,a21436,a21438,a21440,a21442,a21444,a21446,a21448,a21450,a21452,a21454,a21456,a21458,a21460,a21462,
a21464,a21466,a21468,a21470,a21472,a21474,a21476,a21478,a21480,a21482,a21484,a21486,a21488,a21490,a21492,
a21494,a21496,a21498,a21500,a21502,a21504,a21506,a21508,a21510,a21512,a21514,a21516,a21518,a21520,a21522,
a21524,a21526,a21528,a21530,a21532,a21534,a21536,a21538,a21540,a21542,a21544,a21546,a21548,a21550,a21552,
a21554,a21556,a21558,a21560,a21562,a21564,a21566,a21568,a21570,a21572,a21574,a21576,a21578,a21580,a21582,
a21584,a21586,a21588,a21590,a21592,a21594,a21596,a21598,a21600,a21602,a21604,a21606,a21608,a21610,a21612,
a21614,a21616,a21618,a21620,a21622,a21624,a21626,a21628,a21630,a21632,a21634,a21636,a21638,a21640,a21642,
a21644,a21646,a21648,a21650,a21652,a21654,a21656,a21658,a21660,a21662,a21666,a21668,a21672,a21674,a21676,
a21678,a21680,a21682,a21684,a21686,a21688,a21690,a21692,a21694,a21696,a21698,a21700,a21702,a21704,a21706,
a21708,a21710,a21712,a21714,a21716,a21718,a21720,a21722,a21724,a21726,a21728,a21730,a21732,a21734,a21736,
a21738,a21740,a21742,a21744,a21746,a21748,a21750,a21752,a21754,a21756,a21758,a21760,a21762,a21764,a21766,
a21768,a21770,a21772,a21774,a21776,a21778,a21780,a21782,a21784,a21786,a21788,a21790,a21792,a21794,a21796,
a21798,a21802,a21804,a21806,a21808,a21812,a21814,a21816,a21818,a21820,a21822,a21824,a21826,a21830,a21832,
a21834,a21836,a21838,a21840,a21842,a21844,a21846,a21848,a21850,a21852,a21854,a21856,a21858,a21860,a21862,
a21864,a21866,a21868,a21870,a21872,a21874,a21876,a21878,a21882,a21884,a21886,a21888,a21890,a21892,a21894,
a21896,a21898,a21900,a21902,a21904,a21906,a21908,a21910,a21912,a21914,a21916,a21918,a21920,a21922,a21924,
a21926,a21928,a21930,a21932,a21934,a21936,a21938,a21940,a21942,a21944,a21946,a21948,a21952,a21954,a21956,
a21960,a21962,a21964,a21966,a21968,a21972,a21974,a21976,a21978,a21980,a21982,a21984,a21986,a21988,a21990,
a21992,a21994,a21996,a21998,a22000,a22002,a22004,a22006,a22008,a22010,a22012,a22016,a22018,a22020,a22022,
a22024,a22026,a22028,a22030,a22032,a22034,a22036,a22038,a22040,a22042,a22044,a22046,a22048,a22050,a22052,
a22054,a22056,a22058,a22060,a22062,a22064,a22066,a22068,a22070,a22072,a22074,a22076,a22078,a22080,a22082,
a22086,a22088,a22090,a22094,a22096,a22098,a22100,a22102,a22106,a22108,a22110,a22112,a22114,a22116,a22118,
a22120,a22122,a22124,a22126,a22128,a22130,a22132,a22134,a22136,a22138,a22140,a22142,a22144,a22146,a22150,
a22152,a22154,a22156,a22158,a22160,a22162,a22164,a22166,a22168,a22170,a22172,a22174,a22176,a22178,a22180,
a22182,a22184,a22186,a22188,a22190,a22192,a22194,a22196,a22198,a22200,a22202,a22204,a22206,a22208,a22210,
a22212,a22214,a22216,a22220,a22222,a22224,a22228,a22230,a22232,a22234,a22236,a22240,a22242,a22244,a22246,
a22248,a22250,a22252,a22254,a22256,a22258,a22260,a22262,a22264,a22266,a22268,a22270,a22272,a22274,a22276,
a22278,a22280,a22284,a22286,a22288,a22290,a22292,a22294,a22296,a22298,a22300,a22302,a22304,a22306,a22308,
a22310,a22312,a22314,a22316,a22318,a22320,a22322,a22324,a22326,a22328,a22330,a22332,a22334,a22336,a22338,
a22340,a22342,a22344,a22346,a22348,a22350,a22354,a22356,a22358,a22362,a22364,a22366,a22368,a22370,a22374,
a22376,a22378,a22380,a22382,a22384,a22386,a22388,a22390,a22392,a22394,a22396,a22398,a22400,a22402,a22404,
a22406,a22408,a22410,a22412,a22414,a22418,a22420,a22422,a22424,a22426,a22428,a22430,a22432,a22434,a22436,
a22438,a22440,a22442,a22444,a22446,a22448,a22450,a22452,a22454,a22456,a22458,a22460,a22462,a22464,a22466,
a22468,a22470,a22472,a22474,a22476,a22478,a22480,a22482,a22484,a22488,a22490,a22492,a22496,a22498,a22500,
a22502,a22504,a22508,a22510,a22512,a22514,a22516,a22518,a22520,a22522,a22524,a22526,a22528,a22530,a22532,
a22534,a22536,a22538,a22540,a22542,a22544,a22546,a22548,a22552,a22554,a22556,a22558,a22560,a22562,a22564,
a22566,a22568,a22570,a22572,a22574,a22576,a22578,a22580,a22582,a22584,a22586,a22588,a22590,a22592,a22594,
a22596,a22598,a22600,a22602,a22604,a22606,a22608,a22610,a22612,a22614,a22616,a22618,a22622,a22624,a22626,
a22630,a22632,a22634,a22636,a22638,a22640,a22642,a22644,a22646,a22648,a22650,a22652,a22654,a22656,a22658,
a22660,a22662,a22664,a22666,a22668,a22670,a22672,a22674,a22676,a22678,a22680,a22682,a22684,a22686,a22688,
a22690,a22692,a22694,a22696,a22698,a22700,a22702,a22704,a22706,a22708,a22710,a22712,a22714,a22716,a22718,
a22720,a22722,a22724,a22726,a22728,a22730,a22732,a22734,a22736,a22738,a22740,a22742,a22744,a22746,a22748,
a22750,a22752,a22754,a22756,a22758,a22760,a22762,a22764,a22766,a22768,a22770,a22772,a22774,a22776,a22778,
a22780,a22782,a22784,a22786,a22788,a22790,a22792,a22794,a22796,a22798,a22800,a22802,a22804,a22806,a22810,
a22812,a22814,a22816,a22818,a22820,a22822,a22824,a22826,a22828,a22830,a22832,a22834,a22836,a22838,a22840,
a22842,a22844,a22846,a22848,a22850,a22852,a22854,a22856,a22858,a22860,a22862,a22864,a22866,a22868,a22870,
a22872,a22874,a22876,a22878,a22880,a22882,a22884,a22886,a22888,a22890,a22892,a22894,a22896,a22898,a22900,
a22902,a22904,a22906,a22908,a22910,a22912,a22914,a22916,a22918,a22920,a22922,a22924,a22926,a22928,a22930,
a22932,a22934,a22936,a22938,a22940,a22942,a22944,a22946,a22948,a22950,a22952,a22954,a22956,a22958,a22960,
a22962,a22964,a22966,a22968,a22970,a22972,a22974,a22976,a22978,a22980,a22982,a22984,a22986,a22988,a22990,
a22992,a22994,a22996,a22998,a23000,a23002,a23004,a23006,a23008,a23010,a23012,a23014,a23016,a23018,a23020,
a23022,a23024,a23026,a23028,a23030,a23032,a23034,a23036,a23038,a23040,a23042,a23044,a23046,a23048,a23050,
a23052,a23054,a23056,a23058,a23060,a23062,a23064,a23066,a23068,a23070,a23072,a23074,a23076,a23078,a23080,
a23082,a23084,a23086,a23088,a23090,a23092,a23094,a23096,a23098,a23100,a23102,a23104,a23106,a23108,a23110,
a23112,a23114,a23116,a23118,a23120,a23122,a23124,a23126,a23128,a23130,a23132,a23134,a23136,a23138,a23140,
a23142,a23144,a23146,a23148,a23150,a23152,a23154,a23156,a23158,a23160,a23162,a23164,a23166,a23168,a23170,
a23172,a23174,a23176,a23178,a23180,a23182,a23184,a23186,a23188,a23190,a23192,a23194,a23196,a23198,a23200,
a23202,a23204,a23206,a23208,a23210,a23212,a23214,a23216,a23218,a23220,a23222,a23224,a23226,a23228,a23230,
a23232,a23234,a23236,a23238,a23240,a23242,a23244,a23246,a23248,a23250,a23252,a23254,a23256,a23258,a23260,
a23262,a23264,a23266,a23268,a23270,a23272,a23274,a23276,a23278,a23280,a23282,a23284,a23286,a23288,a23290,
a23292,a23294,a23296,a23298,a23300,a23302,a23304,a23306,a23308,a23310,a23312,a23314,a23316,a23318,a23320,
a23322,a23324,a23326,a23328,a23330,a23332,a23334,a23336,a23338,a23340,a23342,a23344,a23346,a23348,a23350,
a23352,a23354,a23356,a23358,a23360,a23362,a23364,a23366,a23368,a23370,a23372,a23374,a23376,a23378,a23380,
a23382,a23384,a23386,a23388,a23390,a23392,a23394,a23396,a23398,a23400,a23402,a23404,a23406,a23408,a23410,
a23412,a23414,a23416,a23418,a23420,a23422,a23424,a23426,a23428,a23430,a23432,a23434,a23436,a23438,a23440,
a23442,a23444,a23446,a23448,a23450,a23452,a23454,a23456,a23458,a23460,a23462,a23464,a23466,a23468,a23470,
a23472,a23474,a23476,a23478,a23480,a23482,a23484,a23486,a23488,a23490,a23492,a23494,a23496,a23498,a23500,
a23502,a23504,a23506,a23508,a23510,a23512,a23514,a23516,a23518,a23520,a23522,a23524,a23526,a23528,a23530,
a23532,a23534,a23536,a23538,a23540,a23542,a23544,a23546,a23548,a23550,a23552,a23554,a23556,a23558,a23560,
a23562,a23564,a23566,a23568,a23570,a23572,a23574,a23576,a23578,a23580,a23582,a23584,a23586,a23588,a23590,
a23592,a23594,a23596,a23598,a23600,a23602,a23604,a23606,a23608,a23610,a23612,a23614,a23616,a23618,a23620,
a23622,a23624,a23626,a23628,a23630,a23632,a23634,a23636,a23638,a23640,a23642,a23644,a23646,a23648,a23650,
a23652,a23654,a23656,a23658,a23660,a23662,a23664,a23666,a23668,a23670,a23672,a23674,a23676,a23678,a23680,
a23682,a23684,a23686,a23688,a23690,a23692,a23694,a23696,a23698,a23700,a23702,a23704,a23706,a23708,a23710,
a23712,a23714,a23716,a23718,a23720,a23722,a23724,a23726,a23728,a23730,a23732,a23734,a23738,a23740,a23744,
a23746,a23748,a23750,a23752,a23754,a23756,a23758,a23760,a23762,a23764,a23766,a23768,a23770,a23772,a23774,
a23776,a23778,a23780,a23782,a23784,a23786,a23788,a23790,a23792,a23794,a23796,a23798,a23800,a23802,a23804,
a23806,a23808,a23810,a23812,a23814,a23816,a23818,a23820,a23822,a23824,a23826,a23828,a23830,a23832,a23834,
a23836,a23838,a23840,a23842,a23844,a23846,a23848,a23850,a23852,a23854,a23856,a23858,a23860,a23862,a23864,
a23866,a23868,a23870,a23872,a23874,a23876,a23878,a23880,a23882,a23884,a23886,a23888,a23890,a23892,a23894,
a23896,a23898,a23900,a23902,a23904,a23906,a23908,a23910,a23912,a23914,a23916,a23918,a23920,a23922,a23924,
a23926,a23928,a23930,a23932,a23934,a23936,a23938,a23940,a23942,a23944,a23946,a23948,a23950,a23952,a23954,
a23956,a23958,a23960,a23962,a23964,a23966,a23968,a23970,a23972,a23974,a23976,a23978,a23980,a23982,a23984,
a23986,a23988,a23990,a23992,a23994,a23996,a23998,a24000,a24002,a24004,a24006,a24008,a24010,a24012,a24014,
a24016,a24018,a24020,a24022,a24024,a24026,a24028,a24030,a24032,a24034,a24036,a24038,a24040,a24042,a24044,
a24046,a24048,a24050,a24052,a24054,a24058,a24060,a24062,a24064,a24066,a24068,a24070,a24072,a24074,a24076,
a24078,a24080,a24082,a24084,a24086,a24088,a24090,a24092,a24094,a24096,a24098,a24100,a24102,a24104,a24106,
a24108,a24110,a24112,a24114,a24116,a24118,a24120,a24122,a24124,a24126,a24128,a24130,a24132,a24134,a24136,
a24138,a24140,a24142,a24144,a24146,a24148,a24150,a24152,a24154,a24156,a24158,a24160,a24162,a24164,a24166,
a24168,a24170,a24172,a24174,a24176,a24178,a24180,a24182,a24184,a24186,a24190,a24192,a24194,a24196,a24198,
a24200,a24202,a24204,a24206,a24208,a24210,a24212,a24214,a24216,a24218,a24220,a24222,a24224,a24226,a24228,
a24230,a24232,a24234,a24236,a24238,a24240,a24242,a24244,a24246,a24248,a24250,a24252,a24254,a24256,a24258,
a24260,a24262,a24264,a24266,a24268,a24270,a24272,a24274,a24276,a24278,a24280,a24282,a24284,a24286,a24288,
a24290,a24292,a24294,a24296,a24298,a24300,a24302,a24304,a24306,a24308,a24310,a24312,a24314,a24316,a24318,
a24320,a24324,a24326,a24328,a24330,a24332,a24334,a24336,a24338,a24340,a24342,a24344,a24346,a24348,a24350,
a24352,a24354,a24356,a24358,a24360,a24362,a24364,a24366,a24368,a24370,a24372,a24374,a24376,a24378,a24380,
a24382,a24384,a24386,a24388,a24390,a24392,a24394,a24396,a24398,a24400,a24402,a24404,a24406,a24408,a24410,
a24412,a24414,a24416,a24418,a24420,a24422,a24424,a24426,a24428,a24430,a24432,a24434,a24436,a24438,a24440,
a24442,a24444,a24446,a24448,a24452,a24454,a24456,a24458,a24460,a24462,a24464,a24466,a24468,a24470,a24472,
a24474,a24476,a24478,a24480,a24482,a24484,a24486,a24488,a24490,a24492,a24494,a24496,a24498,a24500,a24502,
a24504,a24506,a24508,a24510,a24512,a24514,a24516,a24518,a24520,a24522,a24524,a24526,a24528,a24530,a24532,
a24534,a24536,a24538,a24540,a24542,a24544,a24546,a24548,a24550,a24552,a24554,a24556,a24558,a24560,a24562,
a24564,a24566,a24568,a24570,a24572,a24574,a24576,a24578,a24580,a24584,a24586,a24588,a24590,a24592,a24594,
a24596,a24598,a24600,a24602,a24604,a24606,a24608,a24610,a24612,a24614,a24616,a24618,a24620,a24622,a24624,
a24626,a24628,a24630,a24632,a24634,a24636,a24638,a24640,a24642,a24644,a24646,a24648,a24650,a24652,a24654,
a24656,a24658,a24660,a24662,a24664,a24666,a24668,a24670,a24672,a24674,a24676,a24678,a24680,a24682,a24684,
a24686,a24688,a24690,a24692,a24694,a24696,a24698,a24700,a24702,a24704,a24706,a24708,a24710,a24712,a24716,
a24718,a24720,a24722,a24724,a24726,a24728,a24730,a24732,a24734,a24736,a24738,a24740,a24742,a24744,a24746,
a24748,a24750,a24752,a24754,a24756,a24758,a24760,a24762,a24764,a24766,a24768,a24770,a24772,a24774,a24776,
a24778,a24780,a24782,a24784,a24786,a24788,a24790,a24792,a24794,a24796,a24798,a24800,a24802,a24804,a24806,
a24808,a24810,a24812,a24814,a24816,a24818,a24820,a24822,a24824,a24826,a24828,a24830,a24832,a24834,a24836,
a24838,a24840,a24842,a24844,a24848,a24850,a24852,a24854,a24856,a24858,a24860,a24862,a24864,a24866,a24868,
a24870,a24872,a24874,a24876,a24878,a24880,a24882,a24884,a24886,a24888,a24890,a24892,a24894,a24896,a24898,
a24900,a24902,a24904,a24906,a24908,a24910,a24912,a24914,a24916,a24918,a24920,a24922,a24924,a24926,a24928,
a24930,a24932,a24934,a24936,a24938,a24940,a24942,a24944,a24946,a24948,a24950,a24952,a24954,a24956,a24958,
a24960,a24962,a24964,a24966,a24968,a24970,a24972,a24976,a24978,a24980,a24982,a24984,a24986,a24988,a24990,
a24992,a24994,a24996,a24998,a25000,a25002,a25004,a25006,a25008,a25010,a25012,a25014,a25016,a25018,a25020,
a25022,a25024,a25026,a25028,a25030,a25032,a25034,a25036,a25038,a25040,a25042,a25044,a25046,a25048,a25050,
a25052,a25054,a25056,a25058,a25060,a25062,a25064,a25066,a25068,a25070,a25072,a25074,a25076,a25078,a25080,
a25082,a25084,a25086,a25088,a25090,a25092,a25094,a25096,a25098,a25100,a25102,a25104,a25108,a25110,a25112,
a25114,a25116,a25118,a25120,a25122,a25124,a25126,a25128,a25130,a25132,a25134,a25136,a25138,a25140,a25142,
a25144,a25146,a25148,a25150,a25152,a25154,a25156,a25158,a25160,a25162,a25164,a25166,a25168,a25170,a25172,
a25174,a25176,a25178,a25180,a25182,a25184,a25186,a25188,a25190,a25192,a25194,a25196,a25198,a25200,a25202,
a25204,a25206,a25208,a25210,a25212,a25214,a25216,a25218,a25220,a25222,a25224,a25226,a25228,a25230,a25232,
a25234,a25238,a25240,a25244,a25246,a25248,a25250,a25252,a25254,a25256,a25258,a25260,a25262,a25264,a25266,
a25268,a25270,a25272,a25274,a25276,a25278,a25280,a25282,a25284,a25286,a25288,a25290,a25292,a25294,a25296,
a25298,a25300,a25302,a25304,a25306,a25308,a25310,a25312,a25314,a25316,a25318,a25320,a25322,a25324,a25326,
a25328,a25330,a25332,a25334,a25336,a25338,a25340,a25342,a25344,a25346,a25348,a25350,a25352,a25354,a25356,
a25358,a25360,a25362,a25364,a25366,a25368,a25370,a25372,a25374,a25376,a25378,a25380,a25382,a25384,a25386,
a25388,a25390,a25392,a25394,a25396,a25398,a25400,a25402,a25404,a25406,a25408,a25410,a25412,a25414,a25416,
a25418,a25420,a25422,a25424,a25426,a25428,a25430,a25432,a25434,a25436,a25438,a25440,a25442,a25444,a25446,
a25448,a25450,a25452,a25454,a25456,a25458,a25460,a25462,a25464,a25466,a25468,a25470,a25472,a25474,a25476,
a25478,a25480,a25482,a25484,a25486,a25488,a25490,a25492,a25494,a25496,a25498,a25500,a25502,a25504,a25506,
a25508,a25510,a25512,a25514,a25516,a25518,a25520,a25522,a25524,a25526,a25528,a25530,a25532,a25536,a25538,
a25540,a25542,a25544,a25546,a25548,a25550,a25552,a25554,a25556,a25558,a25560,a25562,a25564,a25566,a25568,
a25570,a25572,a25574,a25576,a25580,a25582,a25584,a25586,a25588,a25590,a25592,a25594,a25596,a25598,a25600,
a25602,a25604,a25606,a25608,a25610,a25612,a25614,a25616,a25618,a25620,a25622,a25624,a25626,a25630,a25632,
a25634,a25636,a25638,a25640,a25642,a25644,a25646,a25648,a25650,a25652,a25654,a25656,a25658,a25660,a25662,
a25664,a25666,a25668,a25670,a25674,a25676,a25678,a25680,a25682,a25684,a25686,a25688,a25690,a25692,a25694,
a25696,a25698,a25700,a25702,a25704,a25706,a25708,a25710,a25712,a25714,a25716,a25718,a25720,a25722,a25724,
a25726,a25728,a25730,a25732,a25734,a25736,a25738,a25740,a25742,a25744,a25746,a25748,a25750,a25752,a25754,
a25756,a25758,a25760,a25762,a25764,a25766,a25768,a25770,a25772,a25774,a25776,a25778,a25780,a25782,a25784,
a25786,a25788,a25790,a25792,a25794,a25796,a25798,a25800,a25802,a25804,a25806,a25808,a25810,a25812,a25814,
a25816,a25818,a25820,a25822,a25824,a25826,a25828,a25830,a25832,a25834,a25836,a25840,a25842,a25844,a25848,
a25854,a25856,a25858,a25860,a25862,a25864,a25866,a25868,a25870,a25872,a25874,a25876,a25878,a25880,a25882,
a25884,a25886,a25888,a25890,a25892,a25894,a25896,a25898,a25900,a25902,a25904,a25906,a25908,a25910,a25912,
a25914,a25916,a25918,a25920,a25922,a25924,a25926,a25928,a25930,a25932,a25934,a25936,a25938,a25940,a25942,
a25944,a25946,a25948,a25950,a25952,a25954,a25956,a25958,a25960,a25962,a25964,a25966,a25968,a25970,a25972,
a25974,a25976,a25978,a25980,a25982,a25984,a25986,a25988,a25990,a25992,a25994,a25996,a25998,a26000,a26002,
a26004,a26006,a26008,a26010,a26012,a26014,a26016,a26018,a26020,a26022,a26024,a26026,a26028,a26030,a26032,
a26034,a26036,a26038,a26040,a26042,a26044,a26046,a26048,a26050,a26052,a26054,a26056,a26058,a26060,a26062,
a26064,a26066,a26068,a26070,a26072,a26074,a26076,a26078,a26080,a26082,a26084,a26086,a26088,a26090,a26092,
a26094,a26096,a26098,a26100,a26102,a26104,a26106,a26108,a26110,a26112,a26114,a26116,a26118,a26120,a26122,
a26124,a26126,a26128,a26130,a26132,a26134,a26136,a26138,a26140,a26142,a26144,a26146,a26148,a26150,a26152,
a26154,a26156,a26158,a26160,a26162,a26164,a26166,a26168,a26170,a26172,a26174,a26176,a26178,a26180,a26182,
a26184,a26186,a26188,a26190,a26192,a26194,a26196,a26198,a26200,a26202,a26204,a26206,a26208,a26210,a26212,
a26214,a26216,a26218,a26220,a26222,a26224,a26226,a26228,a26230,a26232,a26234,a26236,a26238,a26240,a26242,
a26244,a26246,a26248,a26250,a26252,a26254,a26256,a26258,a26260,a26262,a26264,a26266,a26268,a26270,a26272,
a26274,a26276,a26278,a26280,a26282,a26284,a26286,a26288,a26290,a26292,a26294,a26296,a26298,a26300,a26302,
a26304,a26306,a26308,a26310,a26312,a26314,a26316,a26318,a26320,a26322,a26324,a26326,a26328,a26330,a26332,
a26334,a26336,a26338,a26340,a26342,a26344,a26346,a26348,a26350,a26352,a26354,a26356,a26358,a26360,a26362,
a26364,a26366,a26368,a26370,a26372,a26374,a26376,a26378,a26380,a26382,a26384,a26386,a26388,a26390,a26392,
a26394,a26396,a26398,a26400,a26402,a26404,a26406,a26408,a26410,a26412,a26414,a26416,a26418,a26420,a26422,
a26424,a26426,a26428,a26430,a26432,a26434,a26436,a26438,a26440,a26442,a26444,a26446,a26448,a26450,a26452,
a26454,a26456,a26458,a26460,a26462,a26464,a26466,a26468,a26470,a26472,a26474,a26476,a26478,a26480,a26482,
a26484,a26486,a26488,a26490,a26492,a26494,a26496,a26498,a26500,a26502,a26504,a26506,a26508,a26510,a26512,
a26514,a26516,a26518,a26520,a26522,a26524,a26526,a26528,a26530,a26532,a26534,a26536,a26538,a26540,a26542,
a26544,a26546,a26548,a26550,a26552,a26554,a26556,a26558,a26560,a26562,a26564,a26566,a26568,a26570,a26572,
a26574,a26576,a26578,a26580,a26582,a26584,a26586,a26588,a26590,a26592,a26594,a26596,a26598,a26600,a26602,
a26604,a26606,a26608,a26610,a26612,a26614,a26616,a26618,a26620,a26622,a26624,a26626,a26628,a26630,a26632,
a26634,a26636,a26638,a26640,a26642,a26644,a26646,a26648,a26650,a26652,a26654,a26656,a26658,a26660,a26662,
a26664,a26666,a26668,a26670,a26672,a26674,a26676,a26678,a26680,a26682,a26684,a26686,a26688,a26690,a26692,
a26694,a26696,a26698,a26700,a26702,a26704,a26706,a26708,a26710,a26712,a26714,a26716,a26718,a26720,a26722,
a26724,a26726,a26728,a26730,a26732,a26734,a26736,a26738,a26740,a26742,a26744,a26746,a26748,a26750,a26752,
a26754,a26756,a26758,a26760,a26762,a26764,a26766,a26768,a26770,a26772,a26774,a26776,a26778,a26780,a26782,
a26784,a26786,a26788,a26790,a26792,a26794,a26796,a26798,a26800,a26802,a26804,a26806,a26808,a26810,a26812,
a26814,a26816,a26818,a26820,a26822,a26824,a26826,a26828,a26830,a26832,a26834,a26836,a26838,a26840,a26842,
a26844,a26846,a26848,a26850,a26852,a26854,a26856,a26858,a26860,a26862,a26864,a26866,a26868,a26870,a26872,
a26874,a26876,a26878,a26880,a26882,a26884,a26886,a26888,a26890,a26892,a26894,a26896,a26898,a26900,a26902,
a26904,a26906,a26908,a26910,a26912,a26914,a26916,a26918,a26920,a26922,a26924,a26926,a26928,a26930,a26932,
a26934,a26936,a26938,a26940,a26942,a26944,a26946,a26948,a26950,a26952,a26954,a26956,a26958,a26960,a26962,
a26964,a26966,a26968,a26970,a26972,a26974,a26976,a26978,a26980,a26982,a26984,a26986,a26988,a26990,a26992,
a26994,a26996,a26998,a27000,a27002,a27004,a27006,a27008,a27010,a27012,a27014,a27016,a27018,a27020,a27022,
a27024,a27026,a27028,a27030,a27032,a27034,a27036,a27038,a27040,a27042,a27044,a27046,a27048,a27050,a27052,
a27054,a27056,a27058,a27060,a27062,a27064,a27066,a27068,a27070,a27072,a27074,a27076,a27078,a27080,a27082,
a27084,a27086,a27088,a27090,a27092,a27094,a27096,a27098,a27100,a27102,a27104,a27106,a27108,a27110,a27112,
a27114,a27116,a27118,a27120,a27122,a27124,a27126,a27128,a27130,a27132,a27134,a27136,a27138,a27140,a27142,
a27144,a27146,a27148,a27150,a27152,a27154,a27156,a27158,a27160,a27162,a27164,a27166,a27168,a27170,a27172,
a27174,a27176,a27178,a27180,a27182,a27184,a27186,a27188,a27190,a27192,a27194,a27196,a27198,a27200,a27202,
a27204,a27206,a27208,a27210,a27212,a27214,a27216,a27218,a27220,a27222,a27224,a27226,a27228,a27230,a27232,
a27234,a27236,a27238,a27240,a27242,a27244,a27246,a27248,a27250,a27252,a27254,a27256,a27258,a27260,a27262,
a27264,a27266,a27268,a27270,a27272,a27274,a27276,a27278,a27280,a27282,a27284,a27286,a27288,a27290,a27292,
a27294,a27296,a27298,a27300,a27302,a27304,a27306,a27308,a27310,a27312,a27314,a27316,a27318,a27320,a27322,
a27324,a27326,a27328,a27330,a27332,a27334,a27336,a27338,a27340,a27342,a27344,a27346,a27348,a27350,a27352,
a27354,a27356,a27358,a27360,a27362,a27364,a27366,a27368,a27370,a27372,a27374,a27376,a27378,a27380,a27382,
a27384,a27386,a27388,a27390,a27392,a27394,a27396,a27398,a27400,a27402,a27404,a27406,a27408,a27410,a27412,
a27414,a27416,a27418,a27420,a27422,a27424,a27426,a27428,a27430,a27432,a27434,a27436,a27438,a27440,a27442,
a27444,a27446,a27448,a27450,a27452,a27454,a27456,a27458,a27460,a27462,a27464,a27466,a27468,a27470,a27472,
a27474,a27476,a27478,a27480,a27482,a27484,a27486,a27488,a27490,a27492,a27494,a27496,a27498,a27500,a27502,
a27504,a27506,a27508,a27510,a27512,a27514,a27516,a27518,a27520,a27522,a27524,a27526,a27528,a27530,a27532,
a27534,a27536,a27538,a27540,a27542,a27544,a27546,a27548,a27550,a27552,a27554,a27556,a27558,a27560,a27562,
a27564,a27566,a27568,a27570,a27572,a27574,a27576,a27578,a27580,a27582,a27584,a27586,a27588,a27590,a27592,
a27594,a27596,a27598,a27600,a27602,a27604,a27606,a27608,a27610,a27612,a27614,a27616,a27618,a27620,a27622,
a27624,a27626,a27628,a27630,a27632,a27634,a27636,a27638,a27640,a27642,a27644,a27646,a27648,a27650,a27652,
a27654,a27656,a27658,a27660,a27662,a27664,a27666,a27668,a27670,a27672,a27674,a27676,a27678,a27680,a27682,
a27684,a27686,a27688,a27690,a27692,a27694,a27696,a27698,a27700,a27702,a27704,a27706,a27708,a27710,a27712,
a27714,a27716,a27718,a27720,a27722,a27724,a27726,a27728,a27730,a27732,a27734,a27736,a27738,a27740,a27742,
a27744,a27746,a27748,a27750,a27752,a27754,a27756,a27758,a27760,a27762,a27764,a27766,a27768,a27770,a27772,
a27774,a27776,a27778,a27780,a27782,a27784,a27786,a27788,a27790,a27792,a27794,a27796,a27798,a27800,a27802,
a27804,a27806,a27808,a27810,a27812,a27814,a27816,a27818,a27820,a27822,a27824,a27826,a27828,a27830,a27832,
a27834,a27836,a27838,a27840,a27842,a27844,a27846,a27848,a27850,a27852,a27854,a27856,a27858,a27860,a27862,
a27864,a27866,a27868,a27870,a27872,a27874,a27876,a27878,a27880,a27882,a27884,a27886,a27888,a27890,a27892,
a27894,a27896,a27898,a27900,a27902,a27904,a27906,a27908,a27910,a27912,a27914,a27916,a27918,a27920,a27922,
a27924,a27926,a27928,a27930,a27932,a27934,a27936,a27938,a27940,a27942,a27944,a27946,a27948,a27950,a27952,
a27954,a27956,a27958,a27960,a27962,a27964,a27966,a27968,a27970,a27972,a27974,a27976,a27978,a27980,a27982,
a27984,a27986,a27988,a27990,a27992,a27994,a27996,a27998,a28000,a28002,a28004,a28006,a28008,a28010,a28012,
a28014,a28016,a28018,a28020,a28022,a28024,a28026,a28028,a28030,a28032,a28034,a28036,a28038,a28040,a28042,
a28044,a28046,a28048,a28050,a28052,a28054,a28056,a28058,a28060,a28062,a28064,a28066,a28068,a28070,a28072,
a28074,a28076,a28078,a28080,a28082,a28084,a28086,a28088,a28090,a28092,a28094,a28096,a28098,a28100,a28102,
a28104,a28106,a28108,a28110,a28112,a28114,a28116,a28118,a28120,a28122,a28124,a28126,a28128,a28130,a28132,
a28134,a28136,a28138,a28140,a28142,a28144,a28146,a28148,a28150,a28152,a28154,a28156,a28158,a28160,a28162,
a28164,a28166,a28168,a28170,a28172,a28174,a28176,a28178,a28180,a28182,a28184,a28186,a28190,a28192,a28196,
a28198,a28200,a28202,a28204,a28206,a28208,a28210,a28212,a28214,a28216,a28218,a28220,a28222,a28224,a28226,
a28228,a28230,a28232,a28234,a28238,a28240,a28242,a28244,a28246,a28248,a28250,a28252,a28254,a28256,a28258,
a28260,a28262,a28264,a28266,a28268,a28270,a28272,a28274,a28276,a28278,a28280,a28282,a28284,a28286,a28288,
a28290,a28292,a28294,a28296,a28298,a28300,a28302,a28304,a28306,a28308,a28310,a28312,a28314,a28316,a28318,
a28320,a28322,a28324,a28326,a28328,a28330,a28332,a28334,a28336,a28338,a28340,a28342,a28344,a28346,a28348,
a28350,a28352,a28354,a28356,a28358,a28360,a28362,a28364,a28366,a28368,a28370,a28372,a28374,a28376,a28378,
a28380,a28382,a28384,a28386,a28388,a28390,a28392,a28394,a28396,a28398,a28400,a28402,a28404,a28406,a28408,
a28410,a28412,a28414,a28416,a28418,a28420,a28422,a28424,a28426,a28428,a28430,a28432,a28434,a28436,a28438,
a28440,a28442,a28444,a28446,a28450,a28452,a28454,a28456,a28458,a28460,a28462,a28464,a28466,a28468,a28470,
a28472,a28474,a28476,a28478,a28480,a28482,a28484,a28486,a28488,a28490,a28492,a28494,a28496,a28498,a28500,
a28502,a28504,a28506,a28508,a28510,a28512,a28514,a28516,a28518,a28520,a28522,a28524,a28526,a28528,a28530,
a28532,a28534,a28536,a28538,a28540,a28542,a28544,a28546,a28548,a28550,a28552,a28554,a28556,a28558,a28560,
a28562,a28564,a28566,a28568,a28570,a28572,a28574,a28576,a28578,a28580,a28582,a28584,a28586,a28588,a28590,
a28592,a28594,a28596,a28598,a28600,a28602,a28604,a28606,a28608,a28610,a28612,a28614,a28616,a28618,a28620,
a28622,a28624,a28626,a28628,a28630,a28632,a28634,a28636,a28638,a28640,a28642,a28644,a28646,a28648,a28650,
a28652,a28654,a28656,a28658,a28660,a28662,a28664,a28666,a28668,a28670,a28672,a28674,a28676,a28678,a28680,
a28682,a28684,a28686,a28688,a28690,a28692,a28694,a28696,a28698,a28700,a28702,a28704,a28708,a28710,a28712,
a28714,a28716,a28718,a28720,a28722,a28724,a28726,a28728,a28730,a28732,a28734,a28736,a28738,a28740,a28742,
a28744,a28746,a28748,a28750,a28752,a28754,a28756,a28758,a28760,a28762,a28764,a28766,a28768,a28770,a28772,
a28774,a28776,a28778,a28780,a28782,a28784,a28786,a28788,a28790,a28792,a28794,a28796,a28798,a28800,a28802,
a28804,a28806,a28808,a28810,a28812,a28814,a28816,a28818,a28820,a28822,a28824,a28826,a28828,a28830,a28832,
a28834,a28836,a28838,a28840,a28842,a28844,a28846,a28848,a28850,a28852,a28854,a28856,a28858,a28860,a28862,
a28864,a28866,a28868,a28870,a28872,a28874,a28876,a28878,a28880,a28882,a28884,a28886,a28888,a28890,a28892,
a28894,a28896,a28898,a28900,a28902,a28904,a28906,a28908,a28910,a28912,a28914,a28916,a28918,a28920,a28922,
a28924,a28926,a28928,a28930,a28932,a28934,a28936,a28938,a28940,a28942,a28946,a28948,a28950,a28952,a28954,
a28956,a28958,a28960,a28962,a28964,a28966,a28968,a28970,a28972,a28974,a28976,a28978,a28980,a28982,a28984,
a28986,a28988,a28990,a28992,a28994,a28996,a28998,a29000,a29002,a29004,a29006,a29008,a29010,a29012,a29014,
a29016,a29018,a29020,a29022,a29024,a29026,a29028,a29030,a29032,a29034,a29036,a29038,a29040,a29042,a29044,
a29046,a29048,a29050,a29052,a29054,a29056,a29058,a29060,a29062,a29064,a29066,a29068,a29070,a29072,a29074,
a29076,a29078,a29080,a29082,a29084,a29086,a29088,a29090,a29092,a29094,a29096,a29098,a29100,a29102,a29104,
a29106,a29108,a29110,a29112,a29114,a29116,a29118,a29120,a29122,a29124,a29126,a29128,a29130,a29132,a29134,
a29136,a29138,a29140,a29142,a29144,a29146,a29148,a29150,a29152,a29154,a29156,a29158,a29160,a29162,a29164,
a29166,a29168,a29170,a29172,a29174,a29176,a29178,a29180,a29182,a29184,a29186,a29188,a29190,a29192,a29194,
a29196,a29198,a29200,a29202,a29204,a29206,a29208,a29212,a29214,a29216,a29218,a29220,a29222,a29224,a29226,
a29228,a29230,a29232,a29234,a29236,a29238,a29240,a29242,a29244,a29246,a29248,a29250,a29252,a29254,a29256,
a29258,a29260,a29262,a29264,a29266,a29268,a29270,a29272,a29274,a29276,a29278,a29280,a29282,a29284,a29286,
a29288,a29290,a29292,a29294,a29296,a29298,a29300,a29302,a29304,a29306,a29308,a29310,a29312,a29314,a29316,
a29318,a29320,a29322,a29324,a29326,a29328,a29330,a29332,a29334,a29336,a29338,a29340,a29342,a29344,a29346,
a29348,a29350,a29352,a29354,a29356,a29358,a29360,a29362,a29364,a29366,a29368,a29370,a29372,a29374,a29376,
a29378,a29380,a29382,a29384,a29386,a29388,a29390,a29392,a29394,a29396,a29398,a29400,a29402,a29404,a29406,
a29408,a29410,a29412,a29414,a29416,a29418,a29420,a29422,a29424,a29426,a29428,a29430,a29432,a29434,a29436,
a29438,a29440,a29442,a29444,a29446,a29448,a29450,a29452,a29454,a29456,a29458,a29460,a29464,a29466,a29468,
a29470,a29472,a29474,a29476,a29478,a29480,a29482,a29484,a29486,a29488,a29490,a29492,a29494,a29496,a29498,
a29500,a29502,a29504,a29506,a29510,a29512,a29514,a29516,a29518,a29520,a29522,a29524,a29526,a29528,a29530,
a29532,a29534,a29536,a29538,a29540,a29542,a29544,a29546,a29550,a29552,a29554,a29556,a29558,a29560,a29562,
a29564,a29566,a29568,a29570,a29572,a29574,a29576,a29578,a29580,a29582,a29584,a29586,a29588,a29590,a29592,
a29594,a29596,a29598,a29600,a29602,a29604,a29606,a29608,a29610,a29612,a29614,a29616,a29618,a29620,a29622,
a29624,a29626,a29628,a29630,a29632,a29634,a29636,a29638,a29640,a29644,a29646,a29648,a29650,a29652,a29654,
a29656,a29658,a29660,a29662,a29664,a29666,a29668,a29670,a29672,a29674,a29676,a29678,a29680,a29682,a29684,
a29686,a29688,a29690,a29692,a29694,a29696,a29698,a29700,a29702,a29704,a29706,a29708,a29710,a29712,a29714,
a29716,a29718,a29720,a29724,a29726,a29730,a29732,a29734,a29736,a29738,a29740,a29742,a29744,a29746,a29748,
a29750,a29752,a29754,a29756,a29758,a29760,a29762,a29764,a29766,a29768,a29770,a29772,a29774,a29776,a29778,
a29780,a29782,a29784,a29786,a29790,a29792,a29796,a29798,a29800,a29802,a29804,a29806,a29808,a29810,a29812,
a29814,a29816,a29818,a29820,a29822,a29824,a29826,a29828,a29830,a29832,a29834,a29836,a29838,a29840,a29842,
a29844,a29846,a29848,a29850,a29852,a29856,a29858,a29862,a29864,a29866,a29868,a29870,a29872,a29874,a29876,
a29878,a29880,a29882,a29884,a29886,a29888,a29890,a29892,a29894,a29896,a29898,a29900,a29902,a29904,a29906,
a29908,a29910,a29912,a29914,a29916,a29918,a29922,a29924,a29928,a29930,a29932,a29934,a29936,a29938,a29940,
a29942,a29944,a29946,a29948,a29950,a29952,a29954,a29956,a29958,a29960,a29962,a29964,a29966,a29968,a29970,
a29972,a29974,a29976,a29978,a29980,a29982,a29984,a29988,a29990,a29992,a29994,a29996,a29998,a30000,a30002,
a30004,a30006,a30008,a30010,a30012,a30014,a30016,a30018,a30020,a30022,a30024,a30026,a30028,a30030,a30032,
a30034,a30036,a30038,a30040,a30042,a30044,a30046,a30048,a30050,a30052,a30054,a30056,a30058,a30060,a30062,
a30064,a30066,a30068,a30070,a30072,a30074,a30076,a30078,a30080,a30082,a30084,a30086,a30088,a30090,a30092,
a30094,a30096,a30098,a30100,a30102,a30104,a30106,a30108,a30110,a30112,a30114,a30116,a30118,a30120,a30122,
a30124,a30126,a30128,a30130,a30132,a30134,a30136,a30138,a30140,a30142,a30144,a30146,a30148,a30150,a30152,
a30154,a30156,a30158,a30160,a30162,a30164,a30166,a30168,a30170,a30172,a30174,a30176,a30178,a30180,a30182,
a30184,a30186,a30188,a30190,a30192,a30194,a30196,a30198,a30200,a30202,a30204,a30206,a30208,a30210,a30212,
a30214,a30216,a30218,a30220,a30222,a30224,a30226,a30228,a30230,a30232,a30234,a30236,a30238,a30240,a30242,
a30244,a30246,a30248,a30250,a30252,a30254,a30256,a30258,a30260,a30262,a30264,a30266,a30268,a30270,a30272,
a30274,a30276,a30278,a30280,a30282,a30284,a30286,a30288,a30290,a30292,a30294,a30296,a30298,a30300,a30302,
a30304,a30306,a30308,a30310,a30312,a30314,a30316,a30318,a30320,a30322,a30324,a30326,a30328,a30330,a30332,
a30334,a30336,a30338,a30340,a30342,a30344,a30346,a30348,a30350,a30352,a30354,a30356,a30358,a30360,a30362,
a30364,a30366,a30368,a30370,a30372,a30374,a30376,a30378,a30380,a30382,a30384,a30386,a30388,a30390,a30392,
a30394,a30396,a30398,a30400,a30402,a30404,a30406,a30408,a30410,a30412,a30414,a30416,a30418,a30420,a30422,
a30424,a30426,a30428,a30430,a30432,a30434,a30436,a30438,a30440,a30442,a30444,a30446,a30448,a30450,a30452,
a30454,a30456,a30458,a30460,a30462,a30464,a30466,a30468,a30470,a30472,a30474,a30476,a30478,a30480,a30482,
a30484,a30486,a30488,a30490,a30492,a30494,a30496,a30498,a30500,a30502,a30504,a30506,a30508,a30510,a30512,
a30514,a30516,a30518,a30520,a30522,a30524,a30526,a30528,a30530,a30532,a30534,a30536,a30538,a30540,a30542,
a30544,a30546,a30548,a30550,a30552,a30554,a30556,a30558,a30560,a30562,a30564,a30566,a30568,a30570,a30572,
a30574,a30576,a30578,a30580,a30582,a30584,a30586,a30588,a30590,a30592,a30594,a30596,a30598,a30600,a30602,
a30604,a30606,a30608,a30610,a30612,a30614,a30616,a30618,a30620,a30622,a30624,a30626,a30628,a30630,a30632,
a30634,a30636,a30638,a30640,a30642,a30644,a30646,a30648,a30650,a30652,a30654,a30656,a30658,a30660,a30662,
a30664,a30666,a30668,a30670,a30672,a30674,a30676,a30678,a30680,a30682,a30684,a30686,a30688,a30690,a30692,
a30694,a30696,a30698,a30700,a30702,a30704,a30706,a30708,a30710,a30712,a30714,a30716,a30718,a30720,a30722,
a30724,a30726,a30728,a30730,a30732,a30734,a30736,a30738,a30740,a30742,a30744,a30746,a30748,a30750,a30752,
a30754,a30756,a30758,a30760,a30762,a30764,a30766,a30768,a30770,a30772,a30774,a30776,a30778,a30780,a30782,
a30784,a30786,a30788,a30790,a30792,a30794,a30796,a30798,a30800,a30802,a30804,a30806,a30808,a30810,a30812,
a30814,a30816,a30818,a30820,a30822,a30824,a30826,a30828,a30830,a30832,a30834,a30836,a30838,a30840,a30842,
a30844,a30846,a30848,a30850,a30852,a30854,a30856,a30858,a30860,a30862,a30864,a30866,a30868,a30870,a30872,
a30874,a30876,a30878,a30880,a30882,a30884,a30886,a30888,a30890,a30892,a30894,a30896,a30898,a30900,a30902,
a30904,a30906,a30908,a30910,a30912,a30914,a30916,a30918,a30920,a30922,a30924,a30926,a30928,a30930,a30932,
a30934,a30936,a30938,a30940,a30942,a30944,a30946,a30948,a30950,a30952,a30954,a30956,a30958,a30960,a30962,
a30964,a30966,a30968,a30970,a30972,a30974,a30976,a30978,a30980,a30982,a30984,a30986,a30988,a30990,a30992,
a30994,a30996,a30998,a31000,a31002,a31004,a31006,a31008,a31010,a31012,a31014,a31016,a31022,a31024,a31026,
a31028,a31030,a31032,a31034,a31036,a31038,a31044,a31046,a31048,a31050,a31052,a31054,a31056,a31058,a31060,
a31062,a31064,a31066,a31068,a31070,a31072,a31074,a31076,a31078,a31080,a31082,a31084,a31086,a31090,a31092,
a31094,a31096,a31098,a31100,a31102,a31104,a31106,a31108,a31110,a31112,a31114,a31116,a31118,a31120,a31122,
a31124,a31126,a31128,a31130,a31132,a31134,a31136,a31138,a31140,a31142,a31144,a31146,a31148,a31150,a31152,
a31154,a31156,a31158,a31162,a31164,a31166,a31168,a31170,a31172,a31174,a31176,a31178,a31180,a31184,a31186,
a31188,a31190,a31192,a31194,a31196,a31198,a31200,a31202,a31204,a31206,a31210,a31212,a31214,a31216,a31218,
a31220,a31222,a31224,a31226,a31228,a31230,a31232,a31234,a31236,a31238,a31240,a31242,a31244,a31246,a31248,
a31250,a31252,a31254,a31256,a31258,a31260,a31262,a31264,a31266,a31268,a31270,a31272,a31274,a31276,a31278,
a31280,a31282,a31284,a31286,a31288,a31290,a31292,a31294,a31296,a31298,a31300,a31302,a31304,a31306,a31308,
a31310,a31312,a31314,a31316,a31318,a31320,a31322,a31324,a31326,a31328,a31330,a31332,a31334,a31336,a31338,
a31340,a31342,a31344,a31346,a31348,a31350,a31352,a31354,a31356,a31358,a31360,a31362,a31364,a31366,a31368,
a31370,a31372,a31374,a31376,a31378,a31380,a31382,a31384,a31386,a31388,a31390,a31392,a31394,a31396,a31398,
a31400,a31402,a31404,a31406,a31408,a31410,a31412,a31414,a31416,a31418,a31420,a31422,a31424,a31426,a31428,
a31430,a31432,a31434,a31436,a31438,a31440,a31442,a31444,a31446,a31448,a31450,a31452,a31454,a31456,a31458,
a31460,a31462,a31464,a31466,a31468,a31470,a31472,a31474,a31476,a31478,a31480,a31482,a31484,a31486,a31488,
a31490,a31492,a31494,a31496,a31498,a31500,a31502,a31504,a31506,a31508,a31510,a31512,a31514,a31516,a31518,
a31520,a31522,a31524,a31526,a31528,a31530,a31532,a31534,a31536,a31538,a31540,a31542,a31544,a31546,a31548,
a31550,a31552,a31554,a31556,a31558,a31560,a31562,a31564,a31566,a31568,a31570,a31572,a31574,a31576,a31578,
a31580,a31582,a31584,a31586,a31588,a31590,a31592,a31594,a31596,a31598,a31600,a31602,a31604,a31606,a31608,
a31610,a31612,a31614,a31616,a31618,a31620,a31622,a31624,a31626,a31628,a31630,a31632,a31634,a31636,a31638,
a31640,a31642,a31644,a31646,a31648,a31650,a31652,a31654,a31656,a31658,a31660,a31662,a31664,a31666,a31668,
a31670,a31672,a31674,a31676,a31678,a31680,a31682,a31684,a31686,a31688,a31690,a31692,a31694,a31696,a31698,
a31700,a31702,a31704,a31706,a31708,a31710,a31712,a31714,a31716,a31718,a31720,a31722,a31724,a31726,a31728,
a31730,a31732,a31734,a31736,a31738,a31740,a31742,a31744,a31746,a31748,a31750,a31752,a31754,a31756,a31758,
a31760,a31762,a31764,a31766,a31768,a31770,a31772,a31774,a31776,a31778,a31780,a31782,a31784,a31786,a31788,
a31790,a31792,a31794,a31796,a31798,a31800,a31802,a31804,a31806,a31808,a31810,a31812,a31814,a31816,a31818,
a31820,a31822,a31824,a31826,a31828,a31830,a31832,a31834,a31836,a31838,a31840,a31842,a31844,a31846,a31848,
a31850,a31852,a31854,a31856,a31858,a31860,a31862,a31864,a31866,a31868,a31870,a31872,a31874,a31876,a31878,
a31880,a31882,a31884,a31886,a31888,a31890,a31892,a31894,a31896,a31898,a31900,a31902,a31904,a31906,a31908,
a31910,a31912,a31914,a31916,a31918,a31920,a31922,a31924,a31926,a31928,a31930,a31932,a31934,a31936,a31938,
a31940,a31942,a31944,a31946,a31948,a31950,a31952,a31954,a31956,a31958,a31960,a31962,a31964,a31966,a31968,
a31970,a31972,a31974,a31976,a31978,a31980,a31982,a31984,a31986,a31988,a31990,a31992,a31994,a31996,a31998,
a32000,a32002,a32004,a32006,a32008,a32010,a32012,a32014,a32016,a32018,a32020,a32022,a32024,a32026,a32028,
a32030,a32032,a32034,a32036,a32038,a32040,a32042,a32044,a32046,a32048,a32050,a32052,a32054,a32056,a32058,
a32060,a32062,a32064,a32066,a32068,a32070,a32072,a32074,a32076,a32078,a32080,a32082,a32084,a32086,a32088,
a32090,a32092,a32094,a32096,a32098,a32100,a32102,a32104,a32106,a32108,a32110,a32112,a32114,a32116,a32118,
a32120,a32122,a32124,a32126,a32128,a32130,a32132,a32134,a32136,a32138,a32140,a32142,a32144,a32146,a32148,
a32150,a32152,a32154,a32156,a32158,a32160,a32162,a32164,a32166,a32168,a32170,a32172,a32174,a32176,a32178,
a32180,a32182,a32184,a32186,a32188,a32190,a32192,a32194,a32196,a32198,a32200,a32202,a32204,a32206,a32208,
a32210,a32212,a32214,a32216,a32218,a32220,a32222,a32224,a32226,a32228,a32230,a32232,a32234,a32236,a32238,
a32240,a32242,a32244,a32246,a32248,a32250,a32252,a32254,a32256,a32258,a32260,a32262,a32264,a32266,a32268,
a32270,a32272,a32274,a32276,a32278,a32280,a32282,a32284,a32286,a32288,a32290,a32292,a32294,a32296,a32298,
a32300,a32302,a32304,a32306,a32308,a32310,a32312,a32314,a32316,a32318,a32320,a32322,a32324,a32326,a32328,
a32330,a32332,a32334,a32336,a32338,a32340,a32342,a32344,a32346,a32348,a32350,a32352,a32354,a32356,a32358,
a32360,a32362,a32364,a32366,a32368,a32372,a32374,a32376,a32378,a32382,a32384,a32388,a32390,a32392,a32394,
a32396,a32398,a32400,a32402,a32404,a32406,a32408,a32410,a32412,a32414,a32416,a32418,a32420,a32422,a32424,
a32426,a32428,a32430,a32432,a32434,a32436,a32438,a32440,a32442,a32444,a32446,a32448,a32450,a32452,a32454,
a32456,a32458,a32460,a32462,a32464,a32466,a32468,a32472,a32474,a32476,a32478,a32480,a32482,a32484,a32488,
a32490,a32492,a32494,a32496,a32498,a32500,a32502,a32506,a32510,a32512,a32514,a32516,a32518,a32520,a32522,
a32524,a32526,a32528,a32530,a32532,a32534,a32536,a32540,a32542,a32544,a32546,a32548,a32550,a32552,a32554,
a32556,a32558,a32560,a32562,a32564,a32566,a32568,a32570,a32572,a32574,a32576,a32578,a32580,a32582,a32584,
a32586,a32588,a32590,a32594,a32596,a32598,a32600,a32602,a32604,a32606,a32608,a32610,a32612,a32614,a32616,
a32618,a32620,a32622,a32624,a32626,a32628,a32630,a32632,a32636,a32638,a32640,a32642,a32644,a32646,a32648,
a32650,a32652,a32654,a32656,a32658,a32660,a32662,a32664,a32666,a32668,a32670,a32672,a32674,a32676,a32678,
a32682,a32684,a32686,a32688,a32690,a32692,a32694,a32696,a32698,a32700,a32702,a32704,a32706,a32708,a32710,
a32712,a32714,a32716,a32718,a32720,a32724,a32726,a32728,a32730,a32732,a32734,a32736,a32738,a32740,a32742,
a32744,a32746,a32748,a32750,a32752,a32754,a32756,a32758,a32760,a32762,a32764,a32766,a32768,a32770,a32774,
a32776,a32778,a32780,a32782,a32784,a32786,a32788,a32790,a32792,a32794,a32796,a32798,a32800,a32802,a32804,
a32806,a32808,a32810,a32812,a32816,a32818,a32820,a32822,a32824,a32826,a32828,a32830,a32832,a32834,a32836,
a32838,a32840,a32842,a32844,a32846,a32848,a32850,a32852,a32854,a32856,a32858,a32862,a32864,a32866,a32868,
a32870,a32872,a32874,a32876,a32878,a32880,a32882,a32884,a32886,a32888,a32890,a32892,a32894,a32896,a32898,
a32900,a32902,a32904,a32906,a32910,a32912,a32914,a32916,a32918,a32920,a32922,a32924,a32926,a32928,a32930,
a32932,a32934,a32936,a32938,a32940,a32942,a32944,a32946,a32948,a32950,a32952,a32954,a32956,a32958,a32960,
a32962,a32964,a32968,a32970,a32972,a32974,a32976,a32980,a32982,a32984,a32986,a32988,a32990,a32992,a32994,
a32996,a33000,a33002,a33004,a33006,a33008,a33010,a33012,a33016,a33018,a33020,a33022,a33024,a33026,a33028,
a33030,a33034,a33036,a33038,a33040,a33042,a33044,a33048,a33050,a33052,a33054,a33056,a33058,a33060,a33062,
a33064,a33068,a33070,a33072,a33074,a33076,a33080,a33082,a33084,a33086,a33088,a33090,a33092,a33096,a33098,
a33100,a33102,a33104,a33108,a33110,a33112,a33114,a33116,a33118,a33120,a33122,a33124,a33126,a33128,a33130,
a33132,a33134,a33136,a33138,a33140,a33142,a33144,a33146,a33148,a33150,a33152,a33154,a33158,a33160,a33162,
a33164,a33166,a33168,a33170,a33172,a33174,a33176,a33178,a33180,a33182,a33184,a33186,a33188,a33190,a33192,
a33194,a33196,a33200,a33202,a33204,a33206,a33208,a33210,a33212,a33214,a33216,a33218,a33220,a33222,a33224,
a33226,a33228,a33230,a33232,a33234,a33236,a33238,a33240,a33242,a33244,a33246,a33248,a33250,a33252,a33254,
a33256,a33258,a33260,a33262,a33264,a33266,a33268,a33270,a33272,a33274,a33276,a33278,a33280,a33282,a33284,
a33286,a33288,a33290,a33292,a33294,a33296,a33298,a33300,a33302,a33304,a33306,a33308,a33310,a33312,a33314,
a33316,a33318,a33320,a33322,a33324,a33326,a33328,a33330,a33332,a33334,a33336,a33338,a33340,a33342,a33344,
a33346,a33348,a33350,a33352,a33354,a33356,a33358,a33360,a33362,a33364,a33366,a33368,a33370,a33372,a33374,
a33376,a33378,a33380,a33382,a33384,a33386,a33388,a33390,a33392,a33394,a33396,a33398,a33400,a33402,a33404,
a33406,a33408,a33410,a33412,a33414,a33416,a33418,a33420,a33422,a33424,a33426,a33428,a33432,a33434,a33436,
a33438,a33440,a33442,a33444,a33446,a33448,a33450,a33452,a33454,a33456,a33460,a33462,a33464,a33466,a33468,
a33470,a33472,a33474,a33476,a33478,a33480,a33482,a33484,a33486,a33488,a33490,a33492,a33494,a33496,a33498,
a33500,a33502,a33504,a33506,a33508,a33510,a33512,a33514,a33516,a33518,a33520,a33522,a33524,a33526,a33528,
a33530,a33532,a33534,a33536,a33538,a33540,a33542,a33544,a33546,a33548,a33550,a33552,a33554,a33556,a33558,
a33560,a33562,a33564,a33566,a33568,a33570,a33572,a33574,a33576,a33578,a33580,a33582,a33584,a33586,a33588,
a33590,a33592,a33594,a33596,a33598,a33600,a33602,a33604,a33606,a33608,a33610,a33612,a33614,a33616,a33618,
a33620,a33622,a33624,a33626,a33628,a33630,a33632,a33634,a33636,a33638,a33640,a33642,a33644,a33646,a33648,
a33650,a33652,a33654,a33656,a33658,a33660,a33662,a33664,a33666,a33668,a33670,a33672,a33674,a33676,a33678,
a33680,a33682,a33684,a33686,a33688,a33690,a33692,a33694,a33696,a33698,a33700,a33702,a33704,a33706,a33708,
a33710,a33712,a33714,a33716,a33718,a33720,a33722,a33724,a33726,a33728,a33730,a33732,a33734,a33736,a33738,
a33740,a33742,a33744,a33746,a33748,a33750,a33752,a33754,a33756,a33758,a33760,a33762,a33764,a33766,a33768,
a33770,a33772,a33774,a33776,a33778,a33780,a33782,a33784,a33786,a33788,a33790,a33792,a33794,a33796,a33798,
a33800,a33802,a33804,a33806,a33808,a33810,a33812,a33814,a33816,a33818,a33820,a33822,a33824,a33826,a33828,
a33830,a33832,a33834,a33836,a33838,a33840,a33842,a33844,a33846,a33848,a33850,a33852,a33854,a33856,a33858,
a33860,a33862,a33864,a33866,a33868,a33870,a33872,a33874,a33876,a33878,a33880,a33882,a33884,a33886,a33888,
a33890,a33892,a33894,a33896,a33898,a33900,a33902,a33904,a33906,a33908,a33910,a33912,a33914,a33916,a33918,
a33920,a33922,a33924,a33926,a33928,a33930,a33932,a33934,a33936,a33938,a33940,a33942,a33944,a33946,a33948,
a33950,a33952,a33954,a33956,a33958,a33960,a33962,a33964,a33966,a33968,a33970,a33972,a33974,a33976,a33978,
a33980,a33982,a33984,a33986,a33988,a33990,a33992,a33994,a33996,a33998,a34000,a34002,a34004,a34006,a34008,
a34010,a34012,a34014,a34016,a34018,a34020,a34022,a34024,a34026,a34028,a34030,a34032,a34034,a34036,a34038,
a34040,a34042,a34044,a34046,a34048,a34050,a34052,a34054,a34056,a34058,a34060,a34062,a34064,a34066,a34068,
a34070,a34072,a34074,a34076,a34078,a34080,a34082,a34084,a34086,a34088,a34090,a34092,a34094,a34096,a34098,
a34100,a34102,a34104,a34106,a34108,a34110,a34112,a34114,a34116,a34118,a34120,a34122,a34124,a34126,a34128,
a34130,a34132,a34134,a34136,a34138,a34140,a34142,a34144,a34146,a34148,a34150,a34152,a34154,a34156,a34158,
a34160,a34162,a34164,a34166,a34168,a34170,a34172,a34174,a34178,a34180,a34182,a34184,a34186,a34188,a34190,
a34192,a34194,a34196,a34198,a34200,a34202,a34204,a34206,a34208,a34210,a34212,a34214,a34216,a34218,a34220,
a34222,a34224,a34226,a34228,a34230,a34232,a34234,a34236,a34238,a34240,a34242,a34244,a34246,a34248,a34250,
a34252,a34254,a34256,a34258,a34260,a34262,a34264,a34266,a34268,a34270,a34272,a34274,a34276,a34278,a34280,
a34282,a34284,a34286,a34288,a34290,a34292,a34294,a34296,a34298,a34300,a34302,a34304,a34306,a34308,a34310,
a34312,a34314,a34316,a34318,a34320,a34322,a34324,a34326,a34328,a34330,a34332,a34334,a34336,a34340,a34342,
a34344,a34346,a34348,a34350,a34352,a34354,a34356,a34358,a34360,a34364,a34366,a34368,a34370,a34372,a34374,
a34376,a34378,a34380,a34382,a34384,a34386,a34388,a34390,a34392,a34394,a34396,a34398,a34400,a34402,a34404,
a34406,a34408,a34410,a34412,a34414,a34416,a34418,a34420,a34422,a34424,a34426,a34428,a34430,a34432,a34434,
a34436,a34438,a34440,a34442,a34444,a34446,a34448,a34450,a34452,a34454,a34456,a34458,a34460,a34462,a34464,
a34466,a34468,a34470,a34472,a34474,a34476,a34478,a34480,a34482,a34484,a34486,a34490,a34492,a34496,a34498,
a34500,a34502,a34504,a34506,a34508,a34510,a34512,a34514,a34516,a34518,a34520,a34522,a34524,a34526,a34528,
a34530,a34532,a34534,a34536,a34538,a34540,a34542,a34544,a34546,a34548,a34550,a34552,a34556,a34558,a34562,
a34564,a34566,a34568,a34570,a34572,a34574,a34576,a34578,a34580,a34582,a34584,a34586,a34588,a34590,a34592,
a34594,a34596,a34598,a34600,a34602,a34604,a34606,a34608,a34610,a34612,a34614,a34616,a34618,a34622,a34624,
a34628,a34630,a34632,a34634,a34636,a34638,a34640,a34642,a34644,a34646,a34648,a34650,a34652,a34654,a34656,
a34658,a34660,a34662,a34664,a34666,a34668,a34670,a34672,a34674,a34676,a34678,a34680,a34682,a34684,a34688,
a34690,a34694,a34696,a34698,a34700,a34702,a34704,a34706,a34708,a34710,a34712,a34714,a34716,a34718,a34720,
a34722,a34724,a34726,a34728,a34730,a34732,a34734,a34736,a34738,a34740,a34742,a34744,a34746,a34748,a34750,
a34754,a34756,a34760,a34762,a34764,a34766,a34768,a34770,a34772,a34774,a34776,a34778,a34780,a34782,a34784,
a34786,a34788,a34790,a34792,a34794,a34796,a34798,a34800,a34802,a34804,a34806,a34808,a34810,a34812,a34814,
a34816,a34820,a34822,a34824,a34826,a34828,a34830,a34832,a34834,a34836,a34838,a34840,a34842,a34844,a34846,
a34848,a34850,a34852,a34854,a34856,a34858,a34860,a34862,a34864,a34866,a34868,a34870,a34872,a34874,a34876,
a34878,a34880,a34882,a34884,a34886,a34888,a34890,a34892,a34906,a34908,a34912,a34914,a34916,a34918,a34920,
a34922,a34924,a34926,a34928,a34930,a34932,a34934,a34936,a34938,a34940,a34942,a34944,a34946,a34948,a34950,
a34952,a34954,a34956,a34958,a34960,a34962,a34964,a34966,a34968,a34970,a34972,a34974,a34976,a34978,a34980,
a34982,a34984,a34986,a34990,a34992,a34994,a34996,a34998,a35002,a35004,a35006,a35008,a35010,a35012,a35014,
a35016,a35018,a35020,a35022,a35024,a35026,a35028,a35030,a35032,a35034,a35036,a35038,a35040,a35042,a35044,
a35046,a35048,a35050,a35052,a35056,a35058,a35060,a35062,a35064,a35068,a35070,a35072,a35074,a35076,a35078,
a35080,a35082,a35084,a35086,a35088,a35090,a35092,a35094,a35096,a35098,a35100,a35102,a35104,a35106,a35108,
a35110,a35112,a35114,a35116,a35118,a35122,a35124,a35126,a35128,a35130,a35134,a35136,a35138,a35140,a35142,
a35144,a35146,a35148,a35150,a35152,a35154,a35156,a35158,a35160,a35162,a35164,a35166,a35168,a35170,a35172,
a35174,a35176,a35178,a35180,a35182,a35184,a35188,a35190,a35192,a35194,a35196,a35200,a35202,a35204,a35206,
a35208,a35210,a35212,a35214,a35216,a35218,a35220,a35222,a35224,a35226,a35228,a35230,a35232,a35234,a35236,
a35238,a35240,a35242,a35244,a35246,a35248,a35250,a35254,a35256,a35258,a35260,a35262,a35266,a35268,a35270,
a35272,a35274,a35276,a35278,a35280,a35282,a35284,a35286,a35288,a35290,a35292,a35294,a35296,a35298,a35300,
a35302,a35304,a35306,a35308,a35310,a35312,a35314,a35316,a35318,a35320,a35322,a35324,a35326,a35328,a35332,
a35334,a35336,a35338,a35340,a35342,a35344,a35346,a35348,a35350,a35352,a35354,a35356,a35358,a35360,a35362,
a35364,a35366,a35368,a35370,a35372,a35374,a35376,a35378,a35380,a35382,a35384,a35386,a35388,a35390,a35392,
a35394,a35396,a35398,a35400,a35402,a35404,a35406,a35408,a35410,a35412,a35414,a35416,a35418,a35420,a35422,
a35424,a35426,a35428,a35430,a35432,a35434,a35436,a35438,a35440,a35442,a35444,a35446,a35448,a35450,a35452,
a35454,a35456,a35458,a35460,a35462,a35464,a35466,a35468,a35470,a35474,a35476,a35478,a35480,a35482,a35484,
a35486,a35488,a35490,a35492,a35494,a35496,a35498,a35500,a35502,a35504,a35506,a35508,a35510,a35512,a35516,
a35518,a35520,a35522,a35524,a35526,a35528,a35530,a35532,a35534,a35536,a35538,a35540,a35542,a35544,a35546,
a35548,a35550,a35552,a35556,a35558,a35560,a35562,a35564,a35566,a35568,a35570,a35572,a35574,a35576,a35578,
a35580,a35582,a35584,a35586,a35590,a35592,a35594,a35596,a35598,a35600,a35602,a35604,a35606,a35608,a35610,
a35612,a35614,a35616,a35618,a35620,a35622,a35624,a35626,a35628,a35630,a35632,a35634,a35638,a35640,a35642,
a35644,a35646,a35648,a35650,a35652,a35654,a35656,a35658,a35660,a35662,a35666,a35668,a35670,a35672,a35674,
a35676,a35678,a35680,a35682,a35684,a35686,a35688,a35690,a35692,a35694,a35696,a35698,a35702,a35704,a35706,
a35708,a35710,a35712,a35714,a35716,a35718,a35722,a35724,a35726,a35728,a35730,a35732,a35734,a35736,a35738,
a35740,a35742,a35744,a35746,a35750,a35752,a35754,a35756,a35758,a35760,a35762,a35764,a35766,a35768,a35770,
a35772,a35774,a35776,a35778,a35780,a35782,a35784,a35786,a35788,a35790,a35792,a35794,a35796,a35798,a35800,
a35802,a35804,a35806,a35808,a35810,a35812,a35814,a35816,a35818,a35820,a35822,a35824,a35826,a35828,a35830,
a35832,a35834,a35836,a35838,a35840,a35842,a35844,a35846,a35848,a35850,a35852,a35854,a35856,a35858,a35860,
a35862,a35864,a35866,a35868,a35870,a35872,a35874,a35876,a35878,a35880,a35882,a35884,a35886,a35888,a35890,
a35892,a35894,a35896,a35898,a35900,a35902,a35904,a35906,a35908,a35910,a35912,a35914,a35916,a35918,a35920,
a35922,a35924,a35926,a35928,a35932,a35934,a35936,a35938,a35940,a35942,a35944,a35948,a35950,a35952,a35954,
a35956,a35958,a35962,a35964,a35966,a35970,a35972,a35974,a35976,a35978,a35980,a35982,a35984,a35986,a35988,
a35990,a35992,a35994,a35996,a35998,a36000,a36002,a36004,a36006,a36008,a36010,a36012,a36014,a36016,a36018,
a36020,a36022,a36024,a36026,a36028,a36030,a36032,a36034,a36036,a36038,a36040,a36042,a36044,a36046,a36048,
a36050,a36052,a36054,a36056,a36058,a36060,a36062,a36064,a36066,a36068,a36070,a36072,a36074,a36076,a36078,
a36080,a36082,a36084,a36086,a36088,a36090,a36092,a36094,a36096,a36098,a36100,a36102,a36104,a36106,a36108,
a36110,a36112,a36114,a36116,a36118,a36120,a36122,a36124,a36126,a36128,a36130,a36132,a36134,a36136,a36138,
a36140,a36142,a36144,a36146,a36148,a36150,a36152,a36154,a36156,a36158,a36160,a36162,a36164,a36166,a36168,
a36170,a36172,a36174,a36176,a36178,a36180,a36182,a36184,a36186,a36188,a36190,a36192,a36194,a36196,a36198,
a36200,a36202,a36204,a36206,a36208,a36210,a36212,a36214,a36216,a36218,a36220,a36222,a36224,a36226,a36228,
a36230,a36232,a36234,a36236,a36238,a36240,a36242,a36244,a36246,a36248,a36250,a36252,a36254,a36256,a36258,
a36260,a36262,a36264,a36266,a36268,a36270,a36272,a36274,a36276,a36278,a36280,a36282,a36284,a36286,a36288,
a36290,a36292,a36294,a36296,a36298,a36300,a36302,a36304,a36306,a36308,a36310,a36312,a36314,a36316,a36318,
a36320,a36322,a36324,a36326,a36328,a36330,a36332,a36334,a36336,a36338,a36340,a36342,a36344,a36346,a36348,
a36350,a36352,a36354,a36356,a36358,a36360,a36362,a36364,a36366,a36368,a36370,a36372,a36374,a36376,a36378,
a36380,a36382,a36384,a36386,a36388,a36390,a36392,a36394,a36396,a36398,a36400,a36402,a36404,a36406,a36408,
a36410,a36412,a36414,a36416,a36418,a36420,a36422,a36424,a36426,a36428,a36430,a36432,a36434,a36436,a36438,
a36440,a36442,a36444,a36446,a36448,a36450,a36452,a36454,a36456,a36458,a36460,a36462,a36464,a36466,a36468,
a36470,a36472,a36474,a36476,a36478,a36480,a36482,a36484,a36486,a36488,a36490,a36492,a36494,a36496,a36498,
a36500,a36502,a36504,a36506,a36508,a36510,a36512,a36514,a36516,a36518,a36520,a36522,a36524,a36526,a36528,
a36530,a36532,a36534,a36536,a36538,a36540,a36542,a36544,a36546,a36548,a36550,a36552,a36554,a36556,a36558,
a36560,a36562,a36564,a36566,a36568,a36570,a36572,a36574,a36576,a36578,a36580,a36582,a36584,a36586,a36588,
a36590,a36592,a36594,a36596,a36598,a36600,a36602,a36604,a36606,a36608,a36610,a36612,a36614,a36616,a36618,
a36620,a36622,a36624,a36626,a36628,a36630,a36632,a36634,a36636,a36638,a36640,a36642,a36644,a36646,a36648,
a36650,a36652,a36654,a36656,a36658,a36660,a36662,a36664,a36666,a36668,a36670,a36672,a36674,a36676,a36678,
a36680,a36682,a36684,a36686,a36688,a36690,a36692,a36694,a36696,a36698,a36700,a36702,a36704,a36706,a36708,
a36710,a36712,a36714,a36716,a36718,a36720,a36722,a36724,a36726,a36728,a36730,a36732,a36734,a36736,a36738,
a36740,a36742,a36744,a36746,a36748,a36750,a36752,a36754,a36756,a36758,a36760,a36762,a36764,a36766,a36768,
a36770,a36772,a36774,a36776,a36778,a36780,a36782,a36784,a36786,a36788,a36790,a36792,a36794,a36796,a36798,
a36800,a36802,a36804,a36806,a36808,a36810,a36812,a36814,a36816,a36818,a36820,a36822,a36824,a36826,a36828,
a36830,a36832,a36834,a36836,a36838,a36840,a36842,a36844,a36846,a36848,a36850,a36852,a36854,a36856,a36858,
a36860,a36862,a36864,a36866,a36868,a36870,a36872,a36874,a36876,a36878,a36880,a36882,a36884,a36886,a36888,
a36890,a36892,a36894,a36896,a36898,a36900,a36902,a36904,a36906,a36908,a36910,a36912,a36914,a36916,a36918,
a36920,a36922,a36924,a36926,a36928,a36930,a36932,a36934,a36936,a36938,a36940,a36942,a36944,a36946,a36948,
a36950,a36952,a36954,a36956,a36958,a36960,a36962,a36964,a36966,a36968,a36970,a36972,a36974,a36976,a36978,
a36980,a36982,a36984,a36986,a36988,a36990,a36992,a36994,a36996,a36998,a37000,a37002,a37004,a37006,a37008,
a37010,a37012,a37014,a37016,a37018,a37020,a37022,a37024,a37026,a37028,a37030,a37032,a37034,a37036,a37038,
a37040,a37042,a37044,a37046,a37048,a37050,a37052,a37054,a37056,a37058,a37060,a37062,a37064,a37066,a37068,
a37070,a37072,a37074,a37076,a37078,a37080,a37082,a37084,a37086,a37088,a37090,a37092,a37094,a37096,a37098,
a37100,a37102,a37104,a37106,a37108,a37110,a37112,a37114,a37116,a37118,a37120,a37122,a37124,a37126,a37128,
a37130,a37132,a37134,a37136,a37138,a37140,a37142,a37144,a37146,a37148,a37150,a37152,a37154,a37156,a37158,
a37160,a37162,a37164,a37166,a37168,a37170,a37172,a37174,a37176,a37178,a37180,a37182,a37184,a37186,a37188,
a37190,a37192,a37194,a37196,a37198,a37200,a37202,a37204,a37206,a37208,a37210,a37212,a37214,a37216,a37218,
a37220,a37222,a37224,a37226,a37228,a37230,a37232,a37234,a37236,a37238,a37240,a37242,a37244,a37246,a37248,
a37250,a37252,a37254,a37256,a37258,a37260,a37262,a37264,a37266,a37268,a37270,a37272,a37274,a37276,a37278,
a37280,a37282,a37284,a37286,a37288,a37290,a37292,a37294,a37296,a37298,a37300,a37302,a37304,a37306,a37308,
a37310,a37312,a37314,a37316,a37318,a37320,a37322,a37324,a37326,a37328,a37330,a37332,a37334,a37336,a37338,
a37340,a37342,a37344,a37346,a37348,a37350,a37352,a37354,a37356,a37358,a37360,a37362,a37364,a37366,a37368,
a37370,a37372,a37374,a37376,a37378,a37380,a37382,a37384,a37386,a37388,a37390,a37392,a37394,a37396,a37398,
a37400,a37402,a37404,a37406,a37408,a37410,a37412,a37414,a37416,a37418,a37420,a37422,a37424,a37426,a37428,
a37430,a37432,a37434,a37436,a37438,a37440,a37442,a37444,a37446,a37448,a37450,a37452,a37454,a37456,a37458,
a37460,a37462,a37464,a37466,a37468,a37470,a37472,a37474,a37476,a37478,a37480,a37482,a37484,a37486,a37488,
a37490,a37492,a37494,a37496,a37498,a37500,a37502,a37504,a37506,a37508,a37510,a37512,a37514,a37516,a37518,
a37520,a37522,a37524,a37526,a37528,a37530,a37532,a37534,a37536,a37538,a37540,a37542,a37544,a37546,a37548,
a37550,a37552,a37554,a37556,a37558,a37560,a37562,a37564,a37566,a37568,a37570,a37572,a37574,a37576,a37578,
a37580,a37582,a37584,a37586,a37588,a37590,a37592,a37594,a37596,a37598,a37600,a37602,a37604,a37606,a37608,
a37610,a37612,a37614,a37616,a37618,a37620,a37622,a37624,a37626,a37628,a37630,a37632,a37634,a37636,a37638,
a37640,a37642,a37644,a37646,a37648,a37650,a37652,a37654,a37656,a37658,a37660,a37662,a37664,a37666,a37668,
a37670,a37672,a37674,a37676,a37678,a37680,a37682,a37684,a37686,a37688,a37690,a37692,a37694,a37696,a37698,
a37700,a37702,a37704,a37706,a37708,a37710,a37712,a37714,a37716,a37718,a37720,a37722,a37724,a37726,a37728,
a37730,a37732,a37734,a37736,a37738,a37740,a37742,a37744,a37746,a37748,a37750,a37752,a37754,a37756,a37758,
a37760,a37762,a37764,a37766,a37768,a37770,a37772,a37774,a37776,a37778,a37780,a37782,a37784,a37786,a37788,
a37790,a37792,a37794,a37796,a37798,a37800,a37802,a37804,a37806,a37808,a37810,a37812,a37814,a37816,a37818,
a37820,a37822,a37824,a37826,a37828,a37830,a37832,a37834,a37836,a37838,a37840,a37842,a37844,a37846,a37848,
a37850,a37852,a37854,a37856,a37858,a37860,a37862,a37864,a37866,a37868,a37870,a37872,a37874,a37876,a37878,
a37880,a37882,a37884,a37886,a37888,a37890,a37892,a37894,a37896,a37898,a37900,a37902,a37904,a37906,a37908,
a37910,a37912,a37914,a37916,a37918,a37920,a37922,a37924,a37926,a37928,a37930,a37932,a37934,a37936,a37938,
a37940,a37942,a37944,a37946,a37948,a37950,a37952,a37954,a37956,a37958,a37960,a37962,a37964,a37966,a37968,
a37970,a37972,a37974,a37976,a37978,a37980,a37982,a37984,a37986,a37988,a37990,a37992,a37994,a37996,a37998,
a38000,a38002,a38004,a38006,a38008,a38010,a38012,a38014,a38016,a38018,a38020,a38022,a38024,a38026,a38028,
a38030,a38032,a38034,a38036,a38038,a38040,a38042,a38044,a38046,a38048,a38050,a38052,a38054,a38056,a38058,
a38060,a38062,a38064,a38066,a38068,a38070,a38072,a38074,a38076,a38078,a38080,a38082,a38084,a38086,a38088,
a38090,a38092,a38094,a38096,a38098,a38100,a38102,a38104,a38106,a38108,a38110,a38112,a38114,a38116,a38118,
a38120,a38122,a38124,a38126,a38128,a38130,a38132,a38134,a38136,a38138,a38140,a38142,a38144,a38146,a38148,
a38150,a38152,a38154,a38156,a38158,a38160,a38162,a38164,a38166,a38168,a38170,a38172,a38174,a38176,a38178,
a38180,a38182,a38184,a38186,a38188,a38190,a38192,a38194,a38196,a38198,a38200,a38202,a38204,a38206,a38208,
a38210,a38212,a38214,a38216,a38218,a38220,a38222,a38224,a38226,a38228,a38230,a38232,a38234,a38236,a38238,
a38240,a38242,a38244,a38246,a38248,a38250,a38252,a38254,a38256,a38258,a38260,a38262,a38264,a38266,a38268,
a38270,a38272,a38274,a38276,a38278,a38280,a38282,a38284,a38286,a38288,a38290,a38292,a38294,a38296,a38298,
a38300,a38302,a38304,a38306,a38308,a38310,a38312,a38314,a38316,a38318,a38320,a38322,a38324,a38326,a38328,
a38330,a38332,a38334,a38336,a38338,a38340,a38342,a38344,a38346,a38348,a38350,a38352,a38354,a38356,a38358,
a38360,a38362,a38364,a38366,a38368,a38370,a38372,a38374,a38376,a38378,a38380,a38382,a38384,a38386,a38388,
a38390,a38392,a38394,a38396,a38398,a38400,a38402,a38404,a38406,a38408,a38410,a38412,a38414,a38416,a38418,
a38420,a38422,a38424,a38426,a38428,a38430,a38432,a38434,a38436,a38438,a38440,a38442,a38444,a38446,a38448,
a38450,a38452,a38454,a38456,a38458,a38460,a38462,a38464,a38466,a38468,a38470,a38472,a38474,a38476,a38478,
a38480,a38482,a38484,a38486,a38488,a38490,a38492,a38494,a38496,a38498,a38500,a38502,a38504,a38506,a38508,
a38510,a38512,a38514,a38516,a38518,a38520,a38522,a38524,a38526,a38528,a38530,a38532,a38534,a38536,a38538,
a38540,a38542,a38544,a38546,a38548,a38550,a38552,a38554,a38556,a38558,a38560,a38562,a38564,a38566,a38568,
a38570,a38572,a38574,a38576,a38578,a38580,a38582,a38584,a38586,a38588,a38590,a38592,a38594,a38596,a38598,
a38600,a38602,a38604,a38606,a38608,a38610,a38612,a38614,a38616,a38618,a38620,a38622,a38624,a38626,a38628,
a38630,a38632,a38634,a38636,a38638,a38640,a38642,a38644,a38646,a38648,a38650,a38652,a38654,a38656,a38658,
a38660,a38662,a38664,a38666,a38668,a38670,a38672,a38674,a38676,a38678,a38680,a38682,a38684,a38686,a38688,
a38690,a38692,a38694,a38696,a38698,a38700,a38702,a38704,a38706,a38708,a38710,a38712,a38714,a38716,a38718,
a38720,a38722,a38724,a38726,a38728,a38730,a38732,a38734,a38736,a38738,a38740,a38742,a38744,a38746,a38748,
a38750,a38752,a38754,a38756,a38758,a38760,a38762,a38764,a38766,a38768,a38770,a38772,a38774,a38776,a38778,
a38780,a38782,a38784,a38786,a38788,a38790,a38792,a38794,a38796,a38798,a38800,a38802,a38804,a38806,a38808,
a38810,a38812,a38814,a38816,a38818,a38820,a38822,a38824,a38826,a38828,a38830,a38832,a38834,a38836,a38838,
a38840,a38842,a38844,a38846,a38848,a38850,a38852,a38854,a38856,a38858,a38860,a38862,a38864,a38866,a38868,
a38870,a38872,a38874,a38876,a38878,a38880,a38882,a38884,a38886,a38888,a38890,a38892,a38894,a38896,a38898,
a38900,a38902,a38904,a38906,a38908,a38910,a38912,a38914,a38916,a38918,a38920,a38922,a38924,a38926,a38928,
a38930,a38932,a38934,a38936,a38938,a38940,a38942,a38944,a38946,a38948,a38950,a38952,a38954,a38956,a38958,
a38960,a38962,a38964,a38966,a38968,a38970,a38972,a38974,a38976,a38978,a38980,a38982,a38984,a38986,a38988,
a38990,a38992,a38994,a38996,a38998,a39000,a39002,a39004,a39006,a39008,a39010,a39012,a39014,a39016,a39018,
a39020,a39022,a39024,a39026,a39028,a39030,a39032,a39034,a39036,a39038,a39040,a39042,a39044,a39046,a39048,
a39050,a39052,a39054,a39056,a39058,a39060,a39062,a39064,a39066,a39068,a39070,a39072,a39074,a39076,a39078,
a39080,a39082,a39084,a39086,a39088,a39090,a39092,a39094,a39096,a39098,a39100,a39102,a39104,a39106,a39108,
a39110,a39112,a39114,a39116,a39118,a39120,a39122,a39124,a39126,a39128,a39130,a39132,a39134,a39136,a39138,
a39140,a39142,a39144,a39146,a39148,a39150,a39152,a39154,a39156,a39158,a39160,a39162,a39164,a39166,a39168,
a39170,a39172,a39174,a39176,a39178,a39180,a39182,a39184,a39186,a39188,a39190,a39192,a39194,a39196,a39198,
a39200,a39202,a39204,a39206,a39208,a39210,a39212,a39214,a39216,a39218,a39220,a39222,a39224,a39226,a39228,
a39230,a39232,a39234,a39236,a39238,a39240,a39242,a39244,a39246,a39248,a39250,a39252,a39254,a39256,a39258,
a39260,a39262,a39264,a39266,a39268,a39270,a39272,a39274,a39276,a39278,a39280,a39282,a39284,a39286,a39288,
a39290,a39292,a39294,a39296,a39298,a39300,a39302,a39304,a39306,a39308,a39310,a39312,a39314,a39316,a39318,
a39320,a39322,a39324,a39326,a39328,a39330,a39332,a39334,a39336,a39338,a39340,a39342,a39344,a39346,a39348,
a39350,a39352,a39354,a39356,a39358,a39360,a39362,a39364,a39366,a39368,a39370,a39372,a39374,a39376,a39378,
a39380,a39382,a39384,a39386,a39388,a39390,a39392,a39394,a39396,a39398,a39400,a39402,a39404,a39406,a39408,
a39410,a39412,a39414,a39416,a39418,a39420,a39422,a39424,a39426,a39428,a39430,a39432,a39434,a39436,a39438,
a39440,a39442,a39444,a39446,a39448,a39450,a39452,a39454,a39456,a39458,a39460,a39462,a39464,a39466,a39468,
a39470,a39472,a39474,a39476,a39478,a39480,a39482,a39484,a39486,a39488,a39490,a39492,a39494,a39496,a39498,
a39500,a39502,a39504,a39506,a39508,a39510,a39512,a39514,a39516,a39518,a39520,a39522,a39524,a39526,a39528,
a39530,a39532,a39534,a39536,a39538,a39540,a39542,a39544,a39546,a39548,a39550,a39552,a39554,a39556,a39558,
a39560,a39562,a39564,a39566,a39568,a39570,a39572,a39574,a39576,a39578,a39580,a39582,a39584,a39586,a39588,
a39590,a39592,a39594,a39596,a39598,a39600,a39602,a39604,a39606,a39608,a39610,a39612,a39614,a39616,a39618,
a39620,a39622,a39624,a39626,a39628,a39630,a39632,a39634,a39636,a39638,a39640,a39642,a39644,a39646,a39648,
a39650,a39652,a39654,a39656,a39658,a39660,a39662,a39664,a39666,a39668,a39670,a39672,a39674,a39676,a39678,
a39680,a39682,a39684,a39686,a39688,a39690,a39692,a39694,a39696,a39698,a39700,a39702,a39704,a39706,a39708,
a39710,a39712,a39714,a39716,a39718,a39720,a39722,a39724,a39726,a39728,a39730,a39732,a39734,a39736,a39738,
a39740,a39742,a39744,a39746,a39748,a39750,a39752,a39754,a39756,a39758,a39760,a39762,a39764,a39766,a39768,
a39770,a39772,a39774,a39776,a39778,a39780,a39782,a39784,a39786,a39788,a39790,a39792,a39794,a39796,a39798,
a39800,a39802,a39804,a39806,a39808,a39810,a39812,a39814,a39816,a39818,a39820,a39822,a39824,a39826,a39828,
a39830,a39832,a39834,a39836,a39838,a39840,a39842,a39844,a39846,a39848,a39850,a39852,a39854,a39856,a39858,
a39860,a39862,a39864,a39866,a39868,a39870,a39872,a39874,a39876,a39878,a39880,a39882,a39884,a39886,a39888,
a39890,a39892,a39894,a39896,a39898,a39900,a39902,a39904,a39906,a39908,a39910,a39912,a39914,a39916,a39918,
a39920,a39922,a39924,a39926,a39928,a39930,a39932,a39934,a39936,a39938,a39940,a39942,a39944,a39946,a39948,
a39950,a39952,a39954,a39956,a39958,a39960,a39962,a39964,a39966,a39968,a39970,a39972,a39974,a39976,a39978,
a39980,a39982,a39984,a39986,a39988,a39990,a39992,a39994,a39996,a39998,a40000,a40002,a40004,a40006,a40008,
a40010,a40012,a40014,a40016,a40018,a40020,a40022,a40024,a40026,a40028,a40030,a40032,a40034,a40036,a40038,
a40040,a40042,a40044,a40046,a40048,a40050,a40052,a40054,a40056,a40058,a40060,a40062,a40064,a40066,a40068,
a40070,a40072,a40074,a40076,a40078,a40080,a40082,a40084,a40086,a40088,a40090,a40092,a40094,a40096,a40098,
a40100,a40102,a40104,a40106,a40108,a40110,a40112,a40114,a40116,a40118,a40120,a40122,a40124,a40126,a40128,
a40130,a40132,a40134,a40136,a40138,a40140,a40142,a40144,a40146,a40148,a40150,a40152,a40154,a40156,a40158,
a40160,a40162,a40164,a40166,a40168,a40170,a40172,a40174,a40176,a40178,a40180,a40182,a40184,a40186,a40188,
a40190,a40192,a40194,a40196,a40198,a40200,a40202,a40204,a40206,a40208,a40210,a40212,a40214,a40216,a40218,
a40220,a40222,a40224,a40226,a40228,a40230,a40232,a40234,a40236,a40238,a40240,a40242,a40244,a40246,a40248,
a40250,a40252,a40254,a40256,a40258,a40260,a40262,a40264,a40266,a40268,a40270,a40272,a40274,a40276,a40278,
a40280,a40282,a40284,a40286,a40288,a40290,a40292,a40294,a40296,a40298,a40300,a40302,a40304,a40306,a40308,
a40310,a40312,a40314,a40316,a40318,a40320,a40322,a40324,a40326,a40328,a40330,a40332,a40334,a40336,a40338,
a40340,a40342,a40344,a40346,a40348,a40350,a40352,a40354,a40356,a40358,a40360,a40362,a40364,a40366,a40368,
a40370,a40372,a40374,a40376,a40378,a40380,a40382,a40384,a40386,a40388,a40390,a40392,a40394,a40396,a40398,
a40400,a40402,a40404,a40406,a40408,a40410,a40412,a40414,a40416,a40418,a40420,a40422,a40424,a40426,a40428,
a40430,a40432,a40434,a40436,a40438,a40440,a40442,a40444,a40446,a40448,a40450,a40452,a40454,a40456,a40458,
a40460,a40462,a40464,a40466,a40468,a40470,a40472,a40474,a40476,a40478,a40480,a40482,a40484,a40486,a40488,
a40490,a40492,a40494,a40496,a40498,a40500,a40502,a40504,a40506,a40508,a40510,a40512,a40514,a40516,a40518,
a40520,a40522,a40524,a40526,a40528,a40530,a40532,a40534,a40536,a40538,a40540,a40542,a40544,a40546,a40548,
a40550,a40552,a40554,a40556,a40558,a40560,a40562,a40564,a40566,a40568,a40570,a40572,a40574,a40576,a40578,
a40580,a40582,a40584,a40586,a40588,a40590,a40592,a40594,a40596,a40598,a40600,a40602,a40604,a40606,a40608,
a40610,a40612,a40614,a40616,a40618,a40620,a40622,a40624,a40626,a40628,a40630,a40632,a40634,a40636,a40638,
a40640,a40644,a40646,a40648,a40650,a40652,a40654,a40656,a40658,a40660,a40662,a40664,a40666,a40668,a40670,
a40672,a40674,a40676,a40678,a40680,a40682,a40684,a40686,a40688,a40690,a40692,a40694,a40696,a40698,a40700,
a40702,a40704,a40706,a40708,a40710,a40712,a40714,a40716,a40718,a40720,a40722,a40724,a40726,a40728,a40730,
a40732,a40734,a40736,a40738,a40740,a40742,a40744,a40746,a40748,a40750,a40752,a40754,a40756,a40758,a40760,
a40762,a40764,a40766,a40768,a40770,a40772,a40774,a40776,a40778,a40780,a40782,a40784,a40786,a40788,a40790,
a40792,a40794,a40796,a40798,a40800,a40802,a40804,a40806,a40808,a40810,a40812,a40814,a40816,a40818,a40820,
a40822,a40824,a40826,a40828,a40830,a40832,a40834,a40836,a40838,a40840,a40842,a40844,a40846,a40848,a40850,
a40852,a40854,a40856,a40858,a40860,a40862,a40864,a40866,a40868,a40870,a40872,a40874,a40876,a40878,a40880,
a40882,a40884,a40886,a40888,a40890,a40892,a40894,a40896,a40898,a40900,a40902,a40904,a40906,a40908,a40910,
a40912,a40914,a40916,a40918,a40920,a40922,a40924,a40926,a40928,a40930,a40932,a40934,a40936,a40938,a40940,
a40942,a40944,a40946,a40948,a40950,a40952,a40954,a40956,a40958,a40960,a40962,a40964,a40966,a40968,a40970,
a40972,a40974,a40976,a40978,a40980,a40982,a40984,a40986,a40988,a40990,a40992,a40994,a40996,a40998,a41000,
a41002,a41004,a41006,a41008,a41010,a41012,a41014,a41016,a41018,a41020,a41022,a41024,a41026,a41028,a41030,
a41032,a41034,a41036,a41038,a41040,a41042,a41044,a41046,a41048,a41050,a41052,a41054,a41056,a41058,a41060,
a41062,a41064,a41066,a41068,a41070,a41072,a41074,a41076,a41078,a41080,a41082,a41084,a41086,a41088,a41090,
a41092,a41094,a41096,a41098,a41100,a41102,a41104,a41106,a41108,a41110,a41112,a41114,a41116,a41118,a41120,
a41122,a41124,a41126,a41128,a41130,a41132,a41134,a41136,a41138,a41140,a41142,a41144,a41146,a41148,a41150,
a41152,a41154,a41156,a41158,a41160,a41162,a41164,a41166,a41168,a41170,a41172,a41174,a41176,a41178,a41180,
a41182,a41184,a41186,a41188,a41190,a41192,a41194,a41196,a41198,a41200,a41202,a41204,a41206,a41208,a41210,
a41212,a41214,a41216,a41218,a41220,a41222,a41224,a41226,a41228,a41230,a41232,a41234,a41236,a41238,a41240,
a41242,a41244,a41246,a41248,a41250,a41252,a41254,a41256,a41258,a41260,a41262,a41264,a41266,a41268,a41270,
a41272,a41274,a41276,a41278,a41280,a41282,a41284,a41286,a41288,a41290,a41292,a41294,a41296,a41298,a41300,
a41302,a41304,a41306,a41308,a41310,a41312,a41314,a41316,a41318,a41320,a41322,a41324,a41326,a41328,a41330,
a41332,a41334,a41336,a41338,a41340,a41342,a41344,a41346,a41348,a41350,a41352,a41354,a41356,a41358,a41360,
a41362,a41364,a41366,a41368,a41370,a41372,a41374,a41376,a41378,a41380,a41382,a41384,a41386,a41388,a41390,
a41392,a41394,a41396,a41398,a41400,a41402,a41404,a41406,a41408,a41410,a41412,a41414,a41416,a41418,a41420,
a41422,a41424,a41426,a41428,a41430,a41432,a41434,a41436,a41438,a41440,a41442,a41444,a41446,a41448,a41450,
a41452,a41454,a41456,a41458,a41460,a41462,a41464,a41466,a41468,a41470,a41472,a41474,a41476,a41478,a41480,
a41482,a41484,a41486,a41488,a41490,a41492,a41494,a41496,a41498,a41500,a41502,a41504,a41506,a41508,a41510,
a41512,a41514,a41516,a41518,a41520,a41522,a41524,a41526,a41528,a41530,a41532,a41534,a41536,a41538,a41540,
a41542,a41544,a41546,a41548,a41550,a41552,a41554,a41556,a41558,a41560,a41562,a41564,a41566,a41568,a41570,
a41572,a41574,a41576,a41578,a41580,a41582,a41584,a41586,a41588,a41590,a41592,a41594,a41596,a41598,a41600,
a41602,a41604,a41606,a41608,a41610,a41612,a41614,a41616,a41618,a41620,a41622,a41624,a41626,a41628,a41630,
a41632,a41634,a41636,a41640,a41642,a41646,a41648,a41650,a41652,a41656,a41658,a41660,a41662,a41664,a41666,
a41668,a41674,a41676,a41678,a41680,a41682,a41684,a41686,a41688,a41690,a41692,a41694,a41696,a41698,a41700,
a41702,a41704,a41706,a41708,a41710,a41712,a41714,a41716,a41718,a41720,a41722,a41724,a41726,a41728,a41730,
a41732,a41734,a41738,a41740,a41742,a41744,a41746,a41748,a41750,a41752,a41754,a41756,a41758,a41760,a41762,
a41764,a41766,a41768,a41770,a41772,a41774,a41776,a41778,a41780,a41782,a41784,a41786,a41788,a41790,a41792,
a41794,a41796,a41798,a41800,a41802,a41804,a41806,a41808,a41810,a41812,a41814,a41816,a41818,a41820,a41822,
a41824,a41826,a41828,a41830,a41832,a41834,a41836,a41838,a41840,a41842,a41844,a41846,a41848,a41850,a41852,
a41854,a41856,a41858,a41860,a41862,a41864,a41866,a41868,a41870,a41872,a41874,a41876,a41878,a41880,a41882,
a41884,a41886,a41888,a41890,a41892,a41894,a41896,a41898,a41900,a41902,a41904,a41906,a41908,a41910,a41912,
a41914,a41916,a41918,a41920,a41922,a41924,a41926,a41928,a41930,a41932,a41934,a41936,a41938,a41940,a41942,
a41944,a41946,a41948,a41950,a41952,a41954,a41956,a41958,a41960,a41962,a41964,a41966,a41968,a41970,a41972,
a41974,a41976,a41978,a41980,a41982,a41984,a41986,a41988,a41990,a41992,a41994,a41996,a41998,a42000,a42002,
a42004,a42006,a42008,a42010,a42012,a42014,a42016,a42018,a42020,a42022,a42024,a42026,a42028,a42030,a42032,
a42034,a42036,a42038,a42040,a42042,a42044,a42046,a42048,a42050,a42052,a42054,a42056,a42058,a42060,a42062,
a42064,a42066,a42068,a42070,a42072,a42074,a42076,a42078,a42080,a42082,a42084,a42086,a42088,a42090,a42092,
a42094,a42096,a42098,a42100,a42102,a42104,a42106,a42108,a42110,a42112,a42114,a42116,a42118,a42120,a42122,
a42124,a42126,a42128,a42130,a42132,a42134,a42136,a42138,a42140,a42142,a42144,a42146,a42148,a42150,a42152,
a42154,a42156,a42158,a42160,a42162,a42164,a42166,a42168,a42170,a42172,a42174,a42176,a42178,a42180,a42182,
a42184,a42186,a42188,a42190,a42192,a42194,a42196,a42198,a42200,a42202,a42204,a42206,a42208,a42210,a42212,
a42214,a42216,a42218,a42220,a42222,a42224,a42226,a42228,a42230,a42232,a42234,a42236,a42238,a42240,a42242,
a42244,a42246,a42248,a42250,a42252,a42254,a42256,a42258,a42260,a42262,a42264,a42266,a42268,a42270,a42272,
a42274,a42276,a42278,a42280,a42282,a42284,a42286,a42288,a42290,a42292,a42294,a42296,a42298,a42300,a42302,
a42304,a42306,a42308,a42310,a42312,a42314,a42316,a42318,a42320,a42322,a42324,a42326,a42328,a42330,a42332,
a42334,a42336,a42338,a42340,a42342,a42344,a42346,a42348,a42350,a42352,a42354,a42356,a42358,a42360,a42362,
a42364,a42366,a42368,a42370,a42372,a42374,a42376,a42378,a42380,a42382,a42384,a42386,a42388,a42390,a42392,
a42394,a42396,a42398,a42400,a42402,a42404,a42406,a42408,a42410,a42412,a42414,a42416,a42418,a42420,a42422,
a42424,a42426,a42428,a42430,a42432,a42434,a42436,a42438,a42440,a42442,a42444,a42446,a42448,a42450,a42452,
a42454,a42456,a42458,a42460,a42462,a42464,a42466,a42468,a42470,a42472,a42474,a42476,a42478,a42480,a42482,
a42484,a42486,a42488,a42490,a42492,a42494,a42496,a42498,a42500,a42502,a42504,a42506,a42508,a42510,a42512,
a42514,a42516,a42518,a42520,a42522,a42524,a42526,a42528,a42530,a42532,a42534,a42536,a42538,a42540,a42542,
a42544,a42546,a42548,a42550,a42552,a42554,a42556,a42558,a42560,a42562,a42564,a42566,a42568,a42570,a42572,
a42574,a42576,a42578,a42580,a42582,a42584,a42586,a42588,a42590,a42592,a42594,a42596,a42598,a42600,a42602,
a42604,a42606,a42608,a42610,a42612,a42614,a42616,a42618,a42620,a42622,a42624,a42626,a42628,a42630,a42632,
a42634,a42636,a42638,a42640,a42642,a42644,a42646,a42648,a42650,a42652,a42654,a42656,a42658,a42660,a42662,
a42664,a42666,a42668,a42670,a42672,a42674,a42676,a42678,a42680,a42682,a42684,a42686,a42688,a42690,a42692,
a42694,a42696,a42698,a42700,a42702,a42704,a42706,a42708,a42710,a42712,a42714,a42716,a42718,a42720,a42722,
a42724,a42726,a42728,a42730,a42732,a42734,a42736,a42738,a42740,a42742,a42744,a42746,a42748,a42750,a42752,
a42754,a42756,a42758,a42760,a42762,a42764,a42766,a42768,a42770,a42772,a42774,a42776,a42778,a42780,a42782,
a42784,a42786,a42788,a42790,a42792,a42794,a42796,a42798,a42800,a42802,a42804,a42806,a42808,a42810,a42812,
a42814,a42816,a42818,a42820,a42822,a42824,a42826,a42828,a42830,a42832,a42834,a42836,a42838,a42840,a42842,
a42844,a42846,a42848,a42850,a42852,a42854,a42856,a42858,a42860,a42862,a42864,a42866,a42868,a42870,a42872,
a42874,a42876,a42878,a42880,a42882,a42884,a42886,a42888,a42890,a42892,a42894,a42896,a42898,a42900,a42902,
a42904,a42906,a42908,a42910,a42912,a42914,a42916,a42918,a42920,a42922,a42924,a42926,a42928,a42930,a42932,
a42934,a42936,a42938,a42940,a42942,a42944,a42946,a42948,a42950,a42952,a42954,a42956,a42958,a42960,a42962,
a42964,a42966,a42968,a42970,a42972,a42974,a42976,a42978,a42980,a42982,a42984,a42986,a42988,a42990,a42992,
a42994,a42996,a42998,a43000,a43002,a43004,a43006,a43008,a43010,a43012,a43014,a43016,a43018,a43020,a43022,
a43024,a43026,a43028,a43030,a43032,a43034,a43036,a43038,a43040,a43042,a43044,a43046,a43048,a43050,a43052,
a43054,a43056,a43058,a43060,a43062,a43064,a43066,a43068,a43070,a43072,a43074,a43076,a43078,a43080,a43082,
a43084,a43086,a43088,a43090,a43092,a43094,a43096,a43098,a43100,a43102,a43104,a43106,a43108,a43110,a43112,
a43114,a43116,a43118,a43120,a43122,a43124,a43126,a43128,a43130,a43132,a43134,a43136,a43138,a43140,a43142,
a43144,a43146,a43148,a43150,a43152,a43154,a43156,a43158,a43160,a43162,a43164,a43166,a43168,a43170,a43172,
a43174,a43176,a43178,a43180,a43182,a43184,a43186,a43188,a43190,a43192,a43194,a43196,a43198,a43200,a43202,
a43204,a43206,a43208,a43210,a43212,a43214,a43216,a43218,a43220,a43222,a43224,a43226,a43228,a43230,a43232,
a43234,a43236,a43238,a43240,a43242,a43244,a43246,a43248,a43250,a43252,a43254,a43256,a43258,a43260,a43262,
a43264,a43266,a43268,a43270,a43272,a43274,a43276,a43278,a43280,a43282,a43284,a43286,a43288,a43290,a43292,
a43294,a43296,a43298,a43300,a43302,a43304,a43306,a43308,a43310,a43312,a43314,a43316,a43318,a43320,a43322,
a43324,a43326,a43328,a43330,a43332,a43334,a43336,a43338,a43340,a43342,a43344,a43346,a43348,a43350,a43352,
a43354,a43356,a43358,a43360,a43362,a43364,a43366,a43368,a43370,a43372,a43374,a43376,a43378,a43380,a43382,
a43384,a43386,a43388,a43390,a43392,a43394,a43396,a43398,a43400,a43402,a43404,a43406,a43408,a43410,a43412,
a43414,a43416,a43418,a43420,a43422,a43424,a43426,a43428,a43430,a43432,a43434,a43436,a43438,a43440,a43442,
a43444,a43446,a43448,a43450,a43452,a43454,a43456,a43458,a43460,a43462,a43464,a43466,a43468,a43470,a43472,
a43474,a43476,a43478,a43480,a43482,a43484,a43486,a43488,a43490,a43492,a43494,a43496,a43498,a43500,a43502,
a43504,a43506,a43508,a43510,a43512,a43514,a43516,a43518,a43520,a43522,a43524,a43526,a43528,a43530,a43532,
a43534,a43536,a43538,a43540,a43542,a43544,a43546,a43548,a43550,a43552,a43554,a43556,a43558,a43560,a43562,
a43564,a43566,a43568,a43570,a43572,a43574,a43576,a43578,a43580,a43582,a43584,a43586,a43588,a43590,a43592,
a43594,a43596,a43598,a43600,a43602,a43604,a43606,a43608,a43610,a43612,a43614,a43616,a43618,a43620,a43622,
a43624,a43626,a43628,a43630,a43632,a43634,a43636,a43638,a43640,a43642,a43644,a43646,a43648,a43650,a43652,
a43654,a43656,a43658,a43660,a43662,a43664,a43666,a43668,a43670,a43672,a43674,a43676,a43678,a43680,a43682,
a43684,a43686,a43688,a43690,a43692,a43694,a43696,a43698,a43700,a43702,a43704,a43706,a43708,a43710,a43712,
a43714,a43716,a43718,a43720,a43722,a43724,a43726,a43728,a43730,a43732,a43734,a43736,a43738,a43740,a43742,
a43744,a43746,a43748,a43750,a43752,a43754,a43756,a43758,a43760,a43762,a43764,a43766,a43768,a43770,a43772,
a43774,a43776,a43778,a43780,a43782,a43784,a43786,a43788,a43790,a43792,a43794,a43796,a43798,a43800,a43802,
a43804,a43806,a43808,a43810,a43812,a43814,a43816,a43818,a43820,a43822,a43824,a43826,a43828,a43830,a43832,
a43834,a43836,a43838,a43840,a43842,a43844,a43846,a43848,a43850,a43852,a43854,a43856,a43858,a43860,a43862,
a43864,a43866,a43868,a43870,a43872,a43874,a43876,a43878,a43880,a43882,a43884,a43886,a43888,a43890,a43892,
a43894,a43896,a43898,a43900,a43902,a43904,a43906,a43908,a43910,a43912,a43914,a43916,a43918,a43920,a43922,
a43924,a43926,a43928,a43930,a43932,a43934,a43936,a43938,a43940,a43942,a43944,a43946,a43948,a43950,a43952,
a43954,a43956,a43958,a43960,a43962,a43964,a43966,a43968,a43970,a43972,a43974,a43976,a43978,a43980,a43982,
a43984,a43986,a43988,a43990,a43992,a43994,a43996,a43998,a44000,a44002,a44004,a44006,a44008,a44010,a44012,
a44014,a44016,a44018,a44020,a44022,a44024,a44026,a44028,a44030,a44032,a44034,a44036,a44038,a44040,a44042,
a44044,a44046,a44048,a44050,a44052,a44054,a44056,a44058,a44060,a44062,a44064,a44066,a44068,a44070,a44072,
a44074,a44076,a44078,a44080,a44082,a44084,a44086,a44088,a44090,a44092,a44094,a44096,a44098,a44100,a44102,
a44104,a44106,a44108,a44110,a44112,a44114,a44116,a44118,a44120,a44122,a44124,a44126,a44128,a44130,a44132,
a44134,a44136,a44138,a44140,a44142,a44144,a44146,a44148,a44150,a44152,a44154,a44156,a44158,a44160,a44162,
a44164,a44166,a44168,a44170,a44172,a44174,a44176,a44178,a44180,a44182,a44184,a44186,a44188,a44190,a44192,
a44194,a44196,a44198,a44200,a44202,a44204,a44206,a44208,a44210,a44212,a44214,a44216,a44218,a44220,a44222,
a44224,a44226,a44228,a44230,a44232,a44234,a44236,a44238,a44240,a44242,a44244,a44246,a44248,a44250,a44252,
a44254,a44256,a44258,a44260,a44262,a44264,a44266,a44268,a44270,a44272,a44274,a44276,a44278,a44280,a44282,
a44284,a44286,a44288,a44290,a44292,a44294,a44296,a44298,a44300,a44302,a44304,a44306,a44308,a44310,a44312,
a44314,a44316,a44318,a44320,a44322,a44324,a44326,a44328,a44330,a44332,a44334,a44336,a44338,a44340,a44342,
a44344,a44346,a44348,a44350,a44352,a44354,a44356,a44358,a44360,a44362,a44364,a44366,a44368,a44370,a44372,
a44374,a44376,a44378,a44380,a44382,a44384,a44386,a44388,a44390,a44392,a44394,a44396,a44398,a44400,a44402,
a44404,a44406,a44410,a44412,a44414,a44416,a44418,a44420,a44422,a44424,a44426,a44430,a44432,a44434,a44436,
a44438,a44440,a44444,a44446,a44448,a44452,a44454,a44456,a44458,a44460,a44464,a44466,a44468,a44470,a44474,
a44476,a44478,a44480,a44484,a44486,a44488,a44492,a44494,a44496,a44500,a44502,a44504,a44508,a44510,a44512,
a44516,a44518,a44522,a44524,a44528,a44530,a44534,a44536,a44540,a44542,a44546,a44548,a44552,a44554,a44558,
a44560,a44564,a44566,a44570,a44572,a44576,a44578,a44582,a44584,a44588,a44590,a44594,a44596,a44600,a44602,
a44606,a44608,a44612,a44614,a44618,a44620,a44624,a44626,a44630,a44632,a44636,a44638,a44642,a44644,a44648,
a44650,a44654,a44656,a44660,a44662,a44666,a44668,a44672,a44674,a44678,a44680,a44684,a44686,a44690,a44692,
a44696,a44698,a44702,a44704,a44708,a44710,a44714,a44716,a44720,a44722,a44726,a44728,a44732,a44734,a44738,
a44740,a44744,a44746,a44750,a44752,a44756,a44758,a44762,a44764,a44768,a44770,a44774,a44776,a44780,a44782,
a44786,a44788,a44792,a44794,a44798,a44800,a44804,a44806,a44810,a44812,a44816,a44818,a44820,a44822,a44824,
a44826,a44828,a44830,a44832,a44836,a44838,a44840,a44842,a44844,a44846,a44848,a44850,a44852,a44854,a44856,
a44858,a44860,a44862,a44864,a44866,a44868,a44870,a44872,a44874,a44876,a44878,a44880,a44882,a44884,a44886,
a44888,a44890,a44892,a44894,a44896,a44898,a44900,a44902,a44904,a44906,a44908,a44910,a44912,a44914,a44916,
a44918,a44920,a44922,a44924,a44926,a44928,a44930,a44932,a44934,a44936,a44938,a44940,a44942,a44944,a44946,
a44948,a44950,a44952,a44954,a44956,a44958,a44960,a44962,a44964,a44966,a44968,a44970,a44972,a44974,a44976,
a44978,a44980,a44982,a44984,a44986,a44988,a44990,a44992,a44994,a44996,a44998,a45000,a45002,a45004,a45006,
a45008,a45010,a45012,a45014,a45016,a45018,a45020,a45022,a45024,a45026,a45028,a45030,a45032,a45034,a45036,
a45038,a45040,a45042,a45044,a45046,a45048,a45050,a45052,a45054,a45056,a45058,a45060,a45062,a45064,a45066,
a45068,a45070,a45072,a45074,a45076,a45078,a45080,a45082,a45084,a45086,a45088,a45090,a45092,a45094,a45096,
a45098,a45100,a45102,a45104,a45106,a45108,a45110,a45112,a45114,a45116,a45118,a45120,a45122,a45124,a45126,
a45128,a45130,a45132,a45134,a45136,a45138,a45140,a45142,a45144,a45146,a45148,a45150,a45152,a45154,a45156,
a45158,a45160,a45162,a45164,a45166,a45168,a45170,a45172,a45174,a45176,a45178,a45180,a45182,a45184,a45186,
a45188,a45190,a45192,a45194,a45196,a45198,a45200,a45202,a45204,a45206,a45208,a45210,a45212,a45214,a45216,
a45218,a45220,a45222,a45224,a45226,a45228,a45230,a45232,a45234,a45236,a45238,a45240,a45242,a45244,a45246,
a45248,a45250,a45252,a45254,a45256,a45258,a45260,a45262,a45264,a45266,a45268,a45270,a45272,a45274,a45276,
a45278,a45280,a45282,a45284,a45286,a45288,a45290,a45292,a45294,a45296,a45298,a45300,a45302,a45304,a45306,
a45308,a45310,a45312,a45314,a45316,a45318,a45320,a45322,a45324,a45326,a45328,a45330,a45332,a45334,a45336,
a45338,a45340,a45342,a45344,a45346,a45348,a45350,a45352,a45354,a45356,a45358,a45360,a45362,a45364,a45366,
a45368,a45370,a45372,a45374,a45376,a45378,a45380,a45382,a45384,a45386,a45388,a45390,a45392,a45394,a45396,
a45398,a45400,a45402,a45404,a45406,a45408,a45410,a45412,a45414,a45416,a45418,a45420,a45422,a45424,a45426,
a45428,a45430,a45432,a45434,a45436,a45438,a45440,a45442,a45444,a45446,a45448,a45450,a45452,a45454,a45456,
a45458,a45460,a45462,a45464,a45466,a45468,a45470,a45472,a45474,a45476,a45478,a45480,a45482,a45484,a45486,
a45488,a45490,a45492,a45494,a45496,a45498,a45500,a45502,a45504,a45506,a45508,a45510,a45512,a45514,a45516,
a45518,a45520,a45522,a45524,a45526,a45528,a45530,a45532,a45534,a45536,a45538,a45540,a45542,a45544,a45546,
a45548,a45550,a45552,a45554,a45556,a45558,a45560,a45562,a45564,a45566,a45568,a45570,a45572,a45574,a45576,
a45578,a45580,a45582,a45584,a45586,a45588,a45590,a45592,a45594,a45598,a45600,a45602,a45604,a45606,a45610,
a45612,a45614,a45616,a45618,a45620,a45624,a45626,a45628,a45630,a45632,a45634,a45636,a45638,a45640,a45642,
a45644,a45646,a45648,a45650,a45652,a45654,a45656,a45658,a45660,a45662,a45664,a45666,a45668,a45670,a45672,
a45674,a45676,a45678,a45680,a45682,a45684,a45686,a45688,a45690,a45692,a45694,a45696,a45698,a45700,a45702,
a45704,a45706,a45708,a45710,a45712,a45714,a45716,a45718,a45720,a45722,a45724,a45726,a45728,a45730,a45732,
a45734,a45736,a45738,a45740,a45742,a45744,a45746,a45748,a45750,a45752,a45754,a45756,a45758,a45760,a45762,
a45764,a45766,a45768,a45770,a45772,a45774,a45776,a45778,a45780,a45782,a45784,a45786,a45788,a45790,a45792,
a45794,a45796,a45798,a45800,a45802,a45804,a45806,a45808,a45810,a45812,a45814,a45816,a45818,a45820,a45822,
a45824,a45826,a45828,a45830,a45832,a45834,a45836,a45838,a45840,a45842,a45844,a45846,a45848,a45850,a45852,
a45854,a45856,a45858,a45860,a45862,a45864,a45866,a45868,a45870,a45872,a45874,a45876,a45878,a45880,a45882,
a45884,a45886,a45888,a45890,a45892,a45894,a45896,a45898,a45900,a45902,a45904,a45906,a45908,a45910,a45912,
a45914,a45916,a45918,a45920,a45922,a45924,a45926,a45928,a45930,a45932,a45934,a45936,a45938,a45940,a45942,
a45944,a45946,a45948,a45950,a45952,a45954,a45956,a45958,a45960,a45962,a45964,a45966,a45968,a45970,a45972,
a45974,a45976,a45978,a45980,a45982,a45984,a45986,a45988,a45990,a45992,a45994,a45996,a45998,a46000,a46002,
a46004,a46006,a46008,a46010,a46012,a46014,a46016,a46018,a46020,a46022,a46024,a46026,a46028,a46030,a46032,
a46034,a46036,a46038,a46040,a46042,a46044,a46046,a46048,a46050,a46052,a46054,a46056,a46058,a46060,a46062,
a46064,a46066,a46068,a46070,a46072,a46074,a46076,a46078,a46080,a46082,a46084,a46086,a46088,a46090,a46092,
a46094,a46096,a46098,a46100,a46102,a46104,a46106,a46108,a46110,a46112,a46114,a46116,a46118,a46120,a46122,
a46124,a46126,a46128,a46130,a46132,a46134,a46136,a46138,a46140,a46142,a46144,a46146,a46148,a46150,a46152,
a46154,a46156,a46158,a46160,a46162,a46164,a46166,a46168,a46170,a46172,a46174,a46178,a46180,a46182,a46184,
a46186,a46188,a46190,a46192,a46194,a46196,a46198,a46200,a46202,a46204,a46206,a46208,a46210,a46212,a46214,
a46216,a46218,a46220,a46222,a46224,a46226,a46228,a46230,a46232,a46234,a46236,a46238,a46240,a46242,a46244,
a46246,a46248,a46250,a46252,a46254,a46256,a46258,a46260,a46262,a46264,a46266,a46268,a46270,a46272,a46274,
a46276,a46278,a46280,a46282,a46284,a46286,a46288,a46290,a46292,a46294,a46296,a46298,a46300,a46302,a46304,
a46306,a46308,a46310,a46312,a46314,a46316,a46318,a46320,a46322,a46324,a46326,a46328,a46330,a46332,a46334,
a46336,a46338,a46340,a46342,a46344,a46346,a46348,a46350,a46352,a46354,a46356,a46358,a46360,a46362,a46364,
a46366,a46368,a46370,a46372,a46374,a46376,a46378,a46380,a46382,a46384,a46386,a46388,a46390,a46392,a46394,
a46396,a46398,a46400,a46402,a46404,a46406,a46408,a46410,a46412,a46414,a46416,a46418,a46420,a46422,a46424,
a46426,a46428,a46430,a46432,a46434,a46436,a46438,a46440,a46442,a46444,a46446,a46448,a46450,a46452,a46454,
a46456,a46458,a46460,a46462,a46464,a46466,a46468,a46470,a46472,a46474,a46476,a46478,a46480,a46482,a46484,
a46486,a46488,a46490,a46492,a46494,a46496,a46498,a46500,a46502,a46504,a46506,a46508,a46510,a46512,a46514,
a46516,a46518,a46520,a46522,a46524,a46526,a46528,a46530,a46532,a46534,a46536,a46538,a46540,a46542,a46544,
a46546,a46548,a46550,a46552,a46554,a46556,a46558,a46560,a46562,a46564,a46566,a46568,a46570,a46572,a46574,
a46576,a46578,a46580,a46582,a46584,a46586,a46588,a46590,a46592,a46594,a46596,a46598,a46600,a46602,a46604,
a46606,a46608,a46610,a46612,a46614,a46616,a46618,a46620,a46622,a46624,a46626,a46628,a46630,a46632,a46634,
a46636,a46638,a46640,a46642,a46644,a46646,a46648,a46650,a46652,a46654,a46656,a46658,a46660,a46662,a46664,
a46666,a46668,a46670,a46672,a46674,a46676,a46678,a46680,a46682,a46684,a46686,a46688,a46690,a46692,a46694,
a46696,a46698,a46700,a46702,a46704,a46706,a46708,a46710,a46712,a46714,a46716,a46718,a46720,a46722,a46724,
a46726,a46728,a46730,a46732,a46734,a46736,a46738,a46740,a46742,a46744,a46746,a46748,a46750,a46752,a46754,
a46756,a46758,a46760,a46762,a46764,a46766,a46768,a46770,a46772,a46774,a46776,a46778,a46780,a46782,a46784,
a46786,a46788,a46790,a46792,a46794,a46796,a46798,a46800,a46802,a46804,a46806,a46808,a46810,a46812,a46814,
a46816,a46818,a46820,a46822,a46824,a46826,a46828,a46830,a46832,a46834,a46836,a46838,a46840,a46842,a46844,
a46846,a46848,a46850,a46852,a46854,a46856,a46858,a46860,a46862,a46864,a46866,a46868,a46870,a46872,a46874,
a46876,a46878,a46880,a46882,a46884,a46886,a46888,a46890,a46892,a46894,a46896,a46898,a46900,a46902,a46904,
a46906,a46908,a46910,a46912,a46914,a46916,a46918,a46920,a46922,a46924,a46926,a46928,a46930,a46932,a46934,
a46936,a46938,a46940,a46942,a46944,a46946,a46948,a46950,a46952,a46954,a46956,a46958,a46960,a46962,a46964,
a46966,a46968,a46970,a46972,a46974,a46976,a46978,a46980,a46982,a46984,a46986,a46988,a46990,a46992,a46994,
a46996,a46998,a47000,a47002,a47004,a47006,a47008,a47010,a47012,a47014,a47016,a47018,a47020,a47022,a47024,
a47026,a47028,a47030,a47032,a47034,a47036,a47038,a47040,a47042,a47044,a47046,a47048,a47050,a47052,a47054,
a47056,a47058,a47060,a47062,a47064,a47066,a47068,a47070,a47072,a47074,a47076,a47078,a47080,a47082,a47084,
a47086,a47088,a47090,a47092,a47094,a47096,a47098,a47100,a47102,a47104,a47106,a47108,a47110,a47112,a47114,
a47116,a47118,a47120,a47122,a47124,a47126,a47128,a47130,a47132,a47134,a47136,a47138,a47140,a47142,a47144,
a47146,a47148,a47150,a47152,a47154,a47156,a47158,a47160,a47162,a47164,a47166,a47168,a47170,a47172,a47174,
a47176,a47178,a47180,a47182,a47184,a47186,a47188,a47190,a47192,a47194,a47196,a47198,a47200,a47202,a47204,
a47206,a47208,a47210,a47212,a47214,a47216,a47218,a47220,a47222,a47224,a47226,a47228,a47230,a47232,a47234,
a47236,a47238,a47240,a47242,a47244,a47246,a47248,a47250,a47252,a47254,a47256,a47258,a47260,a47262,a47264,
a47266,a47268,a47270,a47272,a47274,a47276,a47278,a47280,a47282,a47284,a47286,a47288,a47290,a47292,a47294,
a47296,a47298,a47300,a47302,a47304,a47306,a47308,a47310,a47312,a47314,a47316,a47318,a47320,a47322,a47324,
a47326,a47328,a47330,a47332,a47334,a47336,a47338,a47340,a47342,a47344,a47346,a47348,a47350,a47352,a47354,
a47356,a47358,a47360,a47362,a47364,a47366,a47368,a47370,a47372,a47374,a47376,a47378,a47380,a47382,a47384,
a47386,a47388,a47390,a47392,a47394,a47396,a47398,a47400,a47402,a47404,a47406,a47408,a47410,a47412,a47414,
a47416,a47418,a47420,a47422,a47424,a47426,a47428,a47430,a47432,a47434,a47436,a47438,a47440,a47442,a47444,
a47446,a47448,a47450,a47452,a47454,a47456,a47458,a47460,a47462,a47464,a47466,a47468,a47470,a47472,a47474,
a47476,a47478,a47480,a47482,a47484,a47486,a47488,a47490,a47492,a47494,a47496,a47498,a47500,a47502,a47504,
a47506,a47508,a47510,a47512,a47514,a47516,a47518,a47520,a47522,a47524,a47526,a47528,a47530,a47532,a47534,
a47536,a47538,a47540,a47542,a47544,a47546,a47548,a47550,a47552,a47554,a47556,a47558,a47560,a47562,a47564,
a47566,a47568,a47570,a47572,a47574,a47576,a47578,a47580,a47582,a47584,a47586,a47588,a47590,a47592,a47594,
a47596,a47598,a47600,a47602,a47604,a47606,a47608,a47610,a47612,a47614,a47616,a47618,a47620,a47622,a47624,
a47626,a47628,a47630,a47632,a47634,a47636,a47638,a47640,a47642,a47644,a47646,a47648,a47650,a47652,a47654,
a47656,a47658,a47660,a47662,a47664,a47666,a47668,a47670,a47672,a47674,a47676,a47678,a47680,a47682,a47684,
a47686,a47688,a47690,a47692,a47694,a47696,a47698,a47700,a47702,a47704,a47706,a47708,a47710,a47712,a47714,
a47716,a47718,a47720,a47722,a47724,a47726,a47728,a47730,a47732,a47734,a47736,a47738,a47740,a47742,a47744,
a47746,a47748,a47750,a47752,a47754,a47756,a47758,a47760,a47762,a47764,a47766,a47768,a47770,a47772,a47774,
a47776,a47778,a47780,a47782,a47784,a47786,a47788,a47790,a47792,a47794,a47796,a47798,a47800,a47802,a47804,
a47806,a47808,a47810,a47812,a47814,a47816,a47818,a47820,a47822,a47824,a47826,a47828,a47830,a47832,a47834,
a47836,a47838,a47840,a47842,a47844,a47846,a47848,a47850,a47852,a47854,a47856,a47858,a47860,a47862,a47864,
a47866,a47868,a47870,a47872,a47874,a47876,a47878,a47880,a47882,a47884,a47886,a47888,a47890,a47892,a47894,
a47896,a47898,a47900,a47902,a47904,a47906,a47908,a47910,a47912,a47914,a47916,a47918,a47920,a47922,a47924,
a47926,a47928,a47930,a47932,a47934,a47936,a47938,a47940,a47942,a47944,a47946,a47948,a47950,a47952,a47954,
a47956,a47958,a47960,a47962,a47964,a47966,a47968,a47970,a47972,a47974,a47976,a47978,a47980,a47982,a47984,
a47986,a47988,a47990,a47992,a47994,a47996,a47998,a48000,a48002,a48004,a48006,a48008,a48010,a48012,a48014,
a48016,a48018,a48020,a48024,a48026,a48028,a48030,a48032,a48036,a48038,a48040,a48042,a48044,a48046,a48050,
a48052,a48054,a48056,a48058,a48060,a48062,a48064,a48066,a48068,a48070,a48072,a48074,a48076,a48078,a48080,
a48082,a48084,a48086,a48088,a48090,a48092,a48094,a48096,a48098,a48100,a48102,a48104,a48106,a48108,a48110,
a48112,a48114,a48116,a48118,a48120,a48122,a48124,a48126,a48128,a48130,a48132,a48134,a48136,a48138,a48140,
a48142,a48144,a48146,a48148,a48150,a48152,a48154,a48156,a48158,a48160,a48162,a48164,a48166,a48168,a48170,
a48172,a48174,a48176,a48178,a48180,a48182,a48184,a48186,a48188,a48190,a48192,a48194,a48196,a48198,a48200,
a48202,a48204,a48206,a48208,a48210,a48212,a48214,a48216,a48218,a48220,a48222,a48224,a48226,a48228,a48230,
a48232,a48234,a48236,a48238,a48240,a48242,a48244,a48246,a48248,a48250,a48252,a48254,a48256,a48258,a48260,
a48262,a48264,a48266,a48268,a48270,a48272,a48274,a48276,a48278,a48280,a48282,a48284,a48286,a48288,a48290,
a48292,a48294,a48296,a48298,a48300,a48302,a48304,a48306,a48308,a48310,a48312,a48314,a48316,a48318,a48320,
a48322,a48324,a48326,a48328,a48330,a48332,a48334,a48336,a48338,a48340,a48342,a48344,a48346,a48348,a48350,
a48352,a48354,a48356,a48358,a48360,a48362,a48364,a48366,a48368,a48370,a48372,a48374,a48376,a48378,a48380,
a48382,a48384,a48386,a48388,a48390,a48392,a48394,a48396,a48398,a48400,a48402,a48404,a48406,a48408,a48410,
a48412,a48414,a48416,a48418,a48420,a48422,a48424,a48426,a48428,a48430,a48432,a48434,a48436,a48438,a48440,
a48442,a48444,a48446,a48448,a48450,a48452,a48454,a48456,a48458,a48460,a48462,a48464,a48466,a48468,a48470,
a48472,a48474,a48476,a48478,a48480,a48482,a48484,a48486,a48488,a48490,a48492,a48494,a48496,a48498,a48500,
a48502,a48504,a48506,a48508,a48510,a48512,a48514,a48516,a48518,a48520,a48522,a48524,a48526,a48528,a48530,
a48532,a48534,a48536,a48538,a48540,a48542,a48544,a48546,a48548,a48550,a48552,a48554,a48556,a48558,a48560,
a48562,a48564,a48566,a48568,a48570,a48572,a48574,a48576,a48578,a48580,a48582,a48586,a48588,a48592,a48594,
a48598,a48600,a48604,a48606,a48610,a48612,a48616,a48618,a48622,a48624,a48628,a48630,a48634,a48636,a48640,
a48642,a48646,a48648,a48652,a48654,a48658,a48660,a48664,a48666,a48670,a48672,a48676,a48678,a48682,a48684,
a48688,a48690,a48694,a48696,a48700,a48702,a48706,a48708,a48710,a48712,a48714,a48716,a48718,a48720,a48722,
a48724,a48726,a48730,a48732,a48734,a48736,a48738,a48740,a48742,a48744,a48746,a48748,a48750,a48752,a48754,
a48756,a48758,a48760,a48762,a48764,a48766,a48768,a48770,a48772,a48774,a48776,a48778,a48780,a48782,a48784,
a48786,a48788,a48790,a48794,a48796,a48798,a48800,a48802,a48804,a48806,a48810,a48812,a48814,a48816,a48818,
a48820,a48822,a48824,a48826,a48828,a48830,a48832,a48834,a48836,a48838,a48840,a48842,a48844,a48846,a48848,
a48850,a48852,a48854,a48856,a48858,a48860,a48862,a48864,a48866,a48868,a48870,a48872,a48874,a48876,a48878,
a48880,a48882,a48884,a48886,a48888,a48890,a48892,a48894,a48896,a48898,a48900,a48902,a48904,a48906,a48908,
a48910,a48912,a48914,a48916,a48918,a48920,a48922,a48924,a48926,a48928,a48930,a48932,a48934,a48936,a48938,
a48940,a48942,a48944,a48946,a48948,a48950,a48952,a48954,a48956,a48958,a48960,a48962,a48964,a48966,a48968,
a48970,a48972,a48974,a48976,a48978,a48980,a48982,a48984,a48986,a48988,a48990,a48992,a48994,a48996,a48998,
a49000,a49002,a49004,a49006,a49008,a49010,a49012,a49014,a49016,a49018,a49020,a49022,a49024,a49026,a49028,
a49030,a49032,a49034,a49036,a49038,a49040,a49042,a49044,a49046,a49048,a49050,a49052,a49054,a49056,a49058,
a49060,a49062,a49064,a49066,a49068,a49070,a49072,a49074,a49076,a49078,a49080,a49082,a49084,a49086,a49088,
a49090,a49092,a49094,a49096,a49098,a49100,a49102,a49104,a49106,a49108,a49110,a49112,a49114,a49116,a49118,
a49120,a49122,a49124,a49126,a49128,a49130,a49132,a49134,a49136,a49138,a49140,a49142,a49144,a49146,a49148,
a49150,a49152,a49154,a49156,a49158,a49160,a49162,a49164,a49166,a49168,a49170,a49172,a49174,a49176,a49178,
a49180,a49182,a49184,a49186,a49188,a49190,a49192,a49194,a49196,a49198,a49200,a49202,a49204,a49206,a49208,
a49210,a49212,a49214,a49216,a49218,a49220,a49222,a49224,a49226,a49228,a49230,a49232,a49234,a49236,a49238,
a49240,a49242,a49244,a49246,a49248,a49250,a49252,a49254,a49256,a49258,a49260,a49262,a49264,a49266,a49268,
a49270,a49272,a49274,a49276,a49278,a49280,a49282,a49284,a49286,a49288,a49290,a49292,a49294,a49296,a49298,
a49300,a49302,a49304,a49306,a49308,a49310,a49312,a49314,a49316,a49318,a49320,a49322,a49324,a49326,a49328,
a49330,a49332,a49334,a49336,a49338,a49340,a49342,a49344,a49346,a49348,a49350,a49352,a49354,a49356,a49358,
a49360,a49362,a49364,a49366,a49368,a49370,a49372,a49374,a49376,a49378,a49380,a49382,a49384,a49386,a49388,
a49390,a49392,a49394,a49396,a49398,a49400,a49402,a49404,a49406,a49408,a49410,a49412,a49414,a49416,a49418,
a49420,a49422,a49424,a49426,a49428,a49430,a49432,a49434,a49436,a49438,a49440,a49442,a49444,a49446,a49448,
a49450,a49452,a49454,a49456,a49458,a49460,a49462,a49464,a49466,a49468,a49470,a49472,a49474,a49476,a49478,
a49480,a49482,a49484,a49486,a49488,a49490,a49492,a49494,a49496,a49498,a49500,a49502,a49504,a49506,a49508,
a49510,a49512,a49514,a49516,a49518,a49520,a49522,a49524,a49526,a49528,a49530,a49532,a49534,a49536,a49538,
a49540,a49542,a49544,a49546,a49548,a49550,a49552,a49554,a49556,a49558,a49560,a49562,a49564,a49566,a49568,
a49570,a49572,a49574,a49576,a49578,a49580,a49582,a49584,a49586,a49588,a49590,a49592,a49594,a49596,a49598,
a49600,a49602,a49604,a49606,a49608,a49610,a49612,a49614,a49616,a49618,a49620,a49622,a49624,a49626,a49628,
a49630,a49632,a49634,a49636,a49638,a49640,a49642,a49644,a49646,a49648,a49650,a49652,a49654,a49656,a49658,
a49660,a49662,a49664,a49666,a49668,a49670,a49672,a49674,a49676,a49678,a49680,a49682,a49684,a49686,a49688,
a49690,a49692,a49694,a49696,a49698,a49700,a49702,a49704,a49706,a49708,a49710,a49712,a49714,a49716,a49718,
a49720,a49722,a49724,a49726,a49728,a49730,a49732,a49734,a49736,a49738,a49742,a49744,a49746,a49748,a49750,
a49752,a49754,a49756,a49760,a49762,a49764,a49766,a49768,a49770,a49772,a49774,a49776,a49778,a49780,a49782,
a49786,a49788,a49790,a49792,a49794,a49796,a49798,a49800,a49804,a49806,a49808,a49810,a49812,a49814,a49816,
a49818,a49820,a49822,a49826,a49828,a49830,a49832,a49834,a49836,a49838,a49840,a49844,a49846,a49848,a49850,
a49852,a49854,a49856,a49858,a49860,a49864,a49866,a49868,a49870,a49872,a49874,a49876,a49878,a49882,a49884,
a49886,a49888,a49890,a49892,a49894,a49896,a49898,a49900,a49902,a49904,a49906,a49908,a49910,a49912,a49914,
a49916,a49918,a49920,a49922,a49924,a49926,a49928,a49930,a49934,a49936,a49938,a49940,a49942,a49944,a49946,
a49948,a49950,a49952,a49954,a49956,a49958,a49960,a49962,a49964,a49966,a49968,a49970,a49972,a49974,a49976,
a49978,a49980,a49982,a49984,a49986,a49988,a49990,a49992,a49994,a49998,a50000,a50002,a50004,a50006,a50008,
a50010,a50012,a50014,a50016,a50018,a50020,a50022,a50026,a50028,a50030,a50032,a50034,a50036,a50038,a50040,
a50042,a50044,a50046,a50048,a50050,a50052,a50054,a50056,a50058,a50060,a50062,a50064,a50068,a50070,a50072,
a50074,a50076,a50078,a50080,a50082,a50086,a50088,a50090,a50092,a50094,a50096,a50098,a50100,a50102,a50104,
a50106,a50108,a50110,a50112,a50116,a50118,a50120,a50122,a50124,a50126,a50128,a50130,a50132,a50134,a50138,
a50140,a50142,a50144,a50146,a50148,a50150,a50152,a50154,a50156,a50158,a50160,a50162,a50166,a50168,a50170,
a50172,a50174,a50178,a50180,a50182,a50184,a50186,a50188,a50190,a50192,a50194,a50196,a50198,a50200,a50202,
a50204,a50206,a50208,a50210,a50212,a50214,a50216,a50218,a50220,a50222,a50224,a50226,a50228,a50230,a50232,
a50234,a50236,a50238,a50240,a50242,a50244,a50246,a50248,a50250,a50252,a50254,a50256,a50258,a50260,a50262,
a50264,a50266,a50268,a50270,a50272,a50274,a50276,a50278,a50280,a50282,a50284,a50286,a50288,a50290,a50292,
a50294,a50296,a50298,a50300,a50302,a50304,a50306,a50308,a50310,a50312,a50314,a50316,a50318,a50320,a50322,
a50324,a50326,a50328,a50330,a50332,a50334,a50336,a50338,a50340,a50342,a50344,a50348,a50350,a50352,a50354,
a50356,a50358,a50360,a50362,a50364,a50366,a50368,a50370,a50372,a50374,a50376,a50378,a50380,a50382,a50384,
a50386,a50388,a50390,a50392,a50394,a50396,a50398,a50400,a50402,a50404,a50406,a50408,a50410,a50412,a50414,
a50416,a50418,a50422,a50424,a50426,a50428,a50430,a50432,a50434,a50436,a50438,a50440,a50442,a50444,a50446,
a50448,a50450,a50452,a50454,a50456,a50458,a50460,a50462,a50464,a50466,a50468,a50470,a50472,a50474,a50476,
a50478,a50480,a50482,a50484,a50486,a50488,a50490,a50492,a50494,a50496,a50498,a50500,a50502,a50504,a50506,
a50508,a50510,a50512,a50514,a50516,a50518,a50520,a50522,a50524,a50526,a50528,a50530,a50532,a50534,a50536,
a50538,a50540,a50542,a50544,a50546,a50548,a50550,a50552,a50554,a50556,a50558,a50560,a50562,a50564,a50566,
a50568,a50570,a50572,a50574,a50576,a50578,a50580,a50582,a50584,a50586,a50588,a50590,a50592,a50594,a50596,
a50598,a50600,a50602,a50604,a50606,a50608,a50610,a50612,a50614,a50616,a50618,a50622,a50624,a50626,a50628,
a50630,a50632,a50634,a50636,a50638,a50640,a50642,a50644,a50648,a50650,a50652,a50654,a50656,a50658,a50660,
a50662,a50664,a50666,a50668,a50670,a50674,a50676,a50678,a50680,a50682,a50684,a50686,a50688,a50690,a50692,
a50694,a50696,a50700,a50702,a50704,a50706,a50708,a50710,a50712,a50714,a50716,a50718,a50720,a50722,a50726,
a50728,a50730,a50732,a50734,a50736,a50738,a50740,a50742,a50744,a50746,a50748,a50752,a50754,a50756,a50758,
a50760,a50762,a50764,a50766,a50768,a50770,a50772,a50774,a50778,a50780,a50782,a50784,a50786,a50788,a50790,
a50792,a50794,a50796,a50798,a50800,a50804,a50806,a50808,a50810,a50812,a50814,a50816,a50818,a50820,a50822,
a50824,a50826,a50830,a50832,a50834,a50836,a50838,a50840,a50842,a50844,a50846,a50848,a50850,a50852,a50856,
a50858,a50860,a50862,a50864,a50866,a50868,a50870,a50872,a50874,a50876,a50878,a50880,a50882,a50884,a50886,
a50888,a50890,a50892,a50894,a50896,a50898,a50900,a50902,a50904,a50906,a50908,a50910,a50912,a50914,a50916,
a50918,a50920,a50922,a50924,a50926,a50928,a50930,a50932,a50934,a50936,a50938,a50940,a50942,a50944,a50946,
a50948,a50950,a50952,a50954,a50956,a50958,a50960,a50962,a50964,a50966,a50968,a50970,a50974,a50976,a50978,
a50980,a50982,a50984,a50988,a50992,a50994,a50996,a50998,a51002,a51004,a51006,a51008,a51010,a51012,a51014,
a51016,a51018,a51020,a51022,a51024,a51026,a51028,a51030,a51032,a51034,a51036,a51038,a51040,a51042,a51044,
a51046,a51048,a51050,a51052,a51054,a51056,a51058,a51060,a51062,a51064,a51066,a51068,a51070,a51072,a51074,
a51076,a51078,a51080,a51082,a51084,a51086,a51088,a51090,a51092,a51094,a51096,a51098,a51100,p0;

reg l880,l882,l884,l886,l888,l890,l892,l894,l896,l898,l900,l902,l904,l906,l908,
l910,l912,l914,l916,l918,l920,l922,l924,l926,l928,l930,l932,l934,l936,l938,
l940,l942,l944,l946,l948,l950,l952,l954,l956,l958,l960,l962,l964,l966,l968,
l970,l972,l974,l976,l978,l980,l982,l984,l986,l988,l990,l992,l994,l996,l998,
l1000,l1002,l1004,l1006,l1008,l1010,l1012,l1014,l1016,l1018,l1020,l1022,l1024,l1026,l1028,
l1030,l1032,l1034,l1036,l1038,l1040,l1042,l1044,l1046,l1048,l1050,l1052,l1054,l1056,l1058,
l1060,l1062,l1064,l1066,l1068,l1070,l1072,l1074,l1076,l1078,l1080,l1082,l1084,l1086,l1088,
l1090,l1092,l1094,l1096,l1098,l1100,l1102,l1104,l1106,l1108,l1110,l1112,l1114,l1116,l1118,
l1120,l1122,l1124,l1126,l1128,l1130,l1132,l1134,l1136,l1138,l1140,l1142,l1144,l1146,l1148,
l1150,l1152,l1154,l1156,l1158,l1160,l1162,l1164,l1166,l1168,l1170,l1172,l1174,l1176,l1178,
l1180,l1182,l1184,l1186,l1188,l1190,l1192,l1194,l1196,l1198,l1200,l1202,l1204,l1206,l1208,
l1210,l1212,l1214,l1216,l1218,l1220,l1222,l1224,l1226,l1228,l1230,l1232,l1234,l1236,l1238,
l1240,l1242,l1244,l1246,l1248,l1250,l1252,l1254,l1256,l1258,l1260,l1262,l1264,l1266,l1268,
l1270,l1272,l1274,l1276,l1278,l1280,l1282,l1284,l1286,l1288,l1290,l1292,l1294,l1296,l1298,
l1300,l1302,l1304,l1306,l1308,l1310,l1312,l1314,l1316,l1318,l1320,l1322,l1324,l1326,l1328,
l1330,l1332,l1334,l1336,l1338,l1340,l1342,l1344,l1346,l1348,l1350,l1352,l1354,l1356,l1358,
l1360,l1362,l1364,l1366,l1368,l1370,l1372,l1374,l1376,l1378,l1380,l1382,l1384,l1386,l1388,
l1390,l1392,l1394,l1396,l1398,l1400,l1402,l1404,l1406,l1408,l1410,l1412,l1414,l1416,l1418,
l1420,l1422,l1424,l1426,l1428,l1430,l1432,l1434,l1436,l1438,l1440,l1442,l1444,l1446,l1448,
l1450,l1452,l1454,l1456,l1458,l1460,l1462,l1464,l1466,l1468,l1470,l1472,l1474,l1476,l1478,
l1480,l1482,l1484,l1486,l1488,l1490,l1492,l1494,l1496,l1498,l1500,l1502,l1504,l1506,l1508,
l1510,l1512,l1514,l1516,l1518,l1520,l1522,l1524,l1526,l1528,l1530,l1532,l1534,l1536,l1538,
l1540,l1542,l1544,l1546,l1548,l1550,l1552,l1554,l1556,l1558,l1560,l1562,l1564,l1566,l1568,
l1570,l1572,l1574,l1576,l1578,l1580,l1582,l1584,l1586,l1588,l1590,l1592,l1594,l1596,l1598,
l1600,l1602,l1604,l1606,l1608,l1610,l1612,l1614,l1616,l1618,l1620,l1622,l1624,l1626,l1628,
l1630,l1632,l1634,l1636,l1638,l1640,l1642,l1644,l1646,l1648,l1650,l1652,l1654,l1656,l1658,
l1660,l1662,l1664,l1666,l1668,l1670,l1672,l1674,l1676,l1678,l1680,l1682,l1684,l1686,l1688,
l1690,l1692,l1694,l1696,l1698,l1700,l1702,l1704,l1706,l1708,l1710,l1712,l1714,l1716,l1718,
l1720,l1722,l1724,l1726,l1728,l1730,l1732,l1734,l1736,l1738,l1740,l1742,l1744,l1746,l1748,
l1750,l1752,l1754,l1756,l1758,l1760,l1762,l1764,l1766,l1768,l1770,l1772,l1774,l1776,l1778,
l1780,l1782,l1784,l1786,l1788,l1790,l1792,l1794,l1796,l1798,l1800,l1802,l1804,l1806,l1808,
l1810,l1812,l1814,l1816,l1818,l1820,l1822,l1824,l1826,l1828,l1830,l1832,l1834,l1836,l1838,
l1840,l1842,l1844,l1846,l1848,l1850,l1852,l1854,l1856,l1858,l1860,l1862,l1864,l1866,l1868,
l1870,l1872,l1874,l1876,l1878,l1880,l1882,l1884,l1886,l1888,l1890,l1892,l1894,l1896,l1898,
l1900,l1902,l1904,l1906,l1908,l1910,l1912,l1914,l1916,l1918,l1920,l1922,l1924,l1926,l1928,
l1930,l1932,l1934,l1936,l1938,l1940,l1942,l1944,l1946,l1948,l1950,l1952,l1954,l1956,l1958,
l1960,l1962,l1964,l1966,l1968,l1970,l1972,l1974,l1976,l1978,l1980,l1982,l1984,l1986,l1988,
l1990,l1992,l1994,l1996,l1998,l2000,l2002,l2004,l2006,l2008,l2010,l2012,l2014,l2016,l2018,
l2020,l2022,l2024,l2026,l2028,l2030,l2032,l2034,l2036,l2038,l2040,l2042,l2044,l2046,l2048,
l2050,l2052,l2054,l2056,l2058,l2060,l2062,l2064,l2066,l2068,l2070,l2072,l2074,l2076,l2078,
l2080,l2082,l2084,l2086,l2088,l2090,l2092,l2094,l2096,l2098,l2100,l2102,l2104,l2106,l2108,
l2110,l2112,l2114,l2116,l2118,l2120,l2122,l2124,l2126,l2128,l2130,l2132,l2134,l2136,l2138,
l2140,l2142,l2144,l2146,l2148,l2150,l2152,l2154,l2156,l2158,l2160,l2162,l2164,l2166,l2168,
l2170,l2172,l2174,l2176,l2178,l2180,l2182,l2184,l2186,l2188,l2190,l2192,l2194,l2196,l2198,
l2200,l2202,l2204,l2206,l2208,l2210,l2212,l2214,l2216,l2218,l2220,l2222,l2224,l2226,l2228,
l2230,l2232,l2234,l2236,l2238,l2240,l2242,l2244,l2246,l2248,l2250,l2252,l2254,l2256,l2258,
l2260,l2262,l2264,l2266,l2268,l2270,l2272,l2274,l2276,l2278,l2280,l2282,l2284,l2286,l2288,
l2290,l2292,l2294,l2296,l2298,l2300,l2302,l2304,l2306,l2308,l2310,l2312,l2314,l2316,l2318,
l2320,l2322,l2324,l2326,l2328,l2330,l2332,l2334,l2336,l2338,l2340,l2342,l2344,l2346,l2348,
l2350,l2352,l2354,l2356,l2358,l2360,l2362,l2364,l2366,l2368,l2370,l2372,l2374,l2376,l2378,
l2380,l2382,l2384,l2386,l2388,l2390,l2392,l2394,l2396,l2398,l2400,l2402,l2404,l2406,l2408,
l2410,l2412,l2414,l2416,l2418,l2420,l2422,l2424,l2426,l2428,l2430,l2432,l2434,l2436,l2438,
l2440,l2442,l2444,l2446,l2448,l2450,l2452,l2454,l2456,l2458,l2460,l2462,l2464,l2466,l2468,
l2470,l2472,l2474,l2476,l2478,l2480,l2482,l2484,l2486,l2488,l2490,l2492,l2494,l2496,l2498,
l2500;

initial
begin
   l880 = 0;
   l882 = 0;
   l884 = 0;
   l886 = 0;
   l888 = 0;
   l890 = 0;
   l892 = 0;
   l894 = 0;
   l896 = 0;
   l898 = 0;
   l900 = 0;
   l902 = 0;
   l904 = 0;
   l906 = 0;
   l908 = 0;
   l910 = 0;
   l912 = 0;
   l914 = 0;
   l916 = 0;
   l918 = 0;
   l920 = 0;
   l922 = 0;
   l924 = 0;
   l926 = 0;
   l928 = 0;
   l930 = 0;
   l932 = 0;
   l934 = 0;
   l936 = 0;
   l938 = 0;
   l940 = 0;
   l942 = 0;
   l944 = 0;
   l946 = 0;
   l948 = 0;
   l950 = 0;
   l952 = 0;
   l954 = 0;
   l956 = 0;
   l958 = 0;
   l960 = 0;
   l962 = 0;
   l964 = 0;
   l966 = 0;
   l968 = 0;
   l970 = 0;
   l972 = 0;
   l974 = 0;
   l976 = 0;
   l978 = 0;
   l980 = 0;
   l982 = 0;
   l984 = 0;
   l986 = 0;
   l988 = 0;
   l990 = 0;
   l992 = 0;
   l994 = 0;
   l996 = 0;
   l998 = 0;
   l1000 = 0;
   l1002 = 0;
   l1004 = 0;
   l1006 = 0;
   l1008 = 0;
   l1010 = 0;
   l1012 = 0;
   l1014 = 0;
   l1016 = 0;
   l1018 = 0;
   l1020 = 0;
   l1022 = 0;
   l1024 = 0;
   l1026 = 0;
   l1028 = 0;
   l1030 = 0;
   l1032 = 0;
   l1034 = 0;
   l1036 = 0;
   l1038 = 0;
   l1040 = 0;
   l1042 = 0;
   l1044 = 0;
   l1046 = 0;
   l1048 = 0;
   l1050 = 0;
   l1052 = 0;
   l1054 = 0;
   l1056 = 0;
   l1058 = 0;
   l1060 = 0;
   l1062 = 0;
   l1064 = 0;
   l1066 = 0;
   l1068 = 0;
   l1070 = 0;
   l1072 = 0;
   l1074 = 0;
   l1076 = 0;
   l1078 = 0;
   l1080 = 0;
   l1082 = 0;
   l1084 = 0;
   l1086 = 0;
   l1088 = 0;
   l1090 = 0;
   l1092 = 0;
   l1094 = 0;
   l1096 = 0;
   l1098 = 0;
   l1100 = 0;
   l1102 = 0;
   l1104 = 0;
   l1106 = 0;
   l1108 = 0;
   l1110 = 0;
   l1112 = 0;
   l1114 = 0;
   l1116 = 0;
   l1118 = 0;
   l1120 = 0;
   l1122 = 0;
   l1124 = 0;
   l1126 = 0;
   l1128 = 0;
   l1130 = 0;
   l1132 = 0;
   l1134 = 0;
   l1136 = 0;
   l1138 = 0;
   l1140 = 0;
   l1142 = 0;
   l1144 = 0;
   l1146 = 0;
   l1148 = 0;
   l1150 = 0;
   l1152 = 0;
   l1154 = 0;
   l1156 = 0;
   l1158 = 0;
   l1160 = 0;
   l1162 = 0;
   l1164 = 0;
   l1166 = 0;
   l1168 = 0;
   l1170 = 0;
   l1172 = 0;
   l1174 = 0;
   l1176 = 0;
   l1178 = 0;
   l1180 = 0;
   l1182 = 0;
   l1184 = 0;
   l1186 = 0;
   l1188 = 0;
   l1190 = 0;
   l1192 = 0;
   l1194 = 0;
   l1196 = 0;
   l1198 = 0;
   l1200 = 0;
   l1202 = 0;
   l1204 = 0;
   l1206 = 0;
   l1208 = 0;
   l1210 = 0;
   l1212 = 0;
   l1214 = 0;
   l1216 = 0;
   l1218 = 0;
   l1220 = 0;
   l1222 = 0;
   l1224 = 0;
   l1226 = 0;
   l1228 = 0;
   l1230 = 0;
   l1232 = 0;
   l1234 = 0;
   l1236 = 0;
   l1238 = 0;
   l1240 = 0;
   l1242 = 0;
   l1244 = 0;
   l1246 = 0;
   l1248 = 0;
   l1250 = 0;
   l1252 = 0;
   l1254 = 0;
   l1256 = 0;
   l1258 = 0;
   l1260 = 0;
   l1262 = 0;
   l1264 = 0;
   l1266 = 0;
   l1268 = 0;
   l1270 = 0;
   l1272 = 0;
   l1274 = 0;
   l1276 = 0;
   l1278 = 0;
   l1280 = 0;
   l1282 = 0;
   l1284 = 0;
   l1286 = 0;
   l1288 = 0;
   l1290 = 0;
   l1292 = 0;
   l1294 = 0;
   l1296 = 0;
   l1298 = 0;
   l1300 = 0;
   l1302 = 0;
   l1304 = 0;
   l1306 = 0;
   l1308 = 0;
   l1310 = 0;
   l1312 = 0;
   l1314 = 0;
   l1316 = 0;
   l1318 = 0;
   l1320 = 0;
   l1322 = 0;
   l1324 = 0;
   l1326 = 0;
   l1328 = 0;
   l1330 = 0;
   l1332 = 0;
   l1334 = 0;
   l1336 = 0;
   l1338 = 0;
   l1340 = 0;
   l1342 = 0;
   l1344 = 0;
   l1346 = 0;
   l1348 = 0;
   l1350 = 0;
   l1352 = 0;
   l1354 = 0;
   l1356 = 0;
   l1358 = 0;
   l1360 = 0;
   l1362 = 0;
   l1364 = 0;
   l1366 = 0;
   l1368 = 0;
   l1370 = 0;
   l1372 = 0;
   l1374 = 0;
   l1376 = 0;
   l1378 = 0;
   l1380 = 0;
   l1382 = 0;
   l1384 = 0;
   l1386 = 0;
   l1388 = 0;
   l1390 = 0;
   l1392 = 0;
   l1394 = 0;
   l1396 = 0;
   l1398 = 0;
   l1400 = 0;
   l1402 = 0;
   l1404 = 0;
   l1406 = 0;
   l1408 = 0;
   l1410 = 0;
   l1412 = 0;
   l1414 = 0;
   l1416 = 0;
   l1418 = 0;
   l1420 = 0;
   l1422 = 0;
   l1424 = 0;
   l1426 = 0;
   l1428 = 0;
   l1430 = 0;
   l1432 = 0;
   l1434 = 0;
   l1436 = 0;
   l1438 = 0;
   l1440 = 0;
   l1442 = 0;
   l1444 = 0;
   l1446 = 0;
   l1448 = 0;
   l1450 = 0;
   l1452 = 0;
   l1454 = 0;
   l1456 = 0;
   l1458 = 0;
   l1460 = 0;
   l1462 = 0;
   l1464 = 0;
   l1466 = 0;
   l1468 = 0;
   l1470 = 0;
   l1472 = 0;
   l1474 = 0;
   l1476 = 0;
   l1478 = 0;
   l1480 = 0;
   l1482 = 0;
   l1484 = 0;
   l1486 = 0;
   l1488 = 0;
   l1490 = 0;
   l1492 = 0;
   l1494 = 0;
   l1496 = 0;
   l1498 = 0;
   l1500 = 0;
   l1502 = 0;
   l1504 = 0;
   l1506 = 0;
   l1508 = 0;
   l1510 = 0;
   l1512 = 0;
   l1514 = 0;
   l1516 = 0;
   l1518 = 0;
   l1520 = 0;
   l1522 = 0;
   l1524 = 0;
   l1526 = 0;
   l1528 = 0;
   l1530 = 0;
   l1532 = 0;
   l1534 = 0;
   l1536 = 0;
   l1538 = 0;
   l1540 = 0;
   l1542 = 0;
   l1544 = 0;
   l1546 = 0;
   l1548 = 0;
   l1550 = 0;
   l1552 = 0;
   l1554 = 0;
   l1556 = 0;
   l1558 = 0;
   l1560 = 0;
   l1562 = 0;
   l1564 = 0;
   l1566 = 0;
   l1568 = 0;
   l1570 = 0;
   l1572 = 0;
   l1574 = 0;
   l1576 = 0;
   l1578 = 0;
   l1580 = 0;
   l1582 = 0;
   l1584 = 0;
   l1586 = 0;
   l1588 = 0;
   l1590 = 0;
   l1592 = 0;
   l1594 = 0;
   l1596 = 0;
   l1598 = 0;
   l1600 = 0;
   l1602 = 0;
   l1604 = 0;
   l1606 = 0;
   l1608 = 0;
   l1610 = 0;
   l1612 = 0;
   l1614 = 0;
   l1616 = 0;
   l1618 = 0;
   l1620 = 0;
   l1622 = 0;
   l1624 = 0;
   l1626 = 0;
   l1628 = 0;
   l1630 = 0;
   l1632 = 0;
   l1634 = 0;
   l1636 = 0;
   l1638 = 0;
   l1640 = 0;
   l1642 = 0;
   l1644 = 0;
   l1646 = 0;
   l1648 = 0;
   l1650 = 0;
   l1652 = 0;
   l1654 = 0;
   l1656 = 0;
   l1658 = 0;
   l1660 = 0;
   l1662 = 0;
   l1664 = 0;
   l1666 = 0;
   l1668 = 0;
   l1670 = 0;
   l1672 = 0;
   l1674 = 0;
   l1676 = 0;
   l1678 = 0;
   l1680 = 0;
   l1682 = 0;
   l1684 = 0;
   l1686 = 0;
   l1688 = 0;
   l1690 = 0;
   l1692 = 0;
   l1694 = 0;
   l1696 = 0;
   l1698 = 0;
   l1700 = 0;
   l1702 = 0;
   l1704 = 0;
   l1706 = 0;
   l1708 = 0;
   l1710 = 0;
   l1712 = 0;
   l1714 = 0;
   l1716 = 0;
   l1718 = 0;
   l1720 = 0;
   l1722 = 0;
   l1724 = 0;
   l1726 = 0;
   l1728 = 0;
   l1730 = 0;
   l1732 = 0;
   l1734 = 0;
   l1736 = 0;
   l1738 = 0;
   l1740 = 0;
   l1742 = 0;
   l1744 = 0;
   l1746 = 0;
   l1748 = 0;
   l1750 = 0;
   l1752 = 0;
   l1754 = 0;
   l1756 = 0;
   l1758 = 0;
   l1760 = 0;
   l1762 = 0;
   l1764 = 0;
   l1766 = 0;
   l1768 = 0;
   l1770 = 0;
   l1772 = 0;
   l1774 = 0;
   l1776 = 0;
   l1778 = 0;
   l1780 = 0;
   l1782 = 0;
   l1784 = 0;
   l1786 = 0;
   l1788 = 0;
   l1790 = 0;
   l1792 = 0;
   l1794 = 0;
   l1796 = 0;
   l1798 = 0;
   l1800 = 0;
   l1802 = 0;
   l1804 = 0;
   l1806 = 0;
   l1808 = 0;
   l1810 = 0;
   l1812 = 0;
   l1814 = 0;
   l1816 = 0;
   l1818 = 0;
   l1820 = 0;
   l1822 = 0;
   l1824 = 0;
   l1826 = 0;
   l1828 = 0;
   l1830 = 0;
   l1832 = 0;
   l1834 = 0;
   l1836 = 0;
   l1838 = 0;
   l1840 = 0;
   l1842 = 0;
   l1844 = 0;
   l1846 = 0;
   l1848 = 0;
   l1850 = 0;
   l1852 = 0;
   l1854 = 0;
   l1856 = 0;
   l1858 = 0;
   l1860 = 0;
   l1862 = 0;
   l1864 = 0;
   l1866 = 0;
   l1868 = 0;
   l1870 = 0;
   l1872 = 0;
   l1874 = 0;
   l1876 = 0;
   l1878 = 0;
   l1880 = 0;
   l1882 = 0;
   l1884 = 0;
   l1886 = 0;
   l1888 = 0;
   l1890 = 0;
   l1892 = 0;
   l1894 = 0;
   l1896 = 0;
   l1898 = 0;
   l1900 = 0;
   l1902 = 0;
   l1904 = 0;
   l1906 = 0;
   l1908 = 0;
   l1910 = 0;
   l1912 = 0;
   l1914 = 0;
   l1916 = 0;
   l1918 = 0;
   l1920 = 0;
   l1922 = 0;
   l1924 = 0;
   l1926 = 0;
   l1928 = 0;
   l1930 = 0;
   l1932 = 0;
   l1934 = 0;
   l1936 = 0;
   l1938 = 0;
   l1940 = 0;
   l1942 = 0;
   l1944 = 0;
   l1946 = 0;
   l1948 = 0;
   l1950 = 0;
   l1952 = 0;
   l1954 = 0;
   l1956 = 0;
   l1958 = 0;
   l1960 = 0;
   l1962 = 0;
   l1964 = 0;
   l1966 = 0;
   l1968 = 0;
   l1970 = 0;
   l1972 = 0;
   l1974 = 0;
   l1976 = 0;
   l1978 = 0;
   l1980 = 0;
   l1982 = 0;
   l1984 = 0;
   l1986 = 0;
   l1988 = 0;
   l1990 = 0;
   l1992 = 0;
   l1994 = 0;
   l1996 = 0;
   l1998 = 0;
   l2000 = 0;
   l2002 = 0;
   l2004 = 0;
   l2006 = 0;
   l2008 = 0;
   l2010 = 0;
   l2012 = 0;
   l2014 = 0;
   l2016 = 0;
   l2018 = 0;
   l2020 = 0;
   l2022 = 0;
   l2024 = 0;
   l2026 = 0;
   l2028 = 0;
   l2030 = 0;
   l2032 = 0;
   l2034 = 0;
   l2036 = 0;
   l2038 = 0;
   l2040 = 0;
   l2042 = 0;
   l2044 = 0;
   l2046 = 0;
   l2048 = 0;
   l2050 = 0;
   l2052 = 0;
   l2054 = 0;
   l2056 = 0;
   l2058 = 0;
   l2060 = 0;
   l2062 = 0;
   l2064 = 0;
   l2066 = 0;
   l2068 = 0;
   l2070 = 0;
   l2072 = 0;
   l2074 = 0;
   l2076 = 0;
   l2078 = 0;
   l2080 = 0;
   l2082 = 0;
   l2084 = 0;
   l2086 = 0;
   l2088 = 0;
   l2090 = 0;
   l2092 = 0;
   l2094 = 0;
   l2096 = 0;
   l2098 = 0;
   l2100 = 0;
   l2102 = 0;
   l2104 = 0;
   l2106 = 0;
   l2108 = 0;
   l2110 = 0;
   l2112 = 0;
   l2114 = 0;
   l2116 = 0;
   l2118 = 0;
   l2120 = 0;
   l2122 = 0;
   l2124 = 0;
   l2126 = 0;
   l2128 = 0;
   l2130 = 0;
   l2132 = 0;
   l2134 = 0;
   l2136 = 0;
   l2138 = 0;
   l2140 = 0;
   l2142 = 0;
   l2144 = 0;
   l2146 = 0;
   l2148 = 0;
   l2150 = 0;
   l2152 = 0;
   l2154 = 0;
   l2156 = 0;
   l2158 = 0;
   l2160 = 0;
   l2162 = 0;
   l2164 = 0;
   l2166 = 0;
   l2168 = 0;
   l2170 = 0;
   l2172 = 0;
   l2174 = 0;
   l2176 = 0;
   l2178 = 0;
   l2180 = 0;
   l2182 = 0;
   l2184 = 0;
   l2186 = 0;
   l2188 = 0;
   l2190 = 0;
   l2192 = 0;
   l2194 = 0;
   l2196 = 0;
   l2198 = 0;
   l2200 = 0;
   l2202 = 0;
   l2204 = 0;
   l2206 = 0;
   l2208 = 0;
   l2210 = 0;
   l2212 = 0;
   l2214 = 0;
   l2216 = 0;
   l2218 = 0;
   l2220 = 0;
   l2222 = 0;
   l2224 = 0;
   l2226 = 0;
   l2228 = 0;
   l2230 = 0;
   l2232 = 0;
   l2234 = 0;
   l2236 = 0;
   l2238 = 0;
   l2240 = 0;
   l2242 = 0;
   l2244 = 0;
   l2246 = 0;
   l2248 = 0;
   l2250 = 0;
   l2252 = 0;
   l2254 = 0;
   l2256 = 0;
   l2258 = 0;
   l2260 = 0;
   l2262 = 0;
   l2264 = 0;
   l2266 = 0;
   l2268 = 0;
   l2270 = 0;
   l2272 = 0;
   l2274 = 0;
   l2276 = 0;
   l2278 = 0;
   l2280 = 0;
   l2282 = 0;
   l2284 = 0;
   l2286 = 0;
   l2288 = 0;
   l2290 = 0;
   l2292 = 0;
   l2294 = 0;
   l2296 = 0;
   l2298 = 0;
   l2300 = 0;
   l2302 = 0;
   l2304 = 0;
   l2306 = 0;
   l2308 = 0;
   l2310 = 0;
   l2312 = 0;
   l2314 = 0;
   l2316 = 0;
   l2318 = 0;
   l2320 = 0;
   l2322 = 0;
   l2324 = 0;
   l2326 = 0;
   l2328 = 0;
   l2330 = 0;
   l2332 = 0;
   l2334 = 0;
   l2336 = 0;
   l2338 = 0;
   l2340 = 0;
   l2342 = 0;
   l2344 = 0;
   l2346 = 0;
   l2348 = 0;
   l2350 = 0;
   l2352 = 0;
   l2354 = 0;
   l2356 = 0;
   l2358 = 0;
   l2360 = 0;
   l2362 = 0;
   l2364 = 0;
   l2366 = 0;
   l2368 = 0;
   l2370 = 0;
   l2372 = 0;
   l2374 = 0;
   l2376 = 0;
   l2378 = 0;
   l2380 = 0;
   l2382 = 0;
   l2384 = 0;
   l2386 = 0;
   l2388 = 0;
   l2390 = 0;
   l2392 = 0;
   l2394 = 0;
   l2396 = 0;
   l2398 = 0;
   l2400 = 0;
   l2402 = 0;
   l2404 = 0;
   l2406 = 0;
   l2408 = 0;
   l2410 = 0;
   l2412 = 0;
   l2414 = 0;
   l2416 = 0;
   l2418 = 0;
   l2420 = 0;
   l2422 = 0;
   l2424 = 0;
   l2426 = 0;
   l2428 = 0;
   l2430 = 0;
   l2432 = 0;
   l2434 = 0;
   l2436 = 0;
   l2438 = 0;
   l2440 = 0;
   l2442 = 0;
   l2444 = 0;
   l2446 = 0;
   l2448 = 0;
   l2450 = 0;
   l2452 = 0;
   l2454 = 0;
   l2456 = 0;
   l2458 = 0;
   l2460 = 0;
   l2462 = 0;
   l2464 = 0;
   l2466 = 0;
   l2468 = 0;
   l2470 = 0;
   l2472 = 0;
   l2474 = 0;
   l2476 = 0;
   l2478 = 0;
   l2480 = 0;
   l2482 = 0;
   l2484 = 0;
   l2486 = 0;
   l2488 = 0;
   l2490 = 0;
   l2492 = 0;
   l2494 = 0;
   l2496 = 0;
   l2498 = 0;
   l2500 = 0;
end

always @(posedge na2504)
   l880 <= na2504;

always @(posedge na2780)
   l882 <= na2780;

always @(posedge l886)
   l884 <= l886;

always @(posedge a5360)
   l886 <= a5360;

always @(posedge a17682)
   l888 <= a17682;

always @(posedge c1)
   l890 <= c1;

always @(posedge l894)
   l892 <= l894;

always @(posedge l896)
   l894 <= l896;

always @(posedge l898)
   l896 <= l898;

always @(posedge l900)
   l898 <= l900;

always @(posedge l902)
   l900 <= l902;

always @(posedge l904)
   l902 <= l904;

always @(posedge a5374)
   l904 <= a5374;

always @(posedge a16196)
   l906 <= a16196;

always @(posedge a18514)
   l908 <= a18514;

always @(posedge na18518)
   l910 <= na18518;

always @(posedge a18520)
   l912 <= a18520;

always @(posedge a18542)
   l914 <= a18542;

always @(posedge a18556)
   l916 <= a18556;

always @(posedge a18562)
   l918 <= a18562;

always @(posedge a19756)
   l920 <= a19756;

always @(posedge a19892)
   l922 <= a19892;

always @(posedge l926)
   l924 <= l926;

always @(posedge na8812)
   l926 <= na8812;

always @(posedge a19894)
   l928 <= a19894;

always @(posedge l932)
   l930 <= l932;

always @(posedge l934)
   l932 <= l934;

always @(posedge a19900)
   l934 <= a19900;

always @(posedge a16186)
   l936 <= a16186;

always @(posedge a21664)
   l938 <= a21664;

always @(posedge a23736)
   l940 <= a23736;

always @(posedge a23742)
   l942 <= a23742;

always @(posedge l946)
   l944 <= l946;

always @(posedge l948)
   l946 <= l948;

always @(posedge z0)
   l948 <= z0;

always @(posedge a8150)
   l950 <= a8150;

always @(posedge a24056)
   l952 <= a24056;

always @(posedge a24188)
   l954 <= a24188;

always @(posedge a24322)
   l956 <= a24322;

always @(posedge a24450)
   l958 <= a24450;

always @(posedge a24582)
   l960 <= a24582;

always @(posedge a24714)
   l962 <= a24714;

always @(posedge a24846)
   l964 <= a24846;

always @(posedge a24974)
   l966 <= a24974;

always @(posedge a25106)
   l968 <= a25106;

always @(posedge a25236)
   l970 <= a25236;

always @(posedge na25240)
   l972 <= na25240;

always @(posedge a25242)
   l974 <= a25242;

always @(posedge na25818)
   l976 <= na25818;

always @(posedge na19408)
   l978 <= na19408;

always @(posedge a5352)
   l980 <= a5352;

always @(posedge z1)
   l982 <= z1;

always @(posedge a25838)
   l984 <= a25838;

always @(posedge a25846)
   l986 <= a25846;

always @(posedge a25850)
   l988 <= a25850;

always @(posedge a25852)
   l990 <= a25852;

always @(posedge na26072)
   l992 <= na26072;

always @(posedge na20174)
   l994 <= na20174;

always @(posedge na26078)
   l996 <= na26078;

always @(posedge na26106)
   l998 <= na26106;

always @(posedge na26594)
   l1000 <= na26594;

always @(posedge na2536)
   l1002 <= na2536;

always @(posedge na2752)
   l1004 <= na2752;

always @(posedge na2516)
   l1006 <= na2516;

always @(posedge na26612)
   l1008 <= na26612;

always @(posedge a28188)
   l1010 <= a28188;

always @(posedge a28194)
   l1012 <= a28194;

always @(posedge a28236)
   l1014 <= a28236;

always @(posedge a20078)
   l1016 <= a20078;

always @(posedge a18850)
   l1018 <= a18850;

always @(posedge a28448)
   l1020 <= a28448;

always @(posedge a16250)
   l1022 <= a16250;

always @(posedge na28452)
   l1024 <= na28452;

always @(posedge na25504)
   l1026 <= na25504;

always @(posedge na25804)
   l1028 <= na25804;

always @(posedge a25534)
   l1030 <= a25534;

always @(posedge na28462)
   l1032 <= na28462;

always @(posedge a25578)
   l1034 <= a25578;

always @(posedge a28706)
   l1036 <= a28706;

always @(posedge a18924)
   l1038 <= a18924;

always @(posedge a28944)
   l1040 <= a28944;

always @(posedge a19004)
   l1042 <= a19004;

always @(posedge a29210)
   l1044 <= a29210;

always @(posedge a19086)
   l1046 <= a19086;

always @(posedge a29462)
   l1048 <= a29462;

always @(posedge a19168)
   l1050 <= a19168;

always @(posedge a29508)
   l1052 <= a29508;

always @(posedge na19250)
   l1054 <= na19250;

always @(posedge a29548)
   l1056 <= a29548;

always @(posedge na19332)
   l1058 <= na19332;

always @(posedge na29552)
   l1060 <= na29552;

always @(posedge a25628)
   l1062 <= a25628;

always @(posedge na29562)
   l1064 <= na29562;

always @(posedge na29572)
   l1066 <= na29572;

always @(posedge a25672)
   l1068 <= a25672;

always @(posedge na29582)
   l1070 <= na29582;

always @(posedge na25716)
   l1072 <= na25716;

always @(posedge na29592)
   l1074 <= na29592;

always @(posedge na25760)
   l1076 <= na25760;

always @(posedge na29602)
   l1078 <= na29602;

always @(posedge a29642)
   l1080 <= a29642;

always @(posedge na16278)
   l1082 <= na16278;

always @(posedge na29646)
   l1084 <= na29646;

always @(posedge na29650)
   l1086 <= na29650;

always @(posedge na29654)
   l1088 <= na29654;

always @(posedge na29658)
   l1090 <= na29658;

always @(posedge na29662)
   l1092 <= na29662;

always @(posedge a16608)
   l1094 <= a16608;

always @(posedge a29722)
   l1096 <= a29722;

always @(posedge a20054)
   l1098 <= a20054;

always @(posedge l1102)
   l1100 <= l1102;

always @(posedge z2)
   l1102 <= z2;

always @(posedge a29728)
   l1104 <= a29728;

always @(posedge a16712)
   l1106 <= a16712;

always @(posedge a29788)
   l1108 <= a29788;

always @(posedge a20028)
   l1110 <= a20028;

always @(posedge a29794)
   l1112 <= a29794;

always @(posedge a16816)
   l1114 <= a16816;

always @(posedge a29854)
   l1116 <= a29854;

always @(posedge a20002)
   l1118 <= a20002;

always @(posedge a29860)
   l1120 <= a29860;

always @(posedge a16920)
   l1122 <= a16920;

always @(posedge a29920)
   l1124 <= a29920;

always @(posedge a19976)
   l1126 <= a19976;

always @(posedge a29926)
   l1128 <= a29926;

always @(posedge na17016)
   l1130 <= na17016;

always @(posedge a29986)
   l1132 <= a29986;

always @(posedge na19950)
   l1134 <= na19950;

always @(posedge na29992)
   l1136 <= na29992;

always @(posedge na17112)
   l1138 <= na17112;

always @(posedge na30052)
   l1140 <= na30052;

always @(posedge na19922)
   l1142 <= na19922;

always @(posedge na30058)
   l1144 <= na30058;

always @(posedge na8954)
   l1146 <= na8954;

always @(posedge na30072)
   l1148 <= na30072;

always @(posedge a31018)
   l1150 <= a31018;

always @(posedge a31020)
   l1152 <= a31020;

always @(posedge a31040)
   l1154 <= a31040;

always @(posedge na31048)
   l1156 <= na31048;

always @(posedge a8946)
   l1158 <= a8946;

always @(posedge na8986)
   l1160 <= na8986;

always @(posedge na31060)
   l1162 <= na31060;

always @(posedge na31072)
   l1164 <= na31072;

always @(posedge na31086)
   l1166 <= na31086;

always @(posedge na8924)
   l1168 <= na8924;

always @(posedge na8870)
   l1170 <= na8870;

always @(posedge l1174)
   l1172 <= l1174;

always @(posedge a31088)
   l1174 <= a31088;

always @(posedge l1178)
   l1176 <= l1178;

always @(posedge l1180)
   l1178 <= l1180;

always @(posedge l1182)
   l1180 <= l1182;

always @(posedge l1184)
   l1182 <= l1184;

always @(posedge na31092)
   l1184 <= na31092;

always @(posedge z3)
   l1186 <= z3;

always @(posedge na31152)
   l1188 <= na31152;

always @(posedge na18526)
   l1190 <= na18526;

always @(posedge a31160)
   l1192 <= a31160;

always @(posedge na17784)
   l1194 <= na17784;

always @(posedge l1198)
   l1196 <= l1198;

always @(posedge z4)
   l1198 <= z4;

always @(posedge l1202)
   l1200 <= l1202;

always @(posedge l1204)
   l1202 <= l1204;

always @(posedge l1206)
   l1204 <= l1206;

always @(posedge l1208)
   l1206 <= l1208;

always @(posedge na31102)
   l1208 <= na31102;

always @(posedge na31176)
   l1210 <= na31176;

always @(posedge a31182)
   l1212 <= a31182;

always @(posedge a8970)
   l1214 <= a8970;

always @(posedge l1218)
   l1216 <= l1218;

always @(posedge l1220)
   l1218 <= l1220;

always @(posedge l1222)
   l1220 <= l1222;

always @(posedge l1224)
   l1222 <= l1224;

always @(posedge na31110)
   l1224 <= na31110;

always @(posedge na31202)
   l1226 <= na31202;

always @(posedge a31208)
   l1228 <= a31208;

always @(posedge a9006)
   l1230 <= a9006;

always @(posedge l1234)
   l1232 <= l1234;

always @(posedge l1236)
   l1234 <= l1236;

always @(posedge l1238)
   l1236 <= l1238;

always @(posedge l1240)
   l1238 <= l1240;

always @(posedge na31118)
   l1240 <= na31118;

always @(posedge na31222)
   l1242 <= na31222;

always @(posedge na31228)
   l1244 <= na31228;

always @(posedge na8906)
   l1246 <= na8906;

always @(posedge a32370)
   l1248 <= a32370;

always @(posedge a32380)
   l1250 <= a32380;

always @(posedge na12366)
   l1252 <= na12366;

always @(posedge na32396)
   l1254 <= na32396;

always @(posedge a32386)
   l1256 <= a32386;

always @(posedge na32402)
   l1258 <= na32402;

always @(posedge na12312)
   l1260 <= na12312;

always @(posedge na32408)
   l1262 <= na32408;

always @(posedge na32414)
   l1264 <= na32414;

always @(posedge na12250)
   l1266 <= na12250;

always @(posedge na32420)
   l1268 <= na32420;

always @(posedge na32426)
   l1270 <= na32426;

always @(posedge na12190)
   l1272 <= na12190;

always @(posedge na32432)
   l1274 <= na32432;

always @(posedge na32438)
   l1276 <= na32438;

always @(posedge na16376)
   l1278 <= na16376;

always @(posedge na17092)
   l1280 <= na17092;

always @(posedge na18282)
   l1282 <= na18282;

always @(posedge a16996)
   l1284 <= a16996;

always @(posedge na18208)
   l1286 <= na18208;

always @(posedge a16892)
   l1288 <= a16892;

always @(posedge na18134)
   l1290 <= na18134;

always @(posedge a16788)
   l1292 <= a16788;

always @(posedge na18060)
   l1294 <= na18060;

always @(posedge a16684)
   l1296 <= a16684;

always @(posedge na17986)
   l1298 <= na17986;

always @(posedge a16580)
   l1300 <= a16580;

always @(posedge na17912)
   l1302 <= na17912;

always @(posedge a16514)
   l1304 <= a16514;

always @(posedge na17844)
   l1306 <= na17844;

always @(posedge na32454)
   l1308 <= na32454;

always @(posedge a32470)
   l1310 <= a32470;

always @(posedge a32486)
   l1312 <= a32486;

always @(posedge na22814)
   l1314 <= na22814;

always @(posedge na22822)
   l1316 <= na22822;

always @(posedge na22834)
   l1318 <= na22834;

always @(posedge na22842)
   l1320 <= na22842;

always @(posedge na22854)
   l1322 <= na22854;

always @(posedge na22862)
   l1324 <= na22862;

always @(posedge na22878)
   l1326 <= na22878;

always @(posedge na22886)
   l1328 <= na22886;

always @(posedge na22898)
   l1330 <= na22898;

always @(posedge na22906)
   l1332 <= na22906;

always @(posedge na21710)
   l1334 <= na21710;

always @(posedge na21720)
   l1336 <= na21720;

always @(posedge na21740)
   l1338 <= na21740;

always @(posedge na21752)
   l1340 <= na21752;

always @(posedge na21766)
   l1342 <= na21766;

always @(posedge na21776)
   l1344 <= na21776;

always @(posedge a21800)
   l1346 <= a21800;

always @(posedge a21810)
   l1348 <= a21810;

always @(posedge a21828)
   l1350 <= a21828;

always @(posedge na21840)
   l1352 <= na21840;

always @(posedge na21886)
   l1354 <= na21886;

always @(posedge na21894)
   l1356 <= na21894;

always @(posedge na21906)
   l1358 <= na21906;

always @(posedge na21914)
   l1360 <= na21914;

always @(posedge na21926)
   l1362 <= na21926;

always @(posedge na21934)
   l1364 <= na21934;

always @(posedge a21950)
   l1366 <= a21950;

always @(posedge a21958)
   l1368 <= a21958;

always @(posedge a21970)
   l1370 <= a21970;

always @(posedge na21978)
   l1372 <= na21978;

always @(posedge na22020)
   l1374 <= na22020;

always @(posedge na22028)
   l1376 <= na22028;

always @(posedge na22040)
   l1378 <= na22040;

always @(posedge na22048)
   l1380 <= na22048;

always @(posedge na22060)
   l1382 <= na22060;

always @(posedge na22068)
   l1384 <= na22068;

always @(posedge a22084)
   l1386 <= a22084;

always @(posedge a22092)
   l1388 <= a22092;

always @(posedge a22104)
   l1390 <= a22104;

always @(posedge na22112)
   l1392 <= na22112;

always @(posedge na22154)
   l1394 <= na22154;

always @(posedge na22162)
   l1396 <= na22162;

always @(posedge na22174)
   l1398 <= na22174;

always @(posedge na22182)
   l1400 <= na22182;

always @(posedge na22194)
   l1402 <= na22194;

always @(posedge na22202)
   l1404 <= na22202;

always @(posedge a22218)
   l1406 <= a22218;

always @(posedge a22226)
   l1408 <= a22226;

always @(posedge a22238)
   l1410 <= a22238;

always @(posedge na22246)
   l1412 <= na22246;

always @(posedge na22288)
   l1414 <= na22288;

always @(posedge na22296)
   l1416 <= na22296;

always @(posedge na22308)
   l1418 <= na22308;

always @(posedge na22316)
   l1420 <= na22316;

always @(posedge na22328)
   l1422 <= na22328;

always @(posedge na22336)
   l1424 <= na22336;

always @(posedge a22352)
   l1426 <= a22352;

always @(posedge a22360)
   l1428 <= a22360;

always @(posedge a22372)
   l1430 <= a22372;

always @(posedge na22380)
   l1432 <= na22380;

always @(posedge na22422)
   l1434 <= na22422;

always @(posedge na22430)
   l1436 <= na22430;

always @(posedge na22442)
   l1438 <= na22442;

always @(posedge na22450)
   l1440 <= na22450;

always @(posedge na22462)
   l1442 <= na22462;

always @(posedge na22470)
   l1444 <= na22470;

always @(posedge a22486)
   l1446 <= a22486;

always @(posedge a22494)
   l1448 <= a22494;

always @(posedge a22506)
   l1450 <= a22506;

always @(posedge na22514)
   l1452 <= na22514;

always @(posedge na22556)
   l1454 <= na22556;

always @(posedge na22564)
   l1456 <= na22564;

always @(posedge na22576)
   l1458 <= na22576;

always @(posedge na22584)
   l1460 <= na22584;

always @(posedge na22596)
   l1462 <= na22596;

always @(posedge na22604)
   l1464 <= na22604;

always @(posedge a22620)
   l1466 <= a22620;

always @(posedge a22628)
   l1468 <= a22628;

always @(posedge na22640)
   l1470 <= na22640;

always @(posedge na22648)
   l1472 <= na22648;

always @(posedge na26200)
   l1474 <= na26200;

always @(posedge na26238)
   l1476 <= na26238;

always @(posedge na26282)
   l1478 <= na26282;

always @(posedge na26326)
   l1480 <= na26326;

always @(posedge na26370)
   l1482 <= na26370;

always @(posedge na26414)
   l1484 <= na26414;

always @(posedge a32504)
   l1486 <= a32504;

always @(posedge a32508)
   l1488 <= a32508;

always @(posedge a32538)
   l1490 <= a32538;

always @(posedge a16440)
   l1492 <= a16440;

always @(posedge na33374)
   l1494 <= na33374;

always @(posedge na33380)
   l1496 <= na33380;

always @(posedge na33402)
   l1498 <= na33402;

always @(posedge na33408)
   l1500 <= na33408;

always @(posedge a33430)
   l1502 <= a33430;

always @(posedge na33436)
   l1504 <= na33436;

always @(posedge a33458)
   l1506 <= a33458;

always @(posedge na33464)
   l1508 <= na33464;

always @(posedge a32966)
   l1510 <= a32966;

always @(posedge na33468)
   l1512 <= na33468;

always @(posedge a32978)
   l1514 <= a32978;

always @(posedge l1518)
   l1516 <= l1518;

always @(posedge l1520)
   l1518 <= l1520;

always @(posedge l1522)
   l1520 <= l1522;

always @(posedge na33506)
   l1522 <= na33506;

always @(posedge na33526)
   l1524 <= na33526;

always @(posedge a31042)
   l1526 <= a31042;

always @(posedge na24030)
   l1528 <= na24030;

always @(posedge na33570)
   l1530 <= na33570;

always @(posedge na33624)
   l1532 <= na33624;

always @(posedge na33636)
   l1534 <= na33636;

always @(posedge na33642)
   l1536 <= na33642;

always @(posedge na33652)
   l1538 <= na33652;

always @(posedge a34176)
   l1540 <= a34176;

always @(posedge a32998)
   l1542 <= a32998;

always @(posedge z5)
   l1544 <= z5;

always @(posedge na23774)
   l1546 <= na23774;

always @(posedge na24826)
   l1548 <= na24826;

always @(posedge na34252)
   l1550 <= na34252;

always @(posedge na34268)
   l1552 <= na34268;

always @(posedge na34290)
   l1554 <= na34290;

always @(posedge na34308)
   l1556 <= na34308;

always @(posedge na34326)
   l1558 <= na34326;

always @(posedge na25216)
   l1560 <= na25216;

always @(posedge a34338)
   l1562 <= a34338;

always @(posedge na24954)
   l1564 <= na24954;

always @(posedge na34350)
   l1566 <= na34350;

always @(posedge a34362)
   l1568 <= a34362;

always @(posedge na24694)
   l1570 <= na24694;

always @(posedge na24562)
   l1572 <= na24562;

always @(posedge na24430)
   l1574 <= na24430;

always @(posedge na24302)
   l1576 <= na24302;

always @(posedge na24168)
   l1578 <= na24168;

always @(posedge na24036)
   l1580 <= na24036;

always @(posedge na25086)
   l1582 <= na25086;

always @(posedge a33014)
   l1584 <= a33014;

always @(posedge a33032)
   l1586 <= a33032;

always @(posedge a33046)
   l1588 <= a33046;

always @(posedge a33066)
   l1590 <= a33066;

always @(posedge a33078)
   l1592 <= a33078;

always @(posedge a33094)
   l1594 <= a33094;

always @(posedge a33106)
   l1596 <= a33106;

always @(posedge na34374)
   l1598 <= na34374;

always @(posedge na34380)
   l1600 <= na34380;

always @(posedge na34386)
   l1602 <= na34386;

always @(posedge na34392)
   l1604 <= na34392;

always @(posedge na34398)
   l1606 <= na34398;

always @(posedge na34404)
   l1608 <= na34404;

always @(posedge na34410)
   l1610 <= na34410;

always @(posedge na34416)
   l1612 <= na34416;

always @(posedge na34422)
   l1614 <= na34422;

always @(posedge na34428)
   l1616 <= na34428;

always @(posedge na34440)
   l1618 <= na34440;

always @(posedge na34446)
   l1620 <= na34446;

always @(posedge na34452)
   l1622 <= na34452;

always @(posedge na34458)
   l1624 <= na34458;

always @(posedge na34464)
   l1626 <= na34464;

always @(posedge na34470)
   l1628 <= na34470;

always @(posedge na34476)
   l1630 <= na34476;

always @(posedge na34482)
   l1632 <= na34482;

always @(posedge a34488)
   l1634 <= a34488;

always @(posedge a34494)
   l1636 <= a34494;

always @(posedge na34506)
   l1638 <= na34506;

always @(posedge na34512)
   l1640 <= na34512;

always @(posedge na34518)
   l1642 <= na34518;

always @(posedge na34524)
   l1644 <= na34524;

always @(posedge na34530)
   l1646 <= na34530;

always @(posedge na34536)
   l1648 <= na34536;

always @(posedge na34542)
   l1650 <= na34542;

always @(posedge na34548)
   l1652 <= na34548;

always @(posedge a34554)
   l1654 <= a34554;

always @(posedge a34560)
   l1656 <= a34560;

always @(posedge na34572)
   l1658 <= na34572;

always @(posedge na34578)
   l1660 <= na34578;

always @(posedge na34584)
   l1662 <= na34584;

always @(posedge na34590)
   l1664 <= na34590;

always @(posedge na34596)
   l1666 <= na34596;

always @(posedge na34602)
   l1668 <= na34602;

always @(posedge na34608)
   l1670 <= na34608;

always @(posedge na34614)
   l1672 <= na34614;

always @(posedge a34620)
   l1674 <= a34620;

always @(posedge a34626)
   l1676 <= a34626;

always @(posedge na34638)
   l1678 <= na34638;

always @(posedge na34644)
   l1680 <= na34644;

always @(posedge na34650)
   l1682 <= na34650;

always @(posedge na34656)
   l1684 <= na34656;

always @(posedge na34662)
   l1686 <= na34662;

always @(posedge na34668)
   l1688 <= na34668;

always @(posedge na34674)
   l1690 <= na34674;

always @(posedge na34680)
   l1692 <= na34680;

always @(posedge a34686)
   l1694 <= a34686;

always @(posedge a34692)
   l1696 <= a34692;

always @(posedge na34704)
   l1698 <= na34704;

always @(posedge na34710)
   l1700 <= na34710;

always @(posedge na34716)
   l1702 <= na34716;

always @(posedge na34722)
   l1704 <= na34722;

always @(posedge na34728)
   l1706 <= na34728;

always @(posedge na34734)
   l1708 <= na34734;

always @(posedge na34740)
   l1710 <= na34740;

always @(posedge na34746)
   l1712 <= na34746;

always @(posedge a34752)
   l1714 <= a34752;

always @(posedge a34758)
   l1716 <= a34758;

always @(posedge na34770)
   l1718 <= na34770;

always @(posedge na34776)
   l1720 <= na34776;

always @(posedge na34782)
   l1722 <= na34782;

always @(posedge na34788)
   l1724 <= na34788;

always @(posedge na34794)
   l1726 <= na34794;

always @(posedge na34800)
   l1728 <= na34800;

always @(posedge na34806)
   l1730 <= na34806;

always @(posedge na34812)
   l1732 <= na34812;

always @(posedge a34818)
   l1734 <= a34818;

always @(posedge na34824)
   l1736 <= na34824;

always @(posedge na34836)
   l1738 <= na34836;

always @(posedge na34842)
   l1740 <= na34842;

always @(posedge na34848)
   l1742 <= na34848;

always @(posedge na34854)
   l1744 <= na34854;

always @(posedge na34860)
   l1746 <= na34860;

always @(posedge na34866)
   l1748 <= na34866;

always @(posedge na34872)
   l1750 <= na34872;

always @(posedge na34878)
   l1752 <= na34878;

always @(posedge na34884)
   l1754 <= na34884;

always @(posedge na34890)
   l1756 <= na34890;

always @(posedge a34894)
   l1758 <= a34894;

always @(posedge z6)
   l1760 <= z6;

always @(posedge z7)
   l1762 <= z7;

always @(posedge z8)
   l1764 <= z8;

always @(posedge na17454)
   l1766 <= na17454;

always @(posedge a34896)
   l1768 <= a34896;

always @(posedge a34898)
   l1770 <= a34898;

always @(posedge a34900)
   l1772 <= a34900;

always @(posedge a34902)
   l1774 <= a34902;

always @(posedge na17592)
   l1776 <= na17592;

always @(posedge a34904)
   l1778 <= a34904;

always @(posedge a34910)
   l1780 <= a34910;

always @(posedge a21670)
   l1782 <= a21670;

always @(posedge na34920)
   l1784 <= na34920;

always @(posedge na34928)
   l1786 <= na34928;

always @(posedge na34936)
   l1788 <= na34936;

always @(posedge na34946)
   l1790 <= na34946;

always @(posedge na34954)
   l1792 <= na34954;

always @(posedge na34962)
   l1794 <= na34962;

always @(posedge na34970)
   l1796 <= na34970;

always @(posedge na34976)
   l1798 <= na34976;

always @(posedge a34988)
   l1800 <= a34988;

always @(posedge a21880)
   l1802 <= a21880;

always @(posedge na34994)
   l1804 <= na34994;

always @(posedge a35000)
   l1806 <= a35000;

always @(posedge na35006)
   l1808 <= na35006;

always @(posedge na35012)
   l1810 <= na35012;

always @(posedge na35018)
   l1812 <= na35018;

always @(posedge na35024)
   l1814 <= na35024;

always @(posedge na35030)
   l1816 <= na35030;

always @(posedge na35036)
   l1818 <= na35036;

always @(posedge na35042)
   l1820 <= na35042;

always @(posedge a35054)
   l1822 <= a35054;

always @(posedge a22014)
   l1824 <= a22014;

always @(posedge na35060)
   l1826 <= na35060;

always @(posedge a35066)
   l1828 <= a35066;

always @(posedge na35072)
   l1830 <= na35072;

always @(posedge na35078)
   l1832 <= na35078;

always @(posedge na35084)
   l1834 <= na35084;

always @(posedge na35090)
   l1836 <= na35090;

always @(posedge na35096)
   l1838 <= na35096;

always @(posedge na35102)
   l1840 <= na35102;

always @(posedge na35108)
   l1842 <= na35108;

always @(posedge a35120)
   l1844 <= a35120;

always @(posedge a22148)
   l1846 <= a22148;

always @(posedge na35126)
   l1848 <= na35126;

always @(posedge a35132)
   l1850 <= a35132;

always @(posedge na35138)
   l1852 <= na35138;

always @(posedge na35144)
   l1854 <= na35144;

always @(posedge na35150)
   l1856 <= na35150;

always @(posedge na35156)
   l1858 <= na35156;

always @(posedge na35162)
   l1860 <= na35162;

always @(posedge na35168)
   l1862 <= na35168;

always @(posedge na35174)
   l1864 <= na35174;

always @(posedge a35186)
   l1866 <= a35186;

always @(posedge a22282)
   l1868 <= a22282;

always @(posedge na35192)
   l1870 <= na35192;

always @(posedge a35198)
   l1872 <= a35198;

always @(posedge na35204)
   l1874 <= na35204;

always @(posedge na35210)
   l1876 <= na35210;

always @(posedge na35216)
   l1878 <= na35216;

always @(posedge na35222)
   l1880 <= na35222;

always @(posedge na35228)
   l1882 <= na35228;

always @(posedge na35234)
   l1884 <= na35234;

always @(posedge na35240)
   l1886 <= na35240;

always @(posedge a35252)
   l1888 <= a35252;

always @(posedge a22416)
   l1890 <= a22416;

always @(posedge na35258)
   l1892 <= na35258;

always @(posedge a35264)
   l1894 <= a35264;

always @(posedge na35270)
   l1896 <= na35270;

always @(posedge na35276)
   l1898 <= na35276;

always @(posedge na35282)
   l1900 <= na35282;

always @(posedge na35288)
   l1902 <= na35288;

always @(posedge na35294)
   l1904 <= na35294;

always @(posedge na35300)
   l1906 <= na35300;

always @(posedge na35306)
   l1908 <= na35306;

always @(posedge na35318)
   l1910 <= na35318;

always @(posedge a22550)
   l1912 <= a22550;

always @(posedge na35324)
   l1914 <= na35324;

always @(posedge a35330)
   l1916 <= a35330;

always @(posedge na35336)
   l1918 <= na35336;

always @(posedge na35342)
   l1920 <= na35342;

always @(posedge na35348)
   l1922 <= na35348;

always @(posedge na35354)
   l1924 <= na35354;

always @(posedge na35360)
   l1926 <= na35360;

always @(posedge na35366)
   l1928 <= na35366;

always @(posedge na35372)
   l1930 <= na35372;

always @(posedge na35386)
   l1932 <= na35386;

always @(posedge a22808)
   l1934 <= a22808;

always @(posedge na35392)
   l1936 <= na35392;

always @(posedge na35398)
   l1938 <= na35398;

always @(posedge na35404)
   l1940 <= na35404;

always @(posedge na35410)
   l1942 <= na35410;

always @(posedge na35416)
   l1944 <= na35416;

always @(posedge na35422)
   l1946 <= na35422;

always @(posedge na35428)
   l1948 <= na35428;

always @(posedge na35434)
   l1950 <= na35434;

always @(posedge na35440)
   l1952 <= na35440;

always @(posedge a35472)
   l1954 <= a35472;

always @(posedge l1958)
   l1956 <= l1958;

always @(posedge na8846)
   l1958 <= na8846;

always @(posedge l1962)
   l1960 <= l1962;

always @(posedge na8836)
   l1962 <= na8836;

always @(posedge l1966)
   l1964 <= l1966;

always @(posedge na8860)
   l1966 <= na8860;

always @(posedge l1970)
   l1968 <= l1970;

always @(posedge na8826)
   l1970 <= na8826;

always @(posedge a35514)
   l1972 <= a35514;

always @(posedge a35554)
   l1974 <= a35554;

always @(posedge a35588)
   l1976 <= a35588;

always @(posedge a35636)
   l1978 <= a35636;

always @(posedge a35664)
   l1980 <= a35664;

always @(posedge a35700)
   l1982 <= a35700;

always @(posedge a35720)
   l1984 <= a35720;

always @(posedge a35748)
   l1986 <= a35748;

always @(posedge na35754)
   l1988 <= na35754;

always @(posedge na35760)
   l1990 <= na35760;

always @(posedge na35766)
   l1992 <= na35766;

always @(posedge na35772)
   l1994 <= na35772;

always @(posedge na35778)
   l1996 <= na35778;

always @(posedge na35784)
   l1998 <= na35784;

always @(posedge na35790)
   l2000 <= na35790;

always @(posedge na35796)
   l2002 <= na35796;

always @(posedge na35802)
   l2004 <= na35802;

always @(posedge a32592)
   l2006 <= a32592;

always @(posedge a32634)
   l2008 <= a32634;

always @(posedge a32680)
   l2010 <= a32680;

always @(posedge a32722)
   l2012 <= a32722;

always @(posedge a32772)
   l2014 <= a32772;

always @(posedge a32814)
   l2016 <= a32814;

always @(posedge a32860)
   l2018 <= a32860;

always @(posedge a32908)
   l2020 <= a32908;

always @(posedge a33156)
   l2022 <= a33156;

always @(posedge a33198)
   l2024 <= a33198;

always @(posedge na35828)
   l2026 <= na35828;

always @(posedge l2030)
   l2028 <= l2030;

always @(posedge z9)
   l2030 <= z9;

always @(posedge l2034)
   l2032 <= l2034;

always @(posedge z10)
   l2034 <= z10;

always @(posedge l2038)
   l2036 <= l2038;

always @(posedge z11)
   l2038 <= z11;

always @(posedge l2042)
   l2040 <= l2042;

always @(posedge z12)
   l2042 <= z12;

always @(posedge na35836)
   l2044 <= na35836;

always @(posedge na35856)
   l2046 <= na35856;

always @(posedge na35862)
   l2048 <= na35862;

always @(posedge na35880)
   l2050 <= na35880;

always @(posedge na35886)
   l2052 <= na35886;

always @(posedge na35896)
   l2054 <= na35896;

always @(posedge na35902)
   l2056 <= na35902;

always @(posedge na35912)
   l2058 <= na35912;

always @(posedge na35922)
   l2060 <= na35922;

always @(posedge na18744)
   l2062 <= na18744;

always @(posedge a35930)
   l2064 <= a35930;

always @(posedge z13)
   l2066 <= z13;

always @(posedge a35946)
   l2068 <= a35946;

always @(posedge a35960)
   l2070 <= a35960;

always @(posedge a35968)
   l2072 <= a35968;

always @(posedge na36056)
   l2074 <= na36056;

always @(posedge na37126)
   l2076 <= na37126;

always @(posedge na37160)
   l2078 <= na37160;

always @(posedge na37184)
   l2080 <= na37184;

always @(posedge na37206)
   l2082 <= na37206;

always @(posedge na37222)
   l2084 <= na37222;

always @(posedge na37246)
   l2086 <= na37246;

always @(posedge na37266)
   l2088 <= na37266;

always @(posedge na37386)
   l2090 <= na37386;

always @(posedge na37400)
   l2092 <= na37400;

always @(posedge na37448)
   l2094 <= na37448;

always @(posedge na37476)
   l2096 <= na37476;

always @(posedge na37482)
   l2098 <= na37482;

always @(posedge i252)
   l2100 <= i252;

always @(posedge a41638)
   l2102 <= a41638;

always @(posedge a41644)
   l2104 <= a41644;

always @(posedge i650)
   l2106 <= i650;

always @(posedge na41660)
   l2108 <= na41660;

always @(posedge a41670)
   l2110 <= a41670;

always @(posedge a41672)
   l2112 <= a41672;

always @(posedge na41678)
   l2114 <= na41678;

always @(posedge a41736)
   l2116 <= a41736;

always @(posedge na41742)
   l2118 <= na41742;

always @(posedge na41800)
   l2120 <= na41800;

always @(posedge na41806)
   l2122 <= na41806;

always @(posedge na41846)
   l2124 <= na41846;

always @(posedge a44408)
   l2126 <= a44408;

always @(posedge a44428)
   l2128 <= a44428;

always @(posedge a41654)
   l2130 <= a41654;

always @(posedge a44442)
   l2132 <= a44442;

always @(posedge a44450)
   l2134 <= a44450;

always @(posedge a44462)
   l2136 <= a44462;

always @(posedge a44472)
   l2138 <= a44472;

always @(posedge a44482)
   l2140 <= a44482;

always @(posedge a44490)
   l2142 <= a44490;

always @(posedge a44498)
   l2144 <= a44498;

always @(posedge a44506)
   l2146 <= a44506;

always @(posedge a44514)
   l2148 <= a44514;

always @(posedge a44520)
   l2150 <= a44520;

always @(posedge a44526)
   l2152 <= a44526;

always @(posedge a44532)
   l2154 <= a44532;

always @(posedge a44538)
   l2156 <= a44538;

always @(posedge a44544)
   l2158 <= a44544;

always @(posedge a44550)
   l2160 <= a44550;

always @(posedge a44556)
   l2162 <= a44556;

always @(posedge a44562)
   l2164 <= a44562;

always @(posedge a44568)
   l2166 <= a44568;

always @(posedge a44574)
   l2168 <= a44574;

always @(posedge a44580)
   l2170 <= a44580;

always @(posedge a44586)
   l2172 <= a44586;

always @(posedge a44592)
   l2174 <= a44592;

always @(posedge a44598)
   l2176 <= a44598;

always @(posedge a44604)
   l2178 <= a44604;

always @(posedge a44610)
   l2180 <= a44610;

always @(posedge a44616)
   l2182 <= a44616;

always @(posedge a44622)
   l2184 <= a44622;

always @(posedge a44628)
   l2186 <= a44628;

always @(posedge a44634)
   l2188 <= a44634;

always @(posedge a44640)
   l2190 <= a44640;

always @(posedge a44646)
   l2192 <= a44646;

always @(posedge a44652)
   l2194 <= a44652;

always @(posedge a44658)
   l2196 <= a44658;

always @(posedge a44664)
   l2198 <= a44664;

always @(posedge a44670)
   l2200 <= a44670;

always @(posedge a44676)
   l2202 <= a44676;

always @(posedge a44682)
   l2204 <= a44682;

always @(posedge a44688)
   l2206 <= a44688;

always @(posedge a44694)
   l2208 <= a44694;

always @(posedge a44700)
   l2210 <= a44700;

always @(posedge a44706)
   l2212 <= a44706;

always @(posedge a44712)
   l2214 <= a44712;

always @(posedge a44718)
   l2216 <= a44718;

always @(posedge a44724)
   l2218 <= a44724;

always @(posedge a44730)
   l2220 <= a44730;

always @(posedge a44736)
   l2222 <= a44736;

always @(posedge a44742)
   l2224 <= a44742;

always @(posedge a44748)
   l2226 <= a44748;

always @(posedge a44754)
   l2228 <= a44754;

always @(posedge a44760)
   l2230 <= a44760;

always @(posedge a44766)
   l2232 <= a44766;

always @(posedge a44772)
   l2234 <= a44772;

always @(posedge a44778)
   l2236 <= a44778;

always @(posedge a44784)
   l2238 <= a44784;

always @(posedge a44790)
   l2240 <= a44790;

always @(posedge a44796)
   l2242 <= a44796;

always @(posedge a44802)
   l2244 <= a44802;

always @(posedge a44808)
   l2246 <= a44808;

always @(posedge a44814)
   l2248 <= a44814;

always @(posedge a44834)
   l2250 <= a44834;

always @(posedge a45596)
   l2252 <= a45596;

always @(posedge na8818)
   l2254 <= na8818;

always @(posedge l2258)
   l2256 <= l2258;

always @(posedge l2260)
   l2258 <= l2260;

always @(posedge l2262)
   l2260 <= l2262;

always @(posedge z14)
   l2262 <= z14;

always @(posedge a8814)
   l2264 <= a8814;

always @(posedge z15)
   l2266 <= z15;

always @(posedge z16)
   l2268 <= z16;

always @(posedge z17)
   l2270 <= z17;

always @(posedge l2274)
   l2272 <= l2274;

always @(posedge l2276)
   l2274 <= l2276;

always @(posedge l2278)
   l2276 <= l2278;

always @(posedge l2280)
   l2278 <= l2280;

always @(posedge l2282)
   l2280 <= l2282;

always @(posedge na40992)
   l2282 <= na40992;

always @(posedge l2286)
   l2284 <= l2286;

always @(posedge l2288)
   l2286 <= l2288;

always @(posedge l2290)
   l2288 <= l2290;

always @(posedge na45602)
   l2290 <= na45602;

always @(posedge a45608)
   l2292 <= a45608;

always @(posedge a40642)
   l2294 <= a40642;

always @(posedge l2298)
   l2296 <= l2298;

always @(posedge l2300)
   l2298 <= l2300;

always @(posedge l2302)
   l2300 <= l2302;

always @(posedge l2304)
   l2302 <= l2304;

always @(posedge l2306)
   l2304 <= l2306;

always @(posedge z18)
   l2306 <= z18;

always @(posedge a45622)
   l2308 <= a45622;

always @(posedge a46176)
   l2310 <= a46176;

always @(posedge a48022)
   l2312 <= a48022;

always @(posedge a48034)
   l2314 <= a48034;

always @(posedge a48048)
   l2316 <= a48048;

always @(posedge na48062)
   l2318 <= na48062;

always @(posedge a48584)
   l2320 <= a48584;

always @(posedge a48590)
   l2322 <= a48590;

always @(posedge a48596)
   l2324 <= a48596;

always @(posedge a48602)
   l2326 <= a48602;

always @(posedge a48608)
   l2328 <= a48608;

always @(posedge a48614)
   l2330 <= a48614;

always @(posedge a48620)
   l2332 <= a48620;

always @(posedge a48626)
   l2334 <= a48626;

always @(posedge a48632)
   l2336 <= a48632;

always @(posedge a48638)
   l2338 <= a48638;

always @(posedge a48644)
   l2340 <= a48644;

always @(posedge a48650)
   l2342 <= a48650;

always @(posedge a48656)
   l2344 <= a48656;

always @(posedge a48662)
   l2346 <= a48662;

always @(posedge a48668)
   l2348 <= a48668;

always @(posedge a48674)
   l2350 <= a48674;

always @(posedge a48680)
   l2352 <= a48680;

always @(posedge a48686)
   l2354 <= a48686;

always @(posedge a48692)
   l2356 <= a48692;

always @(posedge a48698)
   l2358 <= a48698;

always @(posedge a48704)
   l2360 <= a48704;

always @(posedge a48728)
   l2362 <= a48728;

always @(posedge a48792)
   l2364 <= a48792;

always @(posedge a48808)
   l2366 <= a48808;

always @(posedge a49932)
   l2368 <= a49932;

always @(posedge na49946)
   l2370 <= na49946;

always @(posedge na49958)
   l2372 <= na49958;

always @(posedge a49740)
   l2374 <= a49740;

always @(posedge a49996)
   l2376 <= a49996;

always @(posedge a49758)
   l2378 <= a49758;

always @(posedge a50024)
   l2380 <= a50024;

always @(posedge a49784)
   l2382 <= a49784;

always @(posedge a50066)
   l2384 <= a50066;

always @(posedge a50084)
   l2386 <= a50084;

always @(posedge a49802)
   l2388 <= a49802;

always @(posedge a50114)
   l2390 <= a50114;

always @(posedge a49824)
   l2392 <= a49824;

always @(posedge a49842)
   l2394 <= a49842;

always @(posedge a50136)
   l2396 <= a50136;

always @(posedge a49862)
   l2398 <= a49862;

always @(posedge a50164)
   l2400 <= a50164;

always @(posedge a49880)
   l2402 <= a49880;

always @(posedge a50176)
   l2404 <= a50176;

always @(posedge l2408)
   l2406 <= l2408;

always @(posedge z19)
   l2408 <= z19;

always @(posedge l2412)
   l2410 <= l2412;

always @(posedge z20)
   l2412 <= z20;

always @(posedge l2416)
   l2414 <= l2416;

always @(posedge z21)
   l2416 <= z21;

always @(posedge l2420)
   l2418 <= l2420;

always @(posedge z22)
   l2420 <= z22;

always @(posedge na50182)
   l2422 <= na50182;

always @(posedge na50188)
   l2424 <= na50188;

always @(posedge na50194)
   l2426 <= na50194;

always @(posedge na50200)
   l2428 <= na50200;

always @(posedge na50248)
   l2430 <= na50248;

always @(posedge na50254)
   l2432 <= na50254;

always @(posedge na50260)
   l2434 <= na50260;

always @(posedge na50266)
   l2436 <= na50266;

always @(posedge na50272)
   l2438 <= na50272;

always @(posedge na50278)
   l2440 <= na50278;

always @(posedge na50284)
   l2442 <= na50284;

always @(posedge a50346)
   l2444 <= a50346;

always @(posedge a50420)
   l2446 <= a50420;

always @(posedge na50426)
   l2448 <= na50426;

always @(posedge a50620)
   l2450 <= a50620;

always @(posedge a50646)
   l2452 <= a50646;

always @(posedge a50672)
   l2454 <= a50672;

always @(posedge a50698)
   l2456 <= a50698;

always @(posedge a50724)
   l2458 <= a50724;

always @(posedge a50750)
   l2460 <= a50750;

always @(posedge a50776)
   l2462 <= a50776;

always @(posedge a50802)
   l2464 <= a50802;

always @(posedge a50828)
   l2466 <= a50828;

always @(posedge a50854)
   l2468 <= a50854;

always @(posedge na50954)
   l2470 <= na50954;

always @(posedge na50958)
   l2472 <= na50958;

always @(posedge na50962)
   l2474 <= na50962;

always @(posedge na50970)
   l2476 <= na50970;

always @(posedge a50972)
   l2478 <= a50972;

always @(posedge na18534)
   l2480 <= na18534;

always @(posedge a50986)
   l2482 <= a50986;

always @(posedge a50990)
   l2484 <= a50990;

always @(posedge na50996)
   l2486 <= na50996;

always @(posedge a51000)
   l2488 <= a51000;

always @(posedge a5624)
   l2490 <= a5624;

always @(posedge z23)
   l2492 <= z23;

always @(posedge z24)
   l2494 <= z24;

always @(posedge z25)
   l2496 <= z25;

always @(posedge z26)
   l2498 <= z26;

always @(posedge z27)
   l2500 <= z27;


assign na2504 = ~a2504;
assign na2780 = ~a2780;
assign a5360 = ~a5358 & a5352;
assign a17682 = a17680 & a16198;
assign c1 = 1;
assign a5374 = ~a5372 & ~a5364;
assign a16196 = a16194 & a16186;
assign a18514 = a18512 & i154;
assign na18518 = ~a18518;
assign a18520 = ~a18508 & ~a9064;
assign a18542 = a18540 & a18526;
assign a18556 = ~a18554 & ~a18514;
assign a18562 = a18560 & a5408;
assign a19756 = ~a19754 & ~a18740;
assign a19892 = a19890 & ~a19862;
assign na8812 = ~a8812;
assign a19894 = ~a8802 & a8432;
assign a19900 = ~a19898 & ~a19896;
assign a16186 = ~a16184 & a14378;
assign a21664 = a21662 & ~a21660;
assign a23736 = ~a23734 & ~a22678;
assign a23742 = a23740 & ~l944;
assign z0 = l924;
assign a8150 = ~a8148 & i236;
assign a24056 = a24054 & ~a23936;
assign a24188 = a24186 & ~a24074;
assign a24322 = a24320 & ~a24208;
assign a24450 = a24448 & ~a24336;
assign a24582 = a24580 & ~a24468;
assign a24714 = a24712 & ~a24600;
assign a24846 = a24844 & ~a24732;
assign a24974 = a24972 & ~a24860;
assign a25106 = a25104 & ~a24990;
assign a25236 = a25234 & ~a25122;
assign na25240 = ~a25240;
assign a25242 = a12730 & i240;
assign na25818 = ~a25818;
assign na19408 = ~a19408;
assign a5352 = ~a5350 & ~a2782;
assign z1 = l980;
assign a25838 = ~a25836 & ~a25828;
assign a25846 = ~a25844 & ~a16220;
assign a25850 = ~a25848 & ~a25828;
assign a25852 = ~a16220 & ~l990;
assign na26072 = ~a26072;
assign na20174 = ~a20174;
assign na26078 = ~a26078;
assign na26106 = ~a26106;
assign na26594 = ~a26594;
assign na2536 = ~a2536;
assign na2752 = ~a2752;
assign na2516 = ~a2516;
assign na26612 = ~a26612;
assign a28188 = a28186 & ~a28022;
assign a28194 = ~a28192 & ~a28190;
assign a28236 = ~a28234 & ~a28196;
assign a20078 = ~a20076 & ~a20058;
assign a18850 = ~a18848 & ~a18846;
assign a28448 = ~a28446 & ~a17470;
assign a16250 = ~a16248 & ~a16240;
assign na28452 = ~a28452;
assign na25504 = ~a25504;
assign na25804 = ~a25804;
assign a25534 = ~a25532 & ~a25512;
assign na28462 = ~a28462;
assign a25578 = ~a25576 & ~a25544;
assign a28706 = ~a28704 & ~a17488;
assign a18924 = ~a18922 & ~a18920;
assign a28944 = ~a28942 & ~a17512;
assign a19004 = ~a19002 & ~a19000;
assign a29210 = ~a29208 & ~a17536;
assign a19086 = ~a19084 & ~a19082;
assign a29462 = ~a29460 & ~a17560;
assign a19168 = ~a19166 & ~a19164;
assign a29508 = ~a29506 & ~a17584;
assign na19250 = ~a19250;
assign a29548 = ~a29546 & ~a17610;
assign na19332 = ~a19332;
assign na29552 = ~a29552;
assign a25628 = ~a25626 & ~a25594;
assign na29562 = ~a29562;
assign na29572 = ~a29572;
assign a25672 = ~a25670 & ~a25644;
assign na29582 = ~a29582;
assign na25716 = ~a25716;
assign na29592 = ~a29592;
assign na25760 = ~a25760;
assign na29602 = ~a29602;
assign a29642 = ~a29640 & ~a17446;
assign na16278 = ~a16278;
assign na29646 = ~a29646;
assign na29650 = ~a29650;
assign na29654 = ~a29654;
assign na29658 = ~a29658;
assign na29662 = ~a29662;
assign a16608 = ~a16606 & ~a16598;
assign a29722 = ~a29720 & ~a29664;
assign a20054 = ~a20052 & ~a20034;
assign z2 = l908;
assign a29728 = ~a29726 & ~a29724;
assign a16712 = ~a16710 & ~a16702;
assign a29788 = ~a29786 & ~a29730;
assign a20028 = ~a20026 & ~a20008;
assign a29794 = ~a29792 & ~a29790;
assign a16816 = ~a16814 & ~a16806;
assign a29854 = ~a29852 & ~a29796;
assign a20002 = ~a20000 & ~a19982;
assign a29860 = ~a29858 & ~a29856;
assign a16920 = ~a16918 & ~a16910;
assign a29920 = ~a29918 & ~a29862;
assign a19976 = ~a19974 & ~a19956;
assign a29926 = ~a29924 & ~a29922;
assign na17016 = ~a17016;
assign a29986 = ~a29984 & ~a29928;
assign na19950 = ~a19950;
assign na29992 = ~a29992;
assign na17112 = ~a17112;
assign na30052 = ~a30052;
assign na19922 = ~a19922;
assign na30058 = ~a30058;
assign na8954 = ~a8954;
assign na30072 = ~a30072;
assign a31018 = a31016 & ~a30900;
assign a31020 = ~a17476 & ~a5360;
assign a31040 = ~a31038 & ~a31030;
assign na31048 = ~a31048;
assign a8946 = ~a8944 & ~a8908;
assign na8986 = ~a8986;
assign na31060 = ~a31060;
assign na31072 = ~a31072;
assign na31086 = ~a31086;
assign na8924 = ~a8924;
assign na8870 = ~a8870;
assign a31088 = ~a8430 & l930;
assign na31092 = ~a31092;
assign z3 = l884;
assign na31152 = ~a31152;
assign na18526 = ~a18526;
assign a31160 = ~a31158 & ~a18514;
assign na17784 = ~a17784;
assign z4 = l892;
assign na31102 = ~a31102;
assign na31176 = ~a31176;
assign a31182 = ~a31180 & ~a31178;
assign a8970 = ~a8968 & ~a8948;
assign na31110 = ~a31110;
assign na31202 = ~a31202;
assign a31208 = ~a31206 & ~a31204;
assign a9006 = ~a9004 & ~a8972;
assign na31118 = ~a31118;
assign na31222 = ~a31222;
assign na31228 = ~a31228;
assign na8906 = ~a8906;
assign a32370 = a32368 & a18508;
assign a32380 = a32378 & ~a18514;
assign na12366 = ~a12366;
assign na32396 = ~a32396;
assign a32386 = ~a32384 & ~a18514;
assign na32402 = ~a32402;
assign na12312 = ~a12312;
assign na32408 = ~a32408;
assign na32414 = ~a32414;
assign na12250 = ~a12250;
assign na32420 = ~a32420;
assign na32426 = ~a32426;
assign na12190 = ~a12190;
assign na32432 = ~a32432;
assign na32438 = ~a32438;
assign na16376 = ~a16376;
assign na17092 = ~a17092;
assign na18282 = ~a18282;
assign a16996 = ~a16994 & a16986;
assign na18208 = ~a18208;
assign a16892 = ~a16890 & a16882;
assign na18134 = ~a18134;
assign a16788 = ~a16786 & a16778;
assign na18060 = ~a18060;
assign a16684 = ~a16682 & a16674;
assign na17986 = ~a17986;
assign a16580 = ~a16578 & a16570;
assign na17912 = ~a17912;
assign a16514 = ~a16512 & a16504;
assign na17844 = ~a17844;
assign na32454 = ~a32454;
assign a32470 = ~a32468 & ~a8972;
assign a32486 = ~a32484 & ~a8948;
assign na22814 = ~a22814;
assign na22822 = ~a22822;
assign na22834 = ~a22834;
assign na22842 = ~a22842;
assign na22854 = ~a22854;
assign na22862 = ~a22862;
assign na22878 = ~a22878;
assign na22886 = ~a22886;
assign na22898 = ~a22898;
assign na22906 = ~a22906;
assign na21710 = ~a21710;
assign na21720 = ~a21720;
assign na21740 = ~a21740;
assign na21752 = ~a21752;
assign na21766 = ~a21766;
assign na21776 = ~a21776;
assign a21800 = ~a21798 & ~a21796;
assign a21810 = ~a21808 & ~a21806;
assign a21828 = ~a21826 & ~a21824;
assign na21840 = ~a21840;
assign na21886 = ~a21886;
assign na21894 = ~a21894;
assign na21906 = ~a21906;
assign na21914 = ~a21914;
assign na21926 = ~a21926;
assign na21934 = ~a21934;
assign a21950 = ~a21948 & ~a21946;
assign a21958 = ~a21956 & ~a21954;
assign a21970 = ~a21968 & ~a21966;
assign na21978 = ~a21978;
assign na22020 = ~a22020;
assign na22028 = ~a22028;
assign na22040 = ~a22040;
assign na22048 = ~a22048;
assign na22060 = ~a22060;
assign na22068 = ~a22068;
assign a22084 = ~a22082 & ~a22080;
assign a22092 = ~a22090 & ~a22088;
assign a22104 = ~a22102 & ~a22100;
assign na22112 = ~a22112;
assign na22154 = ~a22154;
assign na22162 = ~a22162;
assign na22174 = ~a22174;
assign na22182 = ~a22182;
assign na22194 = ~a22194;
assign na22202 = ~a22202;
assign a22218 = ~a22216 & ~a22214;
assign a22226 = ~a22224 & ~a22222;
assign a22238 = ~a22236 & ~a22234;
assign na22246 = ~a22246;
assign na22288 = ~a22288;
assign na22296 = ~a22296;
assign na22308 = ~a22308;
assign na22316 = ~a22316;
assign na22328 = ~a22328;
assign na22336 = ~a22336;
assign a22352 = ~a22350 & ~a22348;
assign a22360 = ~a22358 & ~a22356;
assign a22372 = ~a22370 & ~a22368;
assign na22380 = ~a22380;
assign na22422 = ~a22422;
assign na22430 = ~a22430;
assign na22442 = ~a22442;
assign na22450 = ~a22450;
assign na22462 = ~a22462;
assign na22470 = ~a22470;
assign a22486 = ~a22484 & ~a22482;
assign a22494 = ~a22492 & ~a22490;
assign a22506 = ~a22504 & ~a22502;
assign na22514 = ~a22514;
assign na22556 = ~a22556;
assign na22564 = ~a22564;
assign na22576 = ~a22576;
assign na22584 = ~a22584;
assign na22596 = ~a22596;
assign na22604 = ~a22604;
assign a22620 = ~a22618 & ~a22616;
assign a22628 = ~a22626 & ~a22624;
assign na22640 = ~a22640;
assign na22648 = ~a22648;
assign na26200 = ~a26200;
assign na26238 = ~a26238;
assign na26282 = ~a26282;
assign na26326 = ~a26326;
assign na26370 = ~a26370;
assign na26414 = ~a26414;
assign a32504 = ~a32502 & ~a32488;
assign a32508 = a32506 & i366;
assign a32538 = a32536 & ~a32510;
assign a16440 = ~a16438 & ~a16436;
assign na33374 = ~a33374;
assign na33380 = ~a33380;
assign na33402 = ~a33402;
assign na33408 = ~a33408;
assign a33430 = ~a33428 & ~a33410;
assign na33436 = ~a33436;
assign a33458 = ~a33456 & ~a33438;
assign na33464 = ~a33464;
assign a32966 = a32964 & l968;
assign na33468 = ~a33468;
assign a32978 = a32976 & a25236;
assign na33506 = ~a33506;
assign na33526 = ~a33526;
assign a31042 = a21692 & a16378;
assign na24030 = ~a24030;
assign na33570 = ~a33570;
assign na33624 = ~a33624;
assign na33636 = ~a33636;
assign na33642 = ~a33642;
assign na33652 = ~a33652;
assign a34176 = a34174 & ~a34096;
assign a32998 = a32996 & a24974;
assign z5 = l1516;
assign na23774 = ~a23774;
assign na24826 = ~a24826;
assign na34252 = ~a34252;
assign na34268 = ~a34268;
assign na34290 = ~a34290;
assign na34308 = ~a34308;
assign na34326 = ~a34326;
assign na25216 = ~a25216;
assign a34338 = ~a34336 & ~a34328;
assign na24954 = ~a24954;
assign na34350 = ~a34350;
assign a34362 = ~a34360 & ~a34354;
assign na24694 = ~a24694;
assign na24562 = ~a24562;
assign na24430 = ~a24430;
assign na24302 = ~a24302;
assign na24168 = ~a24168;
assign na24036 = ~a24036;
assign na25086 = ~a25086;
assign a33014 = a33012 & a24846;
assign a33032 = a33030 & a24714;
assign a33046 = a33044 & a24582;
assign a33066 = a33064 & a24450;
assign a33078 = a33076 & a24322;
assign a33094 = a33092 & a24188;
assign a33106 = a33104 & a24056;
assign na34374 = ~a34374;
assign na34380 = ~a34380;
assign na34386 = ~a34386;
assign na34392 = ~a34392;
assign na34398 = ~a34398;
assign na34404 = ~a34404;
assign na34410 = ~a34410;
assign na34416 = ~a34416;
assign na34422 = ~a34422;
assign na34428 = ~a34428;
assign na34440 = ~a34440;
assign na34446 = ~a34446;
assign na34452 = ~a34452;
assign na34458 = ~a34458;
assign na34464 = ~a34464;
assign na34470 = ~a34470;
assign na34476 = ~a34476;
assign na34482 = ~a34482;
assign a34488 = ~a34486 & ~a34484;
assign a34494 = ~a34492 & ~a34490;
assign na34506 = ~a34506;
assign na34512 = ~a34512;
assign na34518 = ~a34518;
assign na34524 = ~a34524;
assign na34530 = ~a34530;
assign na34536 = ~a34536;
assign na34542 = ~a34542;
assign na34548 = ~a34548;
assign a34554 = ~a34552 & ~a34550;
assign a34560 = ~a34558 & ~a34556;
assign na34572 = ~a34572;
assign na34578 = ~a34578;
assign na34584 = ~a34584;
assign na34590 = ~a34590;
assign na34596 = ~a34596;
assign na34602 = ~a34602;
assign na34608 = ~a34608;
assign na34614 = ~a34614;
assign a34620 = ~a34618 & ~a34616;
assign a34626 = ~a34624 & ~a34622;
assign na34638 = ~a34638;
assign na34644 = ~a34644;
assign na34650 = ~a34650;
assign na34656 = ~a34656;
assign na34662 = ~a34662;
assign na34668 = ~a34668;
assign na34674 = ~a34674;
assign na34680 = ~a34680;
assign a34686 = ~a34684 & ~a34682;
assign a34692 = ~a34690 & ~a34688;
assign na34704 = ~a34704;
assign na34710 = ~a34710;
assign na34716 = ~a34716;
assign na34722 = ~a34722;
assign na34728 = ~a34728;
assign na34734 = ~a34734;
assign na34740 = ~a34740;
assign na34746 = ~a34746;
assign a34752 = ~a34750 & ~a34748;
assign a34758 = ~a34756 & ~a34754;
assign na34770 = ~a34770;
assign na34776 = ~a34776;
assign na34782 = ~a34782;
assign na34788 = ~a34788;
assign na34794 = ~a34794;
assign na34800 = ~a34800;
assign na34806 = ~a34806;
assign na34812 = ~a34812;
assign a34818 = ~a34816 & ~a34814;
assign na34824 = ~a34824;
assign na34836 = ~a34836;
assign na34842 = ~a34842;
assign na34848 = ~a34848;
assign na34854 = ~a34854;
assign na34860 = ~a34860;
assign na34866 = ~a34866;
assign na34872 = ~a34872;
assign na34878 = ~a34878;
assign na34884 = ~a34884;
assign na34890 = ~a34890;
assign a34894 = ~a34892 & ~a14378;
assign z6 = l1196;
assign z7 = l1760;
assign z8 = l1762;
assign na17454 = ~a17454;
assign a34896 = ~a17494 & ~a5360;
assign a34898 = ~a17518 & ~a5360;
assign a34900 = ~a17542 & ~a5360;
assign a34902 = ~a17566 & ~a5360;
assign na17592 = ~a17592;
assign a34904 = ~a17616 & ~a5360;
assign a34910 = ~a34908 & ~a34906;
assign a21670 = ~a21668 & ~a21666;
assign na34920 = ~a34920;
assign na34928 = ~a34928;
assign na34936 = ~a34936;
assign na34946 = ~a34946;
assign na34954 = ~a34954;
assign na34962 = ~a34962;
assign na34970 = ~a34970;
assign na34976 = ~a34976;
assign a34988 = ~a34986 & ~a34978;
assign a21880 = ~a21878 & ~a21876;
assign na34994 = ~a34994;
assign a35000 = ~a34998 & ~a34996;
assign na35006 = ~a35006;
assign na35012 = ~a35012;
assign na35018 = ~a35018;
assign na35024 = ~a35024;
assign na35030 = ~a35030;
assign na35036 = ~a35036;
assign na35042 = ~a35042;
assign a35054 = ~a35052 & ~a35044;
assign a22014 = ~a22012 & ~a22010;
assign na35060 = ~a35060;
assign a35066 = ~a35064 & ~a35062;
assign na35072 = ~a35072;
assign na35078 = ~a35078;
assign na35084 = ~a35084;
assign na35090 = ~a35090;
assign na35096 = ~a35096;
assign na35102 = ~a35102;
assign na35108 = ~a35108;
assign a35120 = ~a35118 & ~a35110;
assign a22148 = ~a22146 & ~a22144;
assign na35126 = ~a35126;
assign a35132 = ~a35130 & ~a35128;
assign na35138 = ~a35138;
assign na35144 = ~a35144;
assign na35150 = ~a35150;
assign na35156 = ~a35156;
assign na35162 = ~a35162;
assign na35168 = ~a35168;
assign na35174 = ~a35174;
assign a35186 = ~a35184 & ~a35176;
assign a22282 = ~a22280 & ~a22278;
assign na35192 = ~a35192;
assign a35198 = ~a35196 & ~a35194;
assign na35204 = ~a35204;
assign na35210 = ~a35210;
assign na35216 = ~a35216;
assign na35222 = ~a35222;
assign na35228 = ~a35228;
assign na35234 = ~a35234;
assign na35240 = ~a35240;
assign a35252 = ~a35250 & ~a35242;
assign a22416 = ~a22414 & ~a22412;
assign na35258 = ~a35258;
assign a35264 = ~a35262 & ~a35260;
assign na35270 = ~a35270;
assign na35276 = ~a35276;
assign na35282 = ~a35282;
assign na35288 = ~a35288;
assign na35294 = ~a35294;
assign na35300 = ~a35300;
assign na35306 = ~a35306;
assign na35318 = ~a35318;
assign a22550 = ~a22548 & ~a22546;
assign na35324 = ~a35324;
assign a35330 = ~a35328 & ~a35326;
assign na35336 = ~a35336;
assign na35342 = ~a35342;
assign na35348 = ~a35348;
assign na35354 = ~a35354;
assign na35360 = ~a35360;
assign na35366 = ~a35366;
assign na35372 = ~a35372;
assign na35386 = ~a35386;
assign a22808 = ~a22806 & ~a22804;
assign na35392 = ~a35392;
assign na35398 = ~a35398;
assign na35404 = ~a35404;
assign na35410 = ~a35410;
assign na35416 = ~a35416;
assign na35422 = ~a35422;
assign na35428 = ~a35428;
assign na35434 = ~a35434;
assign na35440 = ~a35440;
assign a35472 = a35470 & ~a35460;
assign na8846 = ~a8846;
assign na8836 = ~a8836;
assign na8860 = ~a8860;
assign na8826 = ~a8826;
assign a35514 = a35512 & ~a35500;
assign a35554 = a35552 & ~a35544;
assign a35588 = a35586 & ~a35578;
assign a35636 = a35634 & ~a35626;
assign a35664 = a35662 & ~a35650;
assign a35700 = a35698 & ~a35690;
assign a35720 = a35718 & ~a35712;
assign a35748 = a35746 & ~a35738;
assign na35754 = ~a35754;
assign na35760 = ~a35760;
assign na35766 = ~a35766;
assign na35772 = ~a35772;
assign na35778 = ~a35778;
assign na35784 = ~a35784;
assign na35790 = ~a35790;
assign na35796 = ~a35796;
assign na35802 = ~a35802;
assign a32592 = a32590 & l966;
assign a32634 = a32632 & l964;
assign a32680 = a32678 & l962;
assign a32722 = a32720 & l960;
assign a32772 = a32770 & a5606;
assign a32814 = a32812 & a5600;
assign a32860 = a32858 & a5594;
assign a32908 = a32906 & a5568;
assign a33156 = ~a33154 & l968;
assign a33198 = a33196 & l970;
assign na35828 = ~a35828;
assign z9 = l1216;
assign z10 = l1200;
assign z11 = l1176;
assign z12 = l1232;
assign na35836 = ~a35836;
assign na35856 = ~a35856;
assign na35862 = ~a35862;
assign na35880 = ~a35880;
assign na35886 = ~a35886;
assign na35896 = ~a35896;
assign na35902 = ~a35902;
assign na35912 = ~a35912;
assign na35922 = ~a35922;
assign na18744 = ~a18744;
assign a35930 = a35928 & ~l926;
assign z13 = l1190;
assign a35946 = a35944 & ~a14378;
assign a35960 = a35958 & ~a14378;
assign a35968 = a35966 & ~l980;
assign na36056 = ~a36056;
assign na37126 = ~a37126;
assign na37160 = ~a37160;
assign na37184 = ~a37184;
assign na37206 = ~a37206;
assign na37222 = ~a37222;
assign na37246 = ~a37246;
assign na37266 = ~a37266;
assign na37386 = ~a37386;
assign na37400 = ~a37400;
assign na37448 = ~a37448;
assign na37476 = ~a37476;
assign na37482 = ~a37482;
assign a41638 = a41636 & ~a41522;
assign a41644 = ~a41642 & ~a41640;
assign na41660 = ~a41660;
assign a41670 = a41668 & ~i674;
assign a41672 = i678 & ~i674;
assign na41678 = ~a41678;
assign a41736 = a41734 & ~a41680;
assign na41742 = ~a41742;
assign na41800 = ~a41800;
assign na41806 = ~a41806;
assign na41846 = ~a41846;
assign a44408 = a44406 & ~a42234;
assign a44428 = ~a44426 & ~a44424;
assign a41654 = ~a41652 & ~a41646;
assign a44442 = ~a44440 & ~a44438;
assign a44450 = ~a44448 & ~a44446;
assign a44462 = ~a44460 & ~a44458;
assign a44472 = ~a44470 & ~a44468;
assign a44482 = ~a44480 & ~a44478;
assign a44490 = ~a44488 & ~a44486;
assign a44498 = ~a44496 & ~a44494;
assign a44506 = ~a44504 & ~a44502;
assign a44514 = ~a44512 & ~a44510;
assign a44520 = ~a44518 & ~a44516;
assign a44526 = ~a44524 & ~a44522;
assign a44532 = ~a44530 & ~a44528;
assign a44538 = ~a44536 & ~a44534;
assign a44544 = ~a44542 & ~a44540;
assign a44550 = ~a44548 & ~a44546;
assign a44556 = ~a44554 & ~a44552;
assign a44562 = ~a44560 & ~a44558;
assign a44568 = ~a44566 & ~a44564;
assign a44574 = ~a44572 & ~a44570;
assign a44580 = ~a44578 & ~a44576;
assign a44586 = ~a44584 & ~a44582;
assign a44592 = ~a44590 & ~a44588;
assign a44598 = ~a44596 & ~a44594;
assign a44604 = ~a44602 & ~a44600;
assign a44610 = ~a44608 & ~a44606;
assign a44616 = ~a44614 & ~a44612;
assign a44622 = ~a44620 & ~a44618;
assign a44628 = ~a44626 & ~a44624;
assign a44634 = ~a44632 & ~a44630;
assign a44640 = ~a44638 & ~a44636;
assign a44646 = ~a44644 & ~a44642;
assign a44652 = ~a44650 & ~a44648;
assign a44658 = ~a44656 & ~a44654;
assign a44664 = ~a44662 & ~a44660;
assign a44670 = ~a44668 & ~a44666;
assign a44676 = ~a44674 & ~a44672;
assign a44682 = ~a44680 & ~a44678;
assign a44688 = ~a44686 & ~a44684;
assign a44694 = ~a44692 & ~a44690;
assign a44700 = ~a44698 & ~a44696;
assign a44706 = ~a44704 & ~a44702;
assign a44712 = ~a44710 & ~a44708;
assign a44718 = ~a44716 & ~a44714;
assign a44724 = ~a44722 & ~a44720;
assign a44730 = ~a44728 & ~a44726;
assign a44736 = ~a44734 & ~a44732;
assign a44742 = ~a44740 & ~a44738;
assign a44748 = ~a44746 & ~a44744;
assign a44754 = ~a44752 & ~a44750;
assign a44760 = ~a44758 & ~a44756;
assign a44766 = ~a44764 & ~a44762;
assign a44772 = ~a44770 & ~a44768;
assign a44778 = ~a44776 & ~a44774;
assign a44784 = ~a44782 & ~a44780;
assign a44790 = ~a44788 & ~a44786;
assign a44796 = ~a44794 & ~a44792;
assign a44802 = ~a44800 & ~a44798;
assign a44808 = ~a44806 & ~a44804;
assign a44814 = ~a44812 & ~a44810;
assign a44834 = a44832 & ~a44816;
assign a45596 = a45594 & ~i650;
assign na8818 = ~a8818;
assign z14 = l2120;
assign a8814 = ~l1172 & l928;
assign z15 = l2256;
assign z16 = l1172;
assign z17 = l2266;
assign na40992 = ~a40992;
assign na45602 = ~a45602;
assign a45608 = ~a45606 & ~a45604;
assign a40642 = ~a40640 & ~a37484;
assign z18 = l2124;
assign a45622 = a45620 & ~a45610;
assign a46176 = a46174 & ~a45948;
assign a48022 = a48020 & ~a47876;
assign a48034 = a48032 & ~a48026;
assign a48048 = a48046 & ~a48040;
assign na48062 = ~a48062;
assign a48584 = a48582 & ~a48504;
assign a48590 = ~a48588 & ~a48586;
assign a48596 = ~a48594 & ~a48592;
assign a48602 = ~a48600 & ~a48598;
assign a48608 = ~a48606 & ~a48604;
assign a48614 = ~a48612 & ~a48610;
assign a48620 = ~a48618 & ~a48616;
assign a48626 = ~a48624 & ~a48622;
assign a48632 = ~a48630 & ~a48628;
assign a48638 = ~a48636 & ~a48634;
assign a48644 = ~a48642 & ~a48640;
assign a48650 = ~a48648 & ~a48646;
assign a48656 = ~a48654 & ~a48652;
assign a48662 = ~a48660 & ~a48658;
assign a48668 = ~a48666 & ~a48664;
assign a48674 = ~a48672 & ~a48670;
assign a48680 = ~a48678 & ~a48676;
assign a48686 = ~a48684 & ~a48682;
assign a48692 = ~a48690 & ~a48688;
assign a48698 = ~a48696 & ~a48694;
assign a48704 = ~a48702 & ~a48700;
assign a48728 = a48726 & ~a48706;
assign a48792 = a48790 & ~i650;
assign a48808 = a48806 & ~a48794;
assign a49932 = a49930 & ~a49684;
assign na49946 = ~a49946;
assign na49958 = ~a49958;
assign a49740 = a49738 & ~a49724;
assign a49996 = a49994 & ~i650;
assign a49758 = a49756 & ~a49746;
assign a50024 = a50022 & ~a50000;
assign a49784 = a49782 & ~a49764;
assign a50066 = a50064 & ~a50026;
assign a50084 = ~a50082 & ~a50076;
assign a49802 = ~a49800 & a49798;
assign a50114 = ~a50112 & ~a50110;
assign a49824 = ~a49822 & a49820;
assign a49842 = a49840 & ~a49830;
assign a50136 = a50134 & ~a50116;
assign a49862 = a49860 & ~a49848;
assign a50164 = a50162 & ~a50138;
assign a49880 = a49878 & ~a49868;
assign a50176 = a50174 & ~a50170;
assign z19 = l2270;
assign z20 = l2284;
assign z21 = l2272;
assign z22 = l2296;
assign na50182 = ~a50182;
assign na50188 = ~a50188;
assign na50194 = ~a50194;
assign na50200 = ~a50200;
assign na50248 = ~a50248;
assign na50254 = ~a50254;
assign na50260 = ~a50260;
assign na50266 = ~a50266;
assign na50272 = ~a50272;
assign na50278 = ~a50278;
assign na50284 = ~a50284;
assign a50346 = ~a50344 & ~a50342;
assign a50420 = ~a50418 & ~a50416;
assign na50426 = ~a50426;
assign a50620 = ~a50618 & ~a50574;
assign a50646 = ~a50644 & ~a50642;
assign a50672 = ~a50670 & ~a50668;
assign a50698 = ~a50696 & ~a50694;
assign a50724 = ~a50722 & ~a50720;
assign a50750 = ~a50748 & ~a50746;
assign a50776 = ~a50774 & ~a50772;
assign a50802 = ~a50800 & ~a50798;
assign a50828 = ~a50826 & ~a50824;
assign a50854 = ~a50852 & ~a50850;
assign na50954 = ~a50954;
assign na50958 = ~a50958;
assign na50962 = ~a50962;
assign na50970 = ~a50970;
assign a50972 = a16186 & ~l2480;
assign na18534 = ~a18534;
assign a50986 = ~a50984 & ~l924;
assign a50990 = ~a50988 & ~l924;
assign na50996 = ~a50996;
assign a51000 = ~a50998 & ~l2488;
assign a5624 = a5622 & ~a5568;
assign z23 = l2094;
assign z24 = l1148;
assign z25 = l1162;
assign z26 = l1166;
assign z27 = l1164;
assign a2502 = l882 & ~l880;
assign a2504 = ~a2502 & ~l1536;
assign a2506 = l1004 & l880;
assign a2508 = a2506 & l1002;
assign a2510 = l1006 & ~l880;
assign a2512 = ~a2510 & ~a2508;
assign a2514 = ~a2512 & l882;
assign a2516 = ~a2514 & ~l1008;
assign a2518 = ~a2516 & ~l1244;
assign a2520 = a2516 & l1244;
assign a2522 = ~a2520 & ~a2518;
assign a2524 = l1002 & ~l880;
assign a2526 = a2506 & ~l1002;
assign a2528 = ~a2526 & ~a2524;
assign a2530 = ~l1004 & l1002;
assign a2532 = ~a2530 & a2528;
assign a2534 = ~a2532 & l882;
assign a2536 = ~a2534 & ~l1534;
assign a2538 = a2536 & l1156;
assign a2540 = ~a2538 & a2522;
assign a2542 = ~a2536 & ~l1156;
assign a2544 = ~a2542 & a2540;
assign a2546 = ~l1228 & l890;
assign a2548 = i4 & ~i2;
assign a2550 = ~a2548 & ~i2;
assign a2552 = i12 & ~i2;
assign a2554 = a2552 & a2550;
assign a2556 = ~a2550 & ~i12;
assign a2558 = ~a2556 & ~a2554;
assign a2560 = ~a2558 & ~i14;
assign a2562 = a2558 & i14;
assign a2564 = ~a2562 & ~a2560;
assign a2566 = ~a2554 & i16;
assign a2568 = ~a2566 & ~a2554;
assign a2570 = ~i8 & i2;
assign a2572 = a2570 & i12;
assign a2574 = a2572 & i18;
assign a2576 = a2574 & ~a2568;
assign a2578 = a2572 & ~i18;
assign a2580 = a2578 & a2568;
assign a2582 = ~a2580 & ~a2576;
assign a2584 = a2574 & a2568;
assign a2586 = a2578 & ~a2568;
assign a2588 = ~a2586 & ~a2584;
assign a2590 = i8 & i2;
assign a2592 = a2590 & i12;
assign a2594 = a2592 & i18;
assign a2596 = a2594 & ~a2568;
assign a2598 = a2592 & ~i18;
assign a2600 = a2598 & a2568;
assign a2602 = ~a2600 & ~a2596;
assign a2604 = a2552 & ~a2550;
assign a2606 = a2604 & i18;
assign a2608 = a2606 & ~a2568;
assign a2610 = a2604 & ~i18;
assign a2612 = a2610 & a2568;
assign a2614 = ~a2612 & ~a2608;
assign a2616 = a2614 & a2602;
assign a2618 = a2616 & a2582;
assign a2620 = a2618 & i20;
assign a2622 = ~a2620 & a2618;
assign a2624 = a2622 & ~a2588;
assign a2626 = a2616 & ~a2554;
assign a2628 = a2626 & a2582;
assign a2630 = ~a2622 & ~a2588;
assign a2632 = a2606 & a2568;
assign a2634 = a2610 & ~a2568;
assign a2636 = ~a2634 & ~a2632;
assign a2638 = ~a2636 & ~a2622;
assign a2640 = a2594 & a2568;
assign a2642 = a2598 & ~a2568;
assign a2644 = ~a2642 & ~a2640;
assign a2646 = ~a2644 & ~a2622;
assign a2648 = ~a2646 & a2602;
assign a2650 = a2648 & a2614;
assign a2652 = a2650 & ~a2638;
assign a2654 = a2652 & ~a2554;
assign a2656 = a2654 & a2582;
assign a2658 = a2656 & ~a2630;
assign a2660 = a2658 & i22;
assign a2662 = ~a2660 & a2628;
assign a2664 = a2662 & a2624;
assign a2666 = ~a2664 & a2582;
assign a2668 = ~a2644 & a2622;
assign a2670 = a2668 & a2662;
assign a2672 = ~a2670 & a2602;
assign a2674 = ~a2636 & a2622;
assign a2676 = a2674 & a2662;
assign a2678 = ~a2676 & a2614;
assign a2680 = a2678 & a2672;
assign a2682 = a2680 & a2666;
assign a2684 = ~a2662 & a2624;
assign a2686 = ~a2684 & ~a2630;
assign a2688 = a2668 & ~a2662;
assign a2690 = ~a2688 & ~a2646;
assign a2692 = a2674 & ~a2662;
assign a2694 = ~a2692 & ~a2638;
assign a2696 = a2694 & a2690;
assign a2698 = a2696 & a2686;
assign a2700 = a2698 & a2682;
assign a2702 = ~a2700 & ~i14;
assign a2704 = ~i12 & ~i2;
assign a2706 = a2704 & a2550;
assign a2708 = ~a2706 & i14;
assign a2710 = ~a2708 & ~a2702;
assign a2712 = a2710 & a2564;
assign a2714 = ~a2564 & ~i92;
assign a2716 = a2564 & i92;
assign a2718 = ~a2716 & ~a2714;
assign a2720 = ~a2710 & ~i92;
assign a2722 = ~a2710 & ~a2564;
assign a2724 = ~a2722 & ~a2712;
assign a2726 = a2724 & i92;
assign a2728 = ~a2726 & ~a2720;
assign a2730 = a2728 & a2718;
assign a2732 = ~a2728 & ~a2718;
assign a2734 = ~a2732 & ~a2730;
assign a2736 = ~a2734 & ~a2712;
assign a2738 = a2736 & ~l890;
assign a2740 = ~a2738 & ~a2546;
assign a2742 = ~l1006 & l880;
assign a2744 = a2742 & ~l1004;
assign a2746 = l1004 & ~l880;
assign a2748 = ~a2746 & ~a2744;
assign a2750 = ~a2748 & l882;
assign a2752 = ~a2750 & ~l1538;
assign a2754 = a2752 & ~a2740;
assign a2756 = ~a2754 & a2544;
assign a2758 = ~a2752 & a2740;
assign a2760 = ~a2758 & a2756;
assign a2762 = ~l1212 & l890;
assign a2764 = a2718 & ~a2712;
assign a2766 = a2764 & ~l890;
assign a2768 = ~a2766 & ~a2762;
assign a2770 = ~a2768 & a2504;
assign a2772 = ~a2770 & a2760;
assign a2774 = a2768 & ~a2504;
assign a2776 = ~a2774 & a2772;
assign a2778 = ~a2776 & l1540;
assign a2780 = ~a2778 & ~l884;
assign a2782 = l890 & ~l888;
assign a2784 = ~a2550 & i6;
assign a2786 = a2570 & i10;
assign a2788 = i32 & i30;
assign a2790 = a2788 & i28;
assign a2792 = a2790 & i26;
assign a2794 = a2792 & i24;
assign a2796 = ~i36 & ~i34;
assign a2798 = ~a2796 & a2794;
assign a2800 = ~a2798 & ~i38;
assign a2802 = a2550 & i42;
assign a2804 = a2802 & i44;
assign a2806 = a2804 & i46;
assign a2808 = a2806 & i48;
assign a2810 = a2808 & i50;
assign a2812 = ~a2550 & i52;
assign a2814 = ~a2812 & ~a2810;
assign a2816 = a2814 & i40;
assign a2818 = ~a2816 & a2550;
assign a2820 = a2570 & i42;
assign a2822 = a2820 & i44;
assign a2824 = a2822 & i46;
assign a2826 = a2824 & i48;
assign a2828 = a2826 & i50;
assign a2830 = a2590 & i42;
assign a2832 = a2830 & i44;
assign a2834 = a2832 & i46;
assign a2836 = a2834 & i48;
assign a2838 = a2836 & i50;
assign a2840 = a2548 & i42;
assign a2842 = a2840 & i44;
assign a2844 = a2842 & i46;
assign a2846 = a2844 & i48;
assign a2848 = a2846 & i50;
assign a2850 = ~a2848 & ~a2838;
assign a2852 = a2850 & ~a2828;
assign a2854 = a2550 & i56;
assign a2856 = ~a2854 & a2852;
assign a2858 = a2856 & i54;
assign a2860 = ~a2858 & ~a2550;
assign a2862 = ~a2860 & ~a2818;
assign a2864 = ~a2862 & a2560;
assign a2866 = i62 & i38;
assign a2868 = a2866 & i60;
assign a2870 = ~a2868 & i58;
assign a2872 = a2868 & ~i58;
assign a2874 = ~a2872 & ~a2870;
assign a2876 = ~a2874 & ~a2798;
assign a2878 = ~a2876 & a2864;
assign a2880 = a2560 & ~i42;
assign a2882 = a2868 & i58;
assign a2884 = ~a2882 & i36;
assign a2886 = ~a2884 & ~a2798;
assign a2888 = a2882 & ~i36;
assign a2890 = ~a2888 & a2886;
assign a2892 = a2890 & a2864;
assign a2894 = a2882 & i36;
assign a2896 = ~a2894 & i34;
assign a2898 = a2894 & ~i34;
assign a2900 = ~a2898 & ~a2896;
assign a2902 = ~a2900 & ~a2798;
assign a2904 = ~a2902 & a2864;
assign a2906 = a2894 & i34;
assign a2908 = ~a2906 & i30;
assign a2910 = ~a2908 & ~a2798;
assign a2912 = a2906 & ~i30;
assign a2914 = ~a2912 & a2910;
assign a2916 = a2560 & ~i50;
assign a2918 = ~a2916 & a2864;
assign a2920 = a2914 & a2864;
assign a2922 = a2906 & i30;
assign a2924 = ~a2922 & i32;
assign a2926 = ~a2924 & ~a2798;
assign a2928 = a2922 & ~i32;
assign a2930 = ~a2928 & a2926;
assign a2932 = a2560 & ~i48;
assign a2934 = ~a2932 & a2918;
assign a2936 = a2930 & a2864;
assign a2938 = a2922 & i32;
assign a2940 = ~a2938 & i28;
assign a2942 = ~a2940 & ~a2798;
assign a2944 = a2938 & ~i28;
assign a2946 = ~a2944 & a2942;
assign a2948 = a2560 & ~i46;
assign a2950 = ~a2948 & a2934;
assign a2952 = a2946 & a2864;
assign a2954 = a2938 & i28;
assign a2956 = ~a2954 & i26;
assign a2958 = ~a2956 & ~a2798;
assign a2960 = a2954 & ~i26;
assign a2962 = ~a2960 & a2958;
assign a2964 = a2560 & ~i44;
assign a2966 = ~a2964 & a2950;
assign a2968 = a2962 & a2864;
assign a2970 = a2954 & i26;
assign a2972 = a2970 & ~i24;
assign a2974 = ~a2972 & ~i24;
assign a2976 = a2966 & ~a2880;
assign a2978 = a2974 & a2864;
assign a2980 = ~a2978 & a2976;
assign a2982 = ~a2980 & ~a2974;
assign a2984 = ~a2982 & a2880;
assign a2986 = ~a2984 & ~a2968;
assign a2988 = a2982 & ~a2880;
assign a2990 = ~a2988 & ~a2986;
assign a2992 = ~a2990 & a2966;
assign a2994 = ~a2992 & ~a2962;
assign a2996 = ~a2994 & a2880;
assign a2998 = ~a2996 & ~a2952;
assign a3000 = a2994 & ~a2880;
assign a3002 = ~a3000 & ~a2998;
assign a3004 = ~a2916 & a2880;
assign a3006 = a3004 & ~a2932;
assign a3008 = a3006 & ~a2948;
assign a3010 = a3008 & ~a2964;
assign a3012 = a3010 & ~a2990;
assign a3014 = ~a3012 & a2982;
assign a3016 = ~a3014 & a2964;
assign a3018 = ~a3016 & ~a3002;
assign a3020 = a3014 & ~a2964;
assign a3022 = ~a3020 & ~a3018;
assign a3024 = ~a3022 & a2950;
assign a3026 = a3024 & a2946;
assign a3028 = ~a3024 & ~a2946;
assign a3030 = ~a3028 & ~a3026;
assign a3032 = a3030 & a2880;
assign a3034 = ~a3032 & ~a2936;
assign a3036 = ~a3030 & ~a2880;
assign a3038 = ~a3036 & ~a3034;
assign a3040 = ~a3022 & a3008;
assign a3042 = a3040 & ~a2994;
assign a3044 = ~a3040 & a2994;
assign a3046 = ~a3044 & ~a3042;
assign a3048 = ~a3046 & ~a3026;
assign a3050 = ~a3048 & a2964;
assign a3052 = ~a3050 & ~a3038;
assign a3054 = a3048 & ~a2964;
assign a3056 = ~a3054 & ~a3052;
assign a3058 = ~a3042 & a3014;
assign a3060 = a2964 & ~a2916;
assign a3062 = a3060 & ~a2932;
assign a3064 = a3062 & ~a2948;
assign a3066 = a3064 & ~a3022;
assign a3068 = ~a3066 & a3058;
assign a3070 = ~a3068 & a2948;
assign a3072 = ~a3070 & ~a3056;
assign a3074 = a3068 & ~a2948;
assign a3076 = ~a3074 & ~a3072;
assign a3078 = ~a3076 & a2934;
assign a3080 = ~a3078 & ~a2930;
assign a3082 = a3078 & a2930;
assign a3084 = ~a3082 & ~a3080;
assign a3086 = a3084 & a2880;
assign a3088 = ~a3086 & ~a2920;
assign a3090 = ~a3084 & ~a2880;
assign a3092 = ~a3090 & ~a3088;
assign a3094 = ~a3076 & a3006;
assign a3096 = a3094 & a3030;
assign a3098 = ~a3094 & ~a3030;
assign a3100 = ~a3098 & ~a3096;
assign a3102 = ~a3100 & ~a3082;
assign a3104 = a3100 & a3082;
assign a3106 = ~a3104 & ~a3102;
assign a3108 = a3106 & a2964;
assign a3110 = ~a3108 & ~a3092;
assign a3112 = ~a3106 & ~a2964;
assign a3114 = ~a3112 & ~a3110;
assign a3116 = ~a3076 & a3062;
assign a3118 = a3116 & ~a3048;
assign a3120 = ~a3116 & a3048;
assign a3122 = ~a3120 & ~a3118;
assign a3124 = ~a3096 & ~a3082;
assign a3126 = ~a3124 & ~a3098;
assign a3128 = ~a3126 & ~a3122;
assign a3130 = a3126 & a3122;
assign a3132 = ~a3130 & ~a3128;
assign a3134 = a3132 & a2948;
assign a3136 = ~a3134 & ~a3114;
assign a3138 = ~a3132 & ~a2948;
assign a3140 = ~a3138 & ~a3136;
assign a3142 = a2948 & ~a2916;
assign a3144 = a3142 & ~a2932;
assign a3146 = a3144 & ~a3076;
assign a3148 = ~a3146 & a3068;
assign a3150 = ~a3126 & ~a3118;
assign a3152 = ~a3150 & ~a3120;
assign a3154 = ~a3152 & a3148;
assign a3156 = ~a3154 & a2932;
assign a3158 = ~a3156 & ~a3140;
assign a3160 = a3154 & ~a2932;
assign a3162 = ~a3160 & ~a3158;
assign a3164 = ~a3162 & a2918;
assign a3166 = a3164 & a2914;
assign a3168 = ~a3164 & ~a2914;
assign a3170 = ~a3168 & ~a3166;
assign a3172 = a3170 & a2880;
assign a3174 = ~a3172 & ~a2904;
assign a3176 = ~a3170 & ~a2880;
assign a3178 = ~a3176 & ~a3174;
assign a3180 = ~a3162 & a3004;
assign a3182 = a3180 & a3084;
assign a3184 = ~a3180 & ~a3084;
assign a3186 = ~a3184 & ~a3182;
assign a3188 = ~a3186 & ~a3166;
assign a3190 = a3186 & a3166;
assign a3192 = ~a3190 & ~a3188;
assign a3194 = a3192 & a2964;
assign a3196 = ~a3194 & ~a3178;
assign a3198 = ~a3192 & ~a2964;
assign a3200 = ~a3198 & ~a3196;
assign a3202 = ~a3162 & a3060;
assign a3204 = a3202 & a3106;
assign a3206 = ~a3202 & ~a3106;
assign a3208 = ~a3206 & ~a3204;
assign a3210 = ~a3182 & ~a3166;
assign a3212 = ~a3210 & ~a3184;
assign a3214 = ~a3212 & ~a3208;
assign a3216 = a3212 & a3208;
assign a3218 = ~a3216 & ~a3214;
assign a3220 = a3218 & a2948;
assign a3222 = ~a3220 & ~a3200;
assign a3224 = ~a3218 & ~a2948;
assign a3226 = ~a3224 & ~a3222;
assign a3228 = ~a3162 & a3142;
assign a3230 = a3228 & a3132;
assign a3232 = ~a3228 & ~a3132;
assign a3234 = ~a3232 & ~a3230;
assign a3236 = ~a3212 & ~a3204;
assign a3238 = ~a3236 & ~a3206;
assign a3240 = ~a3238 & ~a3234;
assign a3242 = a3238 & a3234;
assign a3244 = ~a3242 & ~a3240;
assign a3246 = a3244 & a2932;
assign a3248 = ~a3246 & ~a3226;
assign a3250 = ~a3244 & ~a2932;
assign a3252 = ~a3250 & ~a3248;
assign a3254 = a2932 & ~a2916;
assign a3256 = a3254 & ~a3162;
assign a3258 = ~a3256 & a3154;
assign a3260 = ~a3238 & ~a3230;
assign a3262 = ~a3260 & ~a3232;
assign a3264 = ~a3262 & a3258;
assign a3266 = ~a3264 & a2916;
assign a3268 = ~a3266 & ~a3252;
assign a3270 = a3264 & ~a2916;
assign a3272 = ~a3270 & ~a3268;
assign a3274 = ~a3272 & a2864;
assign a3276 = a3274 & ~a2902;
assign a3278 = ~a3274 & a2902;
assign a3280 = ~a3278 & ~a3276;
assign a3282 = a3280 & a2880;
assign a3284 = ~a3282 & ~a2892;
assign a3286 = ~a3280 & ~a2880;
assign a3288 = ~a3286 & ~a3284;
assign a3290 = ~a3272 & a2880;
assign a3292 = ~a3290 & ~a3170;
assign a3294 = a3290 & a3170;
assign a3296 = ~a3294 & ~a3292;
assign a3298 = ~a3296 & ~a3276;
assign a3300 = a3296 & a3276;
assign a3302 = ~a3300 & ~a3298;
assign a3304 = a3302 & a2964;
assign a3306 = ~a3304 & ~a3288;
assign a3308 = ~a3302 & ~a2964;
assign a3310 = ~a3308 & ~a3306;
assign a3312 = ~a3272 & a2964;
assign a3314 = a3312 & a3192;
assign a3316 = ~a3312 & ~a3192;
assign a3318 = ~a3316 & ~a3314;
assign a3320 = ~a3294 & ~a3276;
assign a3322 = ~a3320 & ~a3292;
assign a3324 = ~a3322 & ~a3318;
assign a3326 = a3322 & a3318;
assign a3328 = ~a3326 & ~a3324;
assign a3330 = a3328 & a2948;
assign a3332 = ~a3330 & ~a3310;
assign a3334 = ~a3328 & ~a2948;
assign a3336 = ~a3334 & ~a3332;
assign a3338 = ~a3272 & a2948;
assign a3340 = a3338 & a3218;
assign a3342 = ~a3338 & ~a3218;
assign a3344 = ~a3342 & ~a3340;
assign a3346 = ~a3322 & ~a3314;
assign a3348 = ~a3346 & ~a3316;
assign a3350 = ~a3348 & ~a3344;
assign a3352 = a3348 & a3344;
assign a3354 = ~a3352 & ~a3350;
assign a3356 = a3354 & a2932;
assign a3358 = ~a3356 & ~a3336;
assign a3360 = ~a3354 & ~a2932;
assign a3362 = ~a3360 & ~a3358;
assign a3364 = ~a3272 & a2932;
assign a3366 = a3364 & a3244;
assign a3368 = ~a3364 & ~a3244;
assign a3370 = ~a3368 & ~a3366;
assign a3372 = ~a3348 & ~a3340;
assign a3374 = ~a3372 & ~a3342;
assign a3376 = ~a3374 & ~a3370;
assign a3378 = a3374 & a3370;
assign a3380 = ~a3378 & ~a3376;
assign a3382 = a3380 & a2916;
assign a3384 = ~a3382 & ~a3362;
assign a3386 = ~a3380 & ~a2916;
assign a3388 = ~a3386 & ~a3384;
assign a3390 = ~a3272 & a2916;
assign a3392 = ~a3390 & a3264;
assign a3394 = ~a3374 & ~a3366;
assign a3396 = ~a3394 & ~a3368;
assign a3398 = ~a3396 & a3392;
assign a3400 = ~a3398 & a3388;
assign a3402 = ~a3400 & a2864;
assign a3404 = a3402 & a2890;
assign a3406 = ~a3402 & ~a2890;
assign a3408 = ~a3406 & ~a3404;
assign a3410 = a3408 & a2880;
assign a3412 = ~a3410 & ~a2878;
assign a3414 = ~a3408 & ~a2880;
assign a3416 = ~a3414 & ~a3412;
assign a3418 = ~a3400 & a2880;
assign a3420 = ~a3418 & ~a3280;
assign a3422 = a3418 & a3280;
assign a3424 = ~a3422 & ~a3420;
assign a3426 = ~a3424 & ~a3404;
assign a3428 = a3424 & a3404;
assign a3430 = ~a3428 & ~a3426;
assign a3432 = a3430 & a2964;
assign a3434 = ~a3432 & ~a3416;
assign a3436 = ~a3430 & ~a2964;
assign a3438 = ~a3436 & ~a3434;
assign a3440 = ~a3422 & ~a3404;
assign a3442 = ~a3440 & ~a3420;
assign a3444 = ~a3400 & a2964;
assign a3446 = ~a3444 & ~a3302;
assign a3448 = a3444 & a3302;
assign a3450 = ~a3448 & ~a3446;
assign a3452 = ~a3450 & ~a3442;
assign a3454 = a3450 & a3442;
assign a3456 = ~a3454 & ~a3452;
assign a3458 = a3456 & a2948;
assign a3460 = ~a3458 & ~a3438;
assign a3462 = ~a3456 & ~a2948;
assign a3464 = ~a3462 & ~a3460;
assign a3466 = ~a3400 & a2948;
assign a3468 = a3466 & a3328;
assign a3470 = ~a3466 & ~a3328;
assign a3472 = ~a3470 & ~a3468;
assign a3474 = ~a3448 & ~a3442;
assign a3476 = ~a3474 & ~a3446;
assign a3478 = ~a3476 & ~a3472;
assign a3480 = a3476 & a3472;
assign a3482 = ~a3480 & ~a3478;
assign a3484 = a3482 & a2932;
assign a3486 = ~a3484 & ~a3464;
assign a3488 = ~a3482 & ~a2932;
assign a3490 = ~a3488 & ~a3486;
assign a3492 = ~a3400 & a2932;
assign a3494 = a3492 & a3354;
assign a3496 = ~a3492 & ~a3354;
assign a3498 = ~a3496 & ~a3494;
assign a3500 = ~a3476 & ~a3468;
assign a3502 = ~a3500 & ~a3470;
assign a3504 = ~a3502 & ~a3498;
assign a3506 = a3502 & a3498;
assign a3508 = ~a3506 & ~a3504;
assign a3510 = a3508 & a2916;
assign a3512 = ~a3510 & ~a3490;
assign a3514 = ~a3508 & ~a2916;
assign a3516 = ~a3514 & ~a3512;
assign a3518 = ~a3400 & a2916;
assign a3520 = a3518 & a3380;
assign a3522 = ~a3518 & ~a3380;
assign a3524 = ~a3522 & ~a3520;
assign a3526 = ~a3502 & ~a3494;
assign a3528 = ~a3526 & ~a3496;
assign a3530 = ~a3528 & ~a3524;
assign a3532 = a3528 & a3524;
assign a3534 = ~a3532 & ~a3530;
assign a3536 = a3534 & a3516;
assign a3538 = ~a3536 & a2864;
assign a3540 = a3538 & ~a2876;
assign a3542 = ~a3536 & a2880;
assign a3544 = ~a3542 & ~a3408;
assign a3546 = a3542 & a3408;
assign a3548 = ~a3546 & ~a3544;
assign a3550 = ~a3548 & ~a3540;
assign a3552 = a3548 & a3540;
assign a3554 = ~a3552 & ~a3550;
assign a3556 = ~a2866 & i60;
assign a3558 = a2866 & ~i60;
assign a3560 = ~a3558 & ~a3556;
assign a3562 = ~a3560 & ~a2798;
assign a3564 = ~a3562 & a2864;
assign a3566 = ~a3538 & a2876;
assign a3568 = ~a3566 & ~a3540;
assign a3570 = a3568 & a2880;
assign a3572 = ~a3570 & ~a3564;
assign a3574 = ~a3568 & ~a2880;
assign a3576 = ~a3574 & ~a3572;
assign a3578 = a3554 & a2964;
assign a3580 = ~a3578 & ~a3576;
assign a3582 = ~a3554 & ~a2964;
assign a3584 = ~a3582 & ~a3580;
assign a3586 = ~a3546 & ~a3540;
assign a3588 = ~a3586 & ~a3544;
assign a3590 = ~a3536 & a2964;
assign a3592 = ~a3590 & ~a3430;
assign a3594 = a3590 & a3430;
assign a3596 = ~a3594 & ~a3592;
assign a3598 = ~a3596 & ~a3588;
assign a3600 = a3596 & a3588;
assign a3602 = ~a3600 & ~a3598;
assign a3604 = a3602 & a2948;
assign a3606 = ~a3604 & ~a3584;
assign a3608 = ~a3602 & ~a2948;
assign a3610 = ~a3608 & ~a3606;
assign a3612 = ~a3594 & ~a3588;
assign a3614 = ~a3612 & ~a3592;
assign a3616 = ~a3536 & a2948;
assign a3618 = ~a3616 & ~a3456;
assign a3620 = a3616 & a3456;
assign a3622 = ~a3620 & ~a3618;
assign a3624 = ~a3622 & ~a3614;
assign a3626 = a3622 & a3614;
assign a3628 = ~a3626 & ~a3624;
assign a3630 = a3628 & a2932;
assign a3632 = ~a3630 & ~a3610;
assign a3634 = ~a3628 & ~a2932;
assign a3636 = ~a3634 & ~a3632;
assign a3638 = ~a3536 & a2932;
assign a3640 = a3638 & a3482;
assign a3642 = ~a3638 & ~a3482;
assign a3644 = ~a3642 & ~a3640;
assign a3646 = ~a3620 & ~a3614;
assign a3648 = ~a3646 & ~a3618;
assign a3650 = ~a3648 & ~a3644;
assign a3652 = a3648 & a3644;
assign a3654 = ~a3652 & ~a3650;
assign a3656 = a3654 & a2916;
assign a3658 = ~a3656 & ~a3636;
assign a3660 = ~a3654 & ~a2916;
assign a3662 = ~a3660 & ~a3658;
assign a3664 = ~a3536 & a2916;
assign a3666 = a3664 & a3508;
assign a3668 = ~a3664 & ~a3508;
assign a3670 = ~a3668 & ~a3666;
assign a3672 = ~a3648 & ~a3640;
assign a3674 = ~a3672 & ~a3642;
assign a3676 = ~a3674 & ~a3670;
assign a3678 = a3674 & a3670;
assign a3680 = ~a3678 & ~a3676;
assign a3682 = a3680 & a3662;
assign a3684 = ~a3682 & a2964;
assign a3686 = ~a3684 & ~a3554;
assign a3688 = a3684 & a3554;
assign a3690 = ~a3682 & a2880;
assign a3692 = ~a3690 & ~a3568;
assign a3694 = ~a3682 & a2864;
assign a3696 = a3694 & ~a3562;
assign a3698 = a3690 & a3568;
assign a3700 = ~a3698 & ~a3696;
assign a3702 = ~a3700 & ~a3692;
assign a3704 = ~a3702 & ~a3688;
assign a3706 = ~a3704 & ~a3686;
assign a3708 = ~a3682 & a2948;
assign a3710 = ~a3708 & ~a3602;
assign a3712 = a3708 & a3602;
assign a3714 = ~a3712 & ~a3710;
assign a3716 = ~a3714 & ~a3706;
assign a3718 = a3714 & a3706;
assign a3720 = ~a3718 & ~a3716;
assign a3722 = ~a3682 & a2916;
assign a3724 = a3722 & a3654;
assign a3726 = ~a3722 & ~a3654;
assign a3728 = ~a3726 & ~a3724;
assign a3730 = ~a3682 & a2932;
assign a3732 = ~a3730 & ~a3628;
assign a3734 = a3730 & a3628;
assign a3736 = ~a3712 & ~a3706;
assign a3738 = ~a3736 & ~a3710;
assign a3740 = ~a3738 & ~a3734;
assign a3742 = ~a3740 & ~a3732;
assign a3744 = ~a3742 & ~a3728;
assign a3746 = a3742 & a3728;
assign a3748 = ~a3746 & ~a3744;
assign a3750 = i62 & ~i38;
assign a3752 = ~i62 & i38;
assign a3754 = ~a3752 & ~a3750;
assign a3756 = ~a3754 & ~a2798;
assign a3758 = ~a3756 & a2864;
assign a3760 = ~a3694 & a3562;
assign a3762 = ~a3760 & ~a3696;
assign a3764 = a3762 & a2880;
assign a3766 = ~a3764 & ~a3758;
assign a3768 = ~a3762 & ~a2880;
assign a3770 = ~a3768 & ~a3766;
assign a3772 = ~a3698 & ~a3692;
assign a3774 = ~a3772 & ~a3696;
assign a3776 = a3772 & a3696;
assign a3778 = ~a3776 & ~a3774;
assign a3780 = a3778 & a2964;
assign a3782 = ~a3780 & ~a3770;
assign a3784 = ~a3778 & ~a2964;
assign a3786 = ~a3784 & ~a3782;
assign a3788 = ~a3688 & ~a3686;
assign a3790 = ~a3788 & ~a3702;
assign a3792 = a3788 & a3702;
assign a3794 = ~a3792 & ~a3790;
assign a3796 = a3794 & a2948;
assign a3798 = ~a3796 & ~a3786;
assign a3800 = ~a3794 & ~a2948;
assign a3802 = ~a3800 & ~a3798;
assign a3804 = a3720 & a2932;
assign a3806 = ~a3804 & ~a3802;
assign a3808 = ~a3720 & ~a2932;
assign a3810 = ~a3808 & ~a3806;
assign a3812 = ~a3734 & ~a3732;
assign a3814 = ~a3812 & ~a3738;
assign a3816 = a3812 & a3738;
assign a3818 = ~a3816 & ~a3814;
assign a3820 = a3818 & a2916;
assign a3822 = ~a3820 & ~a3810;
assign a3824 = ~a3818 & ~a2916;
assign a3826 = ~a3824 & ~a3822;
assign a3828 = a3826 & a3748;
assign a3830 = ~a3828 & a2932;
assign a3832 = ~a3830 & ~a3720;
assign a3834 = a3830 & a3720;
assign a3836 = ~a3828 & a2948;
assign a3838 = ~a3836 & ~a3794;
assign a3840 = a3836 & a3794;
assign a3842 = ~a3828 & a2964;
assign a3844 = ~a3842 & ~a3778;
assign a3846 = a3842 & a3778;
assign a3848 = ~a3828 & a2880;
assign a3850 = ~a3848 & ~a3762;
assign a3852 = a3848 & a3762;
assign a3854 = ~a3828 & a2864;
assign a3856 = a3854 & ~a3756;
assign a3858 = ~a3856 & ~a3852;
assign a3860 = ~a3858 & ~a3850;
assign a3862 = ~a3860 & ~a3846;
assign a3864 = ~a3862 & ~a3844;
assign a3866 = ~a3864 & ~a3840;
assign a3868 = ~a3866 & ~a3838;
assign a3870 = ~a3868 & ~a3834;
assign a3872 = ~a3870 & ~a3832;
assign a3874 = ~a3828 & a2916;
assign a3876 = ~a3874 & ~a3818;
assign a3878 = a3874 & a3818;
assign a3880 = ~a3878 & ~a3876;
assign a3882 = ~a3880 & ~a3872;
assign a3884 = a3880 & a3872;
assign a3886 = ~a3884 & ~a3882;
assign a3888 = a2864 & ~a2800;
assign a3890 = ~a3854 & a3756;
assign a3892 = ~a3890 & ~a3856;
assign a3894 = a3892 & a2880;
assign a3896 = ~a3894 & ~a3888;
assign a3898 = ~a3892 & ~a2880;
assign a3900 = ~a3898 & ~a3896;
assign a3902 = ~a3852 & ~a3850;
assign a3904 = ~a3902 & ~a3856;
assign a3906 = a3902 & a3856;
assign a3908 = ~a3906 & ~a3904;
assign a3910 = a3908 & a2964;
assign a3912 = ~a3910 & ~a3900;
assign a3914 = ~a3908 & ~a2964;
assign a3916 = ~a3914 & ~a3912;
assign a3918 = ~a3846 & ~a3844;
assign a3920 = ~a3918 & ~a3860;
assign a3922 = a3918 & a3860;
assign a3924 = ~a3922 & ~a3920;
assign a3926 = a3924 & a2948;
assign a3928 = ~a3926 & ~a3916;
assign a3930 = ~a3924 & ~a2948;
assign a3932 = ~a3930 & ~a3928;
assign a3934 = ~a3840 & ~a3838;
assign a3936 = ~a3934 & ~a3864;
assign a3938 = a3934 & a3864;
assign a3940 = ~a3938 & ~a3936;
assign a3942 = a3940 & a2932;
assign a3944 = ~a3942 & ~a3932;
assign a3946 = ~a3940 & ~a2932;
assign a3948 = ~a3946 & ~a3944;
assign a3950 = ~a3834 & ~a3832;
assign a3952 = ~a3950 & ~a3868;
assign a3954 = a3950 & a3868;
assign a3956 = ~a3954 & ~a3952;
assign a3958 = a3956 & a2916;
assign a3960 = ~a3958 & ~a3948;
assign a3962 = ~a3956 & ~a2916;
assign a3964 = ~a3962 & ~a3960;
assign a3966 = a3964 & a3886;
assign a3968 = ~a3966 & a2864;
assign a3970 = a3968 & ~a2800;
assign a3972 = ~a3968 & a2800;
assign a3974 = ~a3972 & ~a3970;
assign a3976 = a3974 & a2560;
assign a3978 = i72 & i70;
assign a3980 = a3978 & i68;
assign a3982 = a3980 & i66;
assign a3984 = a3982 & ~i74;
assign a3986 = ~a3984 & i64;
assign a3988 = a2622 & ~a2550;
assign a3990 = a3988 & a2862;
assign a3992 = a2700 & i78;
assign a3994 = ~a3992 & a2682;
assign a3996 = ~a3994 & a2622;
assign a3998 = a3994 & ~a2622;
assign a4000 = ~a3998 & ~a3996;
assign a4002 = ~a4000 & ~a2550;
assign a4004 = a4002 & i42;
assign a4006 = ~a4004 & ~a3990;
assign a4008 = ~a4002 & ~i42;
assign a4010 = ~a4008 & ~a4006;
assign a4012 = ~a3994 & ~a2622;
assign a4014 = ~a4012 & i18;
assign a4016 = a4012 & ~i18;
assign a4018 = ~a4016 & ~a4014;
assign a4020 = ~a4018 & ~a2550;
assign a4022 = a4020 & i44;
assign a4024 = ~a4022 & ~a4010;
assign a4026 = ~a4020 & ~i44;
assign a4028 = ~a4026 & ~a4024;
assign a4030 = a4012 & i18;
assign a4032 = ~a4030 & i80;
assign a4034 = a4030 & ~i80;
assign a4036 = ~a4034 & ~a4032;
assign a4038 = ~a4036 & ~a2550;
assign a4040 = a4038 & i46;
assign a4042 = ~a4040 & ~a4028;
assign a4044 = ~a4038 & ~i46;
assign a4046 = ~a4044 & ~a4042;
assign a4048 = a4030 & i80;
assign a4050 = ~a4048 & i82;
assign a4052 = a4048 & ~i82;
assign a4054 = ~a4052 & ~a4050;
assign a4056 = ~a4054 & ~a2550;
assign a4058 = a4056 & i48;
assign a4060 = ~a4058 & ~a4046;
assign a4062 = ~a4056 & ~i48;
assign a4064 = ~a4062 & ~a4060;
assign a4066 = a4048 & i82;
assign a4068 = a4066 & ~a2550;
assign a4070 = a4068 & i50;
assign a4072 = ~a4070 & ~a4064;
assign a4074 = ~a4068 & ~i50;
assign a4076 = ~a4074 & ~a4072;
assign a4078 = ~a4076 & ~a2700;
assign a4080 = a4078 & i76;
assign a4082 = ~a2674 & ~a2668;
assign a4084 = a4082 & ~a2624;
assign a4086 = ~a2558 & i14;
assign a4088 = a3988 & ~i84;
assign a4090 = ~a3988 & i84;
assign a4092 = ~a4090 & ~a4088;
assign a4094 = a4092 & i12;
assign a4096 = a3988 & ~i12;
assign a4098 = ~a4096 & ~a4094;
assign a4100 = ~a4098 & i14;
assign a4102 = i86 & ~i14;
assign a4104 = ~a4102 & ~a4100;
assign a4106 = ~a4104 & a4086;
assign a4108 = ~a4106 & a4084;
assign a4110 = ~a4108 & a4080;
assign a4112 = a4110 & a3986;
assign a4114 = ~a4110 & ~a3986;
assign a4116 = ~a4114 & ~a4112;
assign a4118 = ~a4116 & a2706;
assign a4120 = a4076 & i88;
assign a4122 = a4120 & ~i90;
assign a4124 = a3986 & ~a2862;
assign a4126 = ~a3986 & a2862;
assign a4128 = ~a4126 & ~a4124;
assign a4130 = ~a4128 & a4122;
assign a4132 = ~a4122 & ~a2862;
assign a4134 = ~a4132 & ~a4130;
assign a4136 = ~a4134 & ~a2706;
assign a4138 = ~a4136 & ~a4118;
assign a4140 = a2722 & i92;
assign a4142 = ~a4140 & a2730;
assign a4144 = ~a4142 & a2712;
assign a4146 = ~a4144 & ~a2764;
assign a4148 = a4146 & ~a2736;
assign a4150 = a4148 & ~a4122;
assign a4152 = a4150 & ~a2712;
assign a4154 = a4152 & ~a4138;
assign a4156 = a4122 & a2862;
assign a4158 = ~a4122 & i94;
assign a4160 = ~a4158 & ~a4156;
assign a4162 = a4160 & a4122;
assign a4164 = ~a4162 & ~a4110;
assign a4166 = a4164 & ~a4154;
assign a4168 = ~a4098 & ~i96;
assign a4170 = a4098 & i96;
assign a4172 = ~a4170 & ~a4168;
assign a4174 = a4172 & i14;
assign a4176 = ~a4098 & ~i14;
assign a4178 = ~a4176 & ~a4174;
assign a4180 = ~a4178 & a2700;
assign a4182 = ~a4180 & a4084;
assign a4184 = ~a4182 & a4166;
assign a4186 = a4110 & ~a3986;
assign a4188 = a3988 & i84;
assign a4190 = a4002 & ~i98;
assign a4192 = ~a4002 & i98;
assign a4194 = ~a4192 & ~a4190;
assign a4196 = ~a4194 & ~a4188;
assign a4198 = a4194 & a4188;
assign a4200 = ~a4198 & ~a4196;
assign a4202 = ~a4200 & a4092;
assign a4204 = a4200 & ~a4092;
assign a4206 = ~a4204 & ~a4202;
assign a4208 = ~a4206 & i12;
assign a4210 = a4002 & ~i12;
assign a4212 = ~a4210 & ~a4208;
assign a4214 = ~a4212 & i14;
assign a4216 = i100 & ~i14;
assign a4218 = ~a4216 & ~a4214;
assign a4220 = ~a4218 & a4086;
assign a4222 = a4002 & i12;
assign a4224 = ~a4222 & ~a4220;
assign a4226 = ~a4224 & a4080;
assign a4228 = a4226 & i66;
assign a4230 = ~a4226 & ~i66;
assign a4232 = ~a4230 & ~a4228;
assign a4234 = ~a4232 & ~a4186;
assign a4236 = a4232 & a4186;
assign a4238 = ~a4236 & ~a4234;
assign a4240 = ~a4238 & a2706;
assign a4242 = ~a3986 & ~a2862;
assign a4244 = i66 & ~i42;
assign a4246 = ~i66 & i42;
assign a4248 = ~a4246 & ~a4244;
assign a4250 = ~a4248 & ~a4242;
assign a4252 = a4248 & a4242;
assign a4254 = ~a4252 & ~a4250;
assign a4256 = ~a4254 & a4122;
assign a4258 = ~a4122 & ~i42;
assign a4260 = ~a4258 & ~a4256;
assign a4262 = ~a4260 & ~a2706;
assign a4264 = ~a4262 & ~a4240;
assign a4266 = ~a4264 & a4152;
assign a4268 = a4122 & i42;
assign a4270 = ~a4122 & i102;
assign a4272 = ~a4270 & ~a4268;
assign a4274 = a4272 & a4122;
assign a4276 = ~a4274 & ~a4226;
assign a4278 = a4276 & ~a4266;
assign a4280 = ~a4098 & i96;
assign a4282 = ~a4212 & ~i104;
assign a4284 = a4212 & i104;
assign a4286 = ~a4284 & ~a4282;
assign a4288 = ~a4286 & ~a4280;
assign a4290 = a4286 & a4280;
assign a4292 = ~a4290 & ~a4288;
assign a4294 = ~a4292 & a4172;
assign a4296 = a4292 & ~a4172;
assign a4298 = ~a4296 & ~a4294;
assign a4300 = ~a4298 & i14;
assign a4302 = ~a4212 & ~i14;
assign a4304 = ~a4302 & ~a4300;
assign a4306 = ~a4304 & a2700;
assign a4308 = ~a4306 & ~a4222;
assign a4310 = ~a4308 & a4278;
assign a4312 = ~a4310 & ~a4184;
assign a4314 = a4308 & ~a4278;
assign a4316 = ~a4314 & ~a4312;
assign a4318 = a4226 & ~i66;
assign a4320 = ~a4318 & ~a4186;
assign a4322 = ~a4226 & i66;
assign a4324 = ~a4322 & ~a4320;
assign a4326 = ~a4200 & ~a4092;
assign a4328 = a4002 & i98;
assign a4330 = ~a4328 & ~a4188;
assign a4332 = ~a4002 & ~i98;
assign a4334 = ~a4332 & ~a4330;
assign a4336 = a4020 & ~i106;
assign a4338 = ~a4020 & i106;
assign a4340 = ~a4338 & ~a4336;
assign a4342 = ~a4340 & ~a4334;
assign a4344 = a4340 & a4334;
assign a4346 = ~a4344 & ~a4342;
assign a4348 = ~a4346 & ~a4326;
assign a4350 = a4346 & a4326;
assign a4352 = ~a4350 & ~a4348;
assign a4354 = ~a4352 & i12;
assign a4356 = a4020 & ~i12;
assign a4358 = ~a4356 & ~a4354;
assign a4360 = ~a4358 & i14;
assign a4362 = i108 & ~i14;
assign a4364 = ~a4362 & ~a4360;
assign a4366 = ~a4364 & a4086;
assign a4368 = a4020 & i12;
assign a4370 = ~a4368 & ~a4366;
assign a4372 = ~a4370 & a4080;
assign a4374 = a4372 & i68;
assign a4376 = ~a4372 & ~i68;
assign a4378 = ~a4376 & ~a4374;
assign a4380 = ~a4378 & ~a4324;
assign a4382 = a4378 & a4324;
assign a4384 = ~a4382 & ~a4380;
assign a4386 = ~a4384 & a2706;
assign a4388 = ~i66 & ~i42;
assign a4390 = ~a4388 & ~a4242;
assign a4392 = i66 & i42;
assign a4394 = ~a4392 & ~a4390;
assign a4396 = i68 & ~i44;
assign a4398 = ~i68 & i44;
assign a4400 = ~a4398 & ~a4396;
assign a4402 = ~a4400 & ~a4394;
assign a4404 = a4400 & a4394;
assign a4406 = ~a4404 & ~a4402;
assign a4408 = ~a4406 & a4122;
assign a4410 = ~a4122 & ~i44;
assign a4412 = ~a4410 & ~a4408;
assign a4414 = ~a4412 & ~a2706;
assign a4416 = ~a4414 & ~a4386;
assign a4418 = ~a4416 & a4152;
assign a4420 = a4122 & i44;
assign a4422 = ~a4122 & i110;
assign a4424 = ~a4422 & ~a4420;
assign a4426 = a4424 & a4122;
assign a4428 = ~a4426 & ~a4372;
assign a4430 = a4428 & ~a4418;
assign a4432 = ~a4292 & ~a4172;
assign a4434 = ~a4212 & i104;
assign a4436 = ~a4434 & ~a4280;
assign a4438 = a4212 & ~i104;
assign a4440 = ~a4438 & ~a4436;
assign a4442 = ~a4358 & ~i112;
assign a4444 = a4358 & i112;
assign a4446 = ~a4444 & ~a4442;
assign a4448 = ~a4446 & ~a4440;
assign a4450 = a4446 & a4440;
assign a4452 = ~a4450 & ~a4448;
assign a4454 = ~a4452 & ~a4432;
assign a4456 = a4452 & a4432;
assign a4458 = ~a4456 & ~a4454;
assign a4460 = ~a4458 & i14;
assign a4462 = ~a4358 & ~i14;
assign a4464 = ~a4462 & ~a4460;
assign a4466 = ~a4464 & a2700;
assign a4468 = ~a4466 & ~a4368;
assign a4470 = ~a4468 & a4430;
assign a4472 = ~a4470 & ~a4316;
assign a4474 = a4468 & ~a4430;
assign a4476 = ~a4474 & ~a4472;
assign a4478 = a4372 & ~i68;
assign a4480 = ~a4478 & ~a4324;
assign a4482 = ~a4372 & i68;
assign a4484 = ~a4482 & ~a4480;
assign a4486 = ~a4346 & a4326;
assign a4488 = a4020 & i106;
assign a4490 = ~a4488 & ~a4334;
assign a4492 = ~a4020 & ~i106;
assign a4494 = ~a4492 & ~a4490;
assign a4496 = a4038 & ~i114;
assign a4498 = ~a4038 & i114;
assign a4500 = ~a4498 & ~a4496;
assign a4502 = ~a4500 & ~a4494;
assign a4504 = a4500 & a4494;
assign a4506 = ~a4504 & ~a4502;
assign a4508 = ~a4506 & ~a4486;
assign a4510 = a4506 & a4486;
assign a4512 = ~a4510 & ~a4508;
assign a4514 = ~a4512 & i12;
assign a4516 = a4038 & ~i12;
assign a4518 = ~a4516 & ~a4514;
assign a4520 = ~a4518 & i14;
assign a4522 = i116 & ~i14;
assign a4524 = ~a4522 & ~a4520;
assign a4526 = ~a4524 & a4086;
assign a4528 = a4038 & i12;
assign a4530 = ~a4528 & ~a4526;
assign a4532 = ~a4530 & a4080;
assign a4534 = a4532 & i72;
assign a4536 = ~a4532 & ~i72;
assign a4538 = ~a4536 & ~a4534;
assign a4540 = ~a4538 & ~a4484;
assign a4542 = a4538 & a4484;
assign a4544 = ~a4542 & ~a4540;
assign a4546 = ~a4544 & a2706;
assign a4548 = ~i68 & ~i44;
assign a4550 = ~a4548 & ~a4394;
assign a4552 = i68 & i44;
assign a4554 = ~a4552 & ~a4550;
assign a4556 = i72 & ~i46;
assign a4558 = ~i72 & i46;
assign a4560 = ~a4558 & ~a4556;
assign a4562 = ~a4560 & ~a4554;
assign a4564 = a4560 & a4554;
assign a4566 = ~a4564 & ~a4562;
assign a4568 = ~a4566 & a4122;
assign a4570 = ~a4122 & ~i46;
assign a4572 = ~a4570 & ~a4568;
assign a4574 = ~a4572 & ~a2706;
assign a4576 = ~a4574 & ~a4546;
assign a4578 = ~a4576 & a4152;
assign a4580 = a4122 & i46;
assign a4582 = ~a4122 & i118;
assign a4584 = ~a4582 & ~a4580;
assign a4586 = a4584 & a4122;
assign a4588 = ~a4586 & ~a4532;
assign a4590 = a4588 & ~a4578;
assign a4592 = ~a4452 & a4432;
assign a4594 = ~a4358 & i112;
assign a4596 = ~a4594 & ~a4440;
assign a4598 = a4358 & ~i112;
assign a4600 = ~a4598 & ~a4596;
assign a4602 = ~a4518 & ~i120;
assign a4604 = a4518 & i120;
assign a4606 = ~a4604 & ~a4602;
assign a4608 = ~a4606 & ~a4600;
assign a4610 = a4606 & a4600;
assign a4612 = ~a4610 & ~a4608;
assign a4614 = ~a4612 & ~a4592;
assign a4616 = a4612 & a4592;
assign a4618 = ~a4616 & ~a4614;
assign a4620 = ~a4618 & i14;
assign a4622 = ~a4518 & ~i14;
assign a4624 = ~a4622 & ~a4620;
assign a4626 = ~a4624 & a2700;
assign a4628 = ~a4626 & ~a4528;
assign a4630 = ~a4628 & a4590;
assign a4632 = ~a4630 & ~a4476;
assign a4634 = a4628 & ~a4590;
assign a4636 = ~a4634 & ~a4632;
assign a4638 = a4532 & ~i72;
assign a4640 = ~a4638 & ~a4484;
assign a4642 = ~a4532 & i72;
assign a4644 = ~a4642 & ~a4640;
assign a4646 = ~a4506 & a4486;
assign a4648 = a4038 & i114;
assign a4650 = ~a4648 & ~a4494;
assign a4652 = ~a4038 & ~i114;
assign a4654 = ~a4652 & ~a4650;
assign a4656 = a4056 & ~i122;
assign a4658 = ~a4056 & i122;
assign a4660 = ~a4658 & ~a4656;
assign a4662 = ~a4660 & ~a4654;
assign a4664 = a4660 & a4654;
assign a4666 = ~a4664 & ~a4662;
assign a4668 = ~a4666 & ~a4646;
assign a4670 = a4666 & a4646;
assign a4672 = ~a4670 & ~a4668;
assign a4674 = ~a4672 & i12;
assign a4676 = a4056 & ~i12;
assign a4678 = ~a4676 & ~a4674;
assign a4680 = ~a4678 & i14;
assign a4682 = i124 & ~i14;
assign a4684 = ~a4682 & ~a4680;
assign a4686 = ~a4684 & a4086;
assign a4688 = a4056 & i12;
assign a4690 = ~a4688 & ~a4686;
assign a4692 = ~a4690 & a4080;
assign a4694 = a4692 & i70;
assign a4696 = ~a4692 & ~i70;
assign a4698 = ~a4696 & ~a4694;
assign a4700 = ~a4698 & ~a4644;
assign a4702 = a4698 & a4644;
assign a4704 = ~a4702 & ~a4700;
assign a4706 = ~a4704 & a2706;
assign a4708 = ~i72 & ~i46;
assign a4710 = ~a4708 & ~a4554;
assign a4712 = i72 & i46;
assign a4714 = ~a4712 & ~a4710;
assign a4716 = i70 & ~i48;
assign a4718 = ~i70 & i48;
assign a4720 = ~a4718 & ~a4716;
assign a4722 = ~a4720 & ~a4714;
assign a4724 = a4720 & a4714;
assign a4726 = ~a4724 & ~a4722;
assign a4728 = ~a4726 & a4122;
assign a4730 = ~a4122 & ~i48;
assign a4732 = ~a4730 & ~a4728;
assign a4734 = ~a4732 & ~a2706;
assign a4736 = ~a4734 & ~a4706;
assign a4738 = ~a4736 & a4152;
assign a4740 = a4122 & i48;
assign a4742 = ~a4122 & i126;
assign a4744 = ~a4742 & ~a4740;
assign a4746 = a4744 & a4122;
assign a4748 = ~a4746 & ~a4692;
assign a4750 = a4748 & ~a4738;
assign a4752 = ~a4612 & a4592;
assign a4754 = ~a4518 & i120;
assign a4756 = ~a4754 & ~a4600;
assign a4758 = a4518 & ~i120;
assign a4760 = ~a4758 & ~a4756;
assign a4762 = ~a4678 & ~i128;
assign a4764 = a4678 & i128;
assign a4766 = ~a4764 & ~a4762;
assign a4768 = ~a4766 & ~a4760;
assign a4770 = a4766 & a4760;
assign a4772 = ~a4770 & ~a4768;
assign a4774 = ~a4772 & ~a4752;
assign a4776 = a4772 & a4752;
assign a4778 = ~a4776 & ~a4774;
assign a4780 = ~a4778 & i14;
assign a4782 = ~a4678 & ~i14;
assign a4784 = ~a4782 & ~a4780;
assign a4786 = ~a4784 & a2700;
assign a4788 = ~a4786 & ~a4688;
assign a4790 = ~a4788 & a4750;
assign a4792 = ~a4790 & ~a4636;
assign a4794 = a4788 & ~a4750;
assign a4796 = ~a4794 & ~a4792;
assign a4798 = ~a4666 & a4646;
assign a4800 = a4056 & i122;
assign a4802 = ~a4800 & ~a4654;
assign a4804 = ~a4056 & ~i122;
assign a4806 = ~a4804 & ~a4802;
assign a4808 = ~a4806 & ~a4068;
assign a4810 = ~a4808 & ~a4798;
assign a4812 = a4808 & a4798;
assign a4814 = ~a4812 & ~a4810;
assign a4816 = ~a4814 & i12;
assign a4818 = a4068 & ~i12;
assign a4820 = ~a4818 & ~a4816;
assign a4822 = ~a4820 & i14;
assign a4824 = i130 & ~i14;
assign a4826 = ~a4824 & ~a4822;
assign a4828 = ~a4826 & a4086;
assign a4830 = a4068 & i12;
assign a4832 = ~a4830 & ~a4828;
assign a4834 = ~a4832 & a4080;
assign a4836 = a4692 & ~i70;
assign a4838 = ~a4836 & ~a4644;
assign a4840 = ~a4692 & i70;
assign a4842 = ~a4840 & ~a4838;
assign a4844 = a4834 & ~i74;
assign a4846 = ~a4834 & i74;
assign a4848 = ~a4846 & ~a4844;
assign a4850 = ~a4848 & ~a4842;
assign a4852 = a4848 & a4842;
assign a4854 = ~a4852 & ~a4850;
assign a4856 = ~a4854 & a2706;
assign a4858 = ~i70 & ~i48;
assign a4860 = ~a4858 & ~a4714;
assign a4862 = i70 & i48;
assign a4864 = ~a4862 & ~a4860;
assign a4866 = ~i74 & ~i50;
assign a4868 = i74 & i50;
assign a4870 = ~a4868 & ~a4866;
assign a4872 = ~a4870 & ~a4864;
assign a4874 = a4870 & a4864;
assign a4876 = ~a4874 & ~a4872;
assign a4878 = ~a4876 & a4122;
assign a4880 = ~a4878 & i50;
assign a4882 = ~a4880 & ~a2706;
assign a4884 = ~a4882 & ~a4856;
assign a4886 = ~a4884 & a4152;
assign a4888 = ~a4886 & ~a4834;
assign a4890 = ~a4772 & a4752;
assign a4892 = ~a4678 & i128;
assign a4894 = ~a4892 & ~a4760;
assign a4896 = a4678 & ~i128;
assign a4898 = ~a4896 & ~a4894;
assign a4900 = ~a4898 & ~a4820;
assign a4902 = a4898 & a4820;
assign a4904 = ~a4902 & ~a4900;
assign a4906 = ~a4904 & ~a4890;
assign a4908 = a4904 & a4890;
assign a4910 = ~a4908 & ~a4906;
assign a4912 = ~a4910 & i14;
assign a4914 = ~a4820 & ~i14;
assign a4916 = ~a4914 & ~a4912;
assign a4918 = ~a4916 & a2700;
assign a4920 = ~a4918 & ~a4830;
assign a4922 = ~a4920 & a4888;
assign a4924 = ~a4922 & ~a4796;
assign a4926 = a4920 & ~a4888;
assign a4928 = ~a4926 & ~a4924;
assign a4930 = ~a4904 & a4890;
assign a4932 = ~a4808 & a4798;
assign a4934 = a4932 & i12;
assign a4936 = a4898 & ~a4820;
assign a4938 = ~a4936 & ~a4934;
assign a4940 = a4938 & ~a4930;
assign a4942 = ~a4940 & i14;
assign a4944 = a4934 & ~i14;
assign a4946 = ~a4944 & ~a4942;
assign a4948 = ~a4946 & a2700;
assign a4950 = ~a4948 & ~a4928;
assign a4952 = ~a4950 & ~a4166;
assign a4954 = ~a4952 & a3976;
assign a4956 = a4950 & a4182;
assign a4958 = ~a4956 & a4954;
assign a4960 = ~a3966 & a2880;
assign a4962 = ~a4960 & ~a3892;
assign a4964 = a4960 & a3892;
assign a4966 = ~a4964 & ~a4962;
assign a4968 = ~a4966 & ~a3970;
assign a4970 = a4966 & a3970;
assign a4972 = ~a4970 & ~a4968;
assign a4974 = ~a4972 & a3974;
assign a4976 = a4972 & ~a3974;
assign a4978 = ~a4976 & ~a4974;
assign a4980 = ~a4978 & a2560;
assign a4982 = ~a4950 & ~a4278;
assign a4984 = a4308 & a4182;
assign a4986 = ~a4308 & ~a4182;
assign a4988 = ~a4986 & ~a4984;
assign a4990 = ~a4988 & a4950;
assign a4992 = ~a4990 & ~a4982;
assign a4994 = a4992 & a4980;
assign a4996 = ~a4994 & ~a4958;
assign a4998 = ~a4992 & ~a4980;
assign a5000 = ~a4998 & ~a4996;
assign a5002 = ~a4972 & ~a3974;
assign a5004 = ~a4964 & ~a3970;
assign a5006 = ~a5004 & ~a4962;
assign a5008 = ~a3966 & a2964;
assign a5010 = ~a5008 & ~a3908;
assign a5012 = a5008 & a3908;
assign a5014 = ~a5012 & ~a5010;
assign a5016 = ~a5014 & ~a5006;
assign a5018 = a5014 & a5006;
assign a5020 = ~a5018 & ~a5016;
assign a5022 = ~a5020 & ~a5002;
assign a5024 = a5020 & a5002;
assign a5026 = ~a5024 & ~a5022;
assign a5028 = ~a5026 & a2560;
assign a5030 = ~a4950 & ~a4430;
assign a5032 = a4984 & a4468;
assign a5034 = ~a4984 & ~a4468;
assign a5036 = ~a5034 & ~a5032;
assign a5038 = ~a5036 & a4950;
assign a5040 = ~a5038 & ~a5030;
assign a5042 = a5040 & a5028;
assign a5044 = ~a5042 & ~a5000;
assign a5046 = ~a5040 & ~a5028;
assign a5048 = ~a5046 & ~a5044;
assign a5050 = ~a5020 & a5002;
assign a5052 = ~a5012 & ~a5006;
assign a5054 = ~a5052 & ~a5010;
assign a5056 = ~a3966 & a2948;
assign a5058 = ~a5056 & ~a3924;
assign a5060 = a5056 & a3924;
assign a5062 = ~a5060 & ~a5058;
assign a5064 = ~a5062 & ~a5054;
assign a5066 = a5062 & a5054;
assign a5068 = ~a5066 & ~a5064;
assign a5070 = ~a5068 & ~a5050;
assign a5072 = a5068 & a5050;
assign a5074 = ~a5072 & ~a5070;
assign a5076 = ~a5074 & a2560;
assign a5078 = ~a4950 & ~a4590;
assign a5080 = a5032 & a4628;
assign a5082 = ~a5032 & ~a4628;
assign a5084 = ~a5082 & ~a5080;
assign a5086 = ~a5084 & a4950;
assign a5088 = ~a5086 & ~a5078;
assign a5090 = a5088 & a5076;
assign a5092 = ~a5090 & ~a5048;
assign a5094 = ~a5088 & ~a5076;
assign a5096 = ~a5094 & ~a5092;
assign a5098 = ~a5068 & a5050;
assign a5100 = ~a5060 & ~a5054;
assign a5102 = ~a5100 & ~a5058;
assign a5104 = ~a3966 & a2932;
assign a5106 = ~a5104 & ~a3940;
assign a5108 = a5104 & a3940;
assign a5110 = ~a5108 & ~a5106;
assign a5112 = ~a5110 & ~a5102;
assign a5114 = a5110 & a5102;
assign a5116 = ~a5114 & ~a5112;
assign a5118 = ~a5116 & ~a5098;
assign a5120 = a5116 & a5098;
assign a5122 = ~a5120 & ~a5118;
assign a5124 = ~a5122 & a2560;
assign a5126 = ~a4950 & ~a4750;
assign a5128 = a5080 & a4788;
assign a5130 = ~a5080 & ~a4788;
assign a5132 = ~a5130 & ~a5128;
assign a5134 = ~a5132 & a4950;
assign a5136 = ~a5134 & ~a5126;
assign a5138 = a5136 & a5124;
assign a5140 = ~a5138 & ~a5096;
assign a5142 = ~a5136 & ~a5124;
assign a5144 = ~a5142 & ~a5140;
assign a5146 = ~a5116 & a5098;
assign a5148 = ~a5108 & ~a5102;
assign a5150 = ~a5148 & ~a5106;
assign a5152 = ~a3966 & a2916;
assign a5154 = ~a5152 & ~a3956;
assign a5156 = a5152 & a3956;
assign a5158 = ~a5156 & ~a5154;
assign a5160 = ~a5158 & ~a5150;
assign a5162 = a5158 & a5150;
assign a5164 = ~a5162 & ~a5160;
assign a5166 = ~a5164 & ~a5146;
assign a5168 = a5164 & a5146;
assign a5170 = ~a5168 & ~a5166;
assign a5172 = ~a5170 & a2560;
assign a5174 = ~a5172 & ~a5144;
assign a5176 = a5174 & ~a2712;
assign a5178 = a5176 & a2786;
assign a5180 = ~a5178 & a2784;
assign a5182 = i132 & i2;
assign a5184 = ~i136 & ~i134;
assign a5186 = a5184 & ~i138;
assign a5188 = a5186 & ~i140;
assign a5190 = a5188 & ~i142;
assign a5192 = a5190 & ~i144;
assign a5194 = a5192 & ~i146;
assign a5196 = ~a5194 & ~i148;
assign a5198 = ~a4178 & a2710;
assign a5200 = ~a5198 & a4108;
assign a5202 = a5200 & a3976;
assign a5204 = ~a4304 & a2710;
assign a5206 = ~a5204 & a4224;
assign a5208 = a5206 & a4980;
assign a5210 = ~a5208 & ~a5202;
assign a5212 = ~a5206 & ~a4980;
assign a5214 = ~a5212 & ~a5210;
assign a5216 = ~a4464 & a2710;
assign a5218 = ~a5216 & a4370;
assign a5220 = a5218 & a5028;
assign a5222 = ~a5220 & ~a5214;
assign a5224 = ~a5218 & ~a5028;
assign a5226 = ~a5224 & ~a5222;
assign a5228 = ~a4624 & a2710;
assign a5230 = ~a5228 & a4530;
assign a5232 = a5230 & a5076;
assign a5234 = ~a5232 & ~a5226;
assign a5236 = ~a5230 & ~a5076;
assign a5238 = ~a5236 & ~a5234;
assign a5240 = ~a4784 & a2710;
assign a5242 = ~a5240 & a4690;
assign a5244 = a5242 & a5124;
assign a5246 = ~a5244 & ~a5238;
assign a5248 = ~a5242 & ~a5124;
assign a5250 = ~a5248 & ~a5246;
assign a5252 = ~a4916 & a2710;
assign a5254 = ~a5252 & a4832;
assign a5256 = a5254 & a5172;
assign a5258 = ~a5256 & ~a5250;
assign a5260 = ~a5254 & ~a5172;
assign a5262 = ~a5260 & ~a5258;
assign a5264 = ~a5262 & a3976;
assign a5266 = a5262 & ~a5200;
assign a5268 = ~a5266 & ~a5264;
assign a5270 = ~a5268 & ~i134;
assign a5272 = ~a5262 & a4980;
assign a5274 = a5262 & ~a5206;
assign a5276 = ~a5274 & ~a5272;
assign a5278 = ~a5276 & ~i136;
assign a5280 = ~a5278 & ~a5270;
assign a5282 = a5276 & i136;
assign a5284 = ~a5282 & ~a5280;
assign a5286 = ~a5262 & a5028;
assign a5288 = a5262 & ~a5218;
assign a5290 = ~a5288 & ~a5286;
assign a5292 = ~a5290 & ~i138;
assign a5294 = ~a5292 & ~a5284;
assign a5296 = a5290 & i138;
assign a5298 = ~a5296 & ~a5294;
assign a5300 = ~a5262 & a5076;
assign a5302 = a5262 & ~a5230;
assign a5304 = ~a5302 & ~a5300;
assign a5306 = ~a5304 & ~i140;
assign a5308 = ~a5306 & ~a5298;
assign a5310 = a5304 & i140;
assign a5312 = ~a5310 & ~a5308;
assign a5314 = ~a5262 & a5124;
assign a5316 = a5262 & ~a5242;
assign a5318 = ~a5316 & ~a5314;
assign a5320 = ~a5318 & ~i142;
assign a5322 = ~a5320 & ~a5312;
assign a5324 = a5318 & i142;
assign a5326 = ~a5324 & ~a5322;
assign a5328 = ~a5262 & a5172;
assign a5330 = a5262 & ~a5254;
assign a5332 = ~a5330 & ~a5328;
assign a5334 = ~a5332 & ~i144;
assign a5336 = ~a5334 & ~a5326;
assign a5338 = a5332 & i144;
assign a5340 = ~a5338 & ~a5336;
assign a5342 = a5340 & ~i146;
assign a5344 = a5342 & a5196;
assign a5346 = a5344 & a5182;
assign a5348 = ~a5346 & a5180;
assign a5350 = ~a5348 & ~l890;
assign a5354 = ~l920 & l890;
assign a5356 = ~a2706 & ~l890;
assign a5358 = ~a5356 & ~a5354;
assign a5362 = ~l894 & ~l892;
assign a5364 = ~l906 & l890;
assign a5366 = a5178 & a4122;
assign a5368 = a5366 & ~i150;
assign a5370 = a5368 & ~i152;
assign a5372 = ~a5370 & ~l890;
assign a5376 = ~a5374 & ~l896;
assign a5378 = a5376 & ~l1762;
assign a5380 = a5378 & ~l1760;
assign a5382 = a5380 & ~l1196;
assign a5384 = a5382 & ~l1198;
assign a5386 = a5384 & ~l904;
assign a5388 = a5386 & ~l898;
assign a5390 = a5388 & ~l900;
assign a5392 = a5390 & ~l902;
assign a5394 = a5392 & a5362;
assign a5396 = ~l938 & l890;
assign a5398 = ~l890 & ~i180;
assign a5400 = ~a5398 & ~a5396;
assign a5402 = a5400 & ~l908;
assign a5404 = a5402 & ~i252;
assign a5406 = ~a5360 & ~l886;
assign a5408 = a5406 & ~l884;
assign a5410 = ~l918 & l890;
assign a5412 = i160 & ~i2;
assign a5414 = i162 & i2;
assign a5416 = a5414 & a2590;
assign a5418 = ~a5416 & i2;
assign a5420 = a5414 & a2570;
assign a5422 = ~a5420 & a5418;
assign a5424 = a5422 & i164;
assign a5426 = i166 & i2;
assign a5428 = i168 & i2;
assign a5430 = ~a5428 & ~a4108;
assign a5432 = i170 & i2;
assign a5434 = ~a5432 & ~a4224;
assign a5436 = ~a5434 & ~a5430;
assign a5438 = a5432 & a4224;
assign a5440 = ~a5438 & ~a5436;
assign a5442 = i172 & i2;
assign a5444 = ~a5442 & ~a4370;
assign a5446 = ~a5444 & ~a5440;
assign a5448 = a5442 & a4370;
assign a5450 = ~a5448 & ~a5446;
assign a5452 = i174 & i2;
assign a5454 = ~a5452 & ~a4530;
assign a5456 = ~a5454 & ~a5450;
assign a5458 = a5452 & a4530;
assign a5460 = ~a5458 & ~a5456;
assign a5462 = i176 & i2;
assign a5464 = ~a5462 & ~a4690;
assign a5466 = ~a5464 & ~a5460;
assign a5468 = a5462 & a4690;
assign a5470 = ~a5468 & ~a5466;
assign a5472 = i178 & i2;
assign a5474 = ~a5472 & ~a4832;
assign a5476 = ~a5474 & ~a5470;
assign a5478 = a5472 & a4832;
assign a5480 = ~a5478 & ~a5476;
assign a5482 = a5480 & ~a5426;
assign a5484 = a5482 & ~a5424;
assign a5486 = ~a5482 & a5424;
assign a5488 = ~a5486 & ~a5484;
assign a5490 = ~a5488 & ~a4148;
assign a5492 = ~a5428 & ~a4182;
assign a5494 = ~a5432 & ~a4308;
assign a5496 = ~a5494 & ~a5492;
assign a5498 = a5432 & a4308;
assign a5500 = ~a5498 & ~a5496;
assign a5502 = ~a5442 & ~a4468;
assign a5504 = ~a5502 & ~a5500;
assign a5506 = a5442 & a4468;
assign a5508 = ~a5506 & ~a5504;
assign a5510 = ~a5452 & ~a4628;
assign a5512 = ~a5510 & ~a5508;
assign a5514 = a5452 & a4628;
assign a5516 = ~a5514 & ~a5512;
assign a5518 = ~a5462 & ~a4788;
assign a5520 = ~a5518 & ~a5516;
assign a5522 = a5462 & a4788;
assign a5524 = ~a5522 & ~a5520;
assign a5526 = ~a5472 & ~a4920;
assign a5528 = ~a5526 & ~a5524;
assign a5530 = a5472 & a4920;
assign a5532 = ~a5530 & ~a5528;
assign a5534 = ~a5426 & a4948;
assign a5536 = ~a5534 & ~a5532;
assign a5538 = a5426 & ~a4948;
assign a5540 = ~a5538 & ~a5536;
assign a5542 = a5540 & ~a5424;
assign a5544 = ~a5540 & a5424;
assign a5546 = ~a5544 & ~a5542;
assign a5548 = ~a5546 & a4148;
assign a5550 = ~a5548 & ~a5490;
assign a5552 = ~a5550 & a5414;
assign a5554 = ~a5552 & ~a5412;
assign a5556 = ~a5554 & ~a2706;
assign a5558 = ~a5556 & ~i2;
assign a5560 = a5558 & ~l890;
assign a5562 = ~a5560 & ~a5410;
assign a5564 = ~l952 & l890;
assign a5566 = a4142 & ~l890;
assign a5568 = ~a5566 & ~a5564;
assign a5570 = ~l954 & l890;
assign a5572 = ~a2564 & i92;
assign a5574 = i194 & ~i92;
assign a5576 = ~a2710 & i92;
assign a5578 = i196 & ~i92;
assign a5580 = ~a5578 & ~a5576;
assign a5582 = i198 & ~i92;
assign a5584 = ~a5582 & a5580;
assign a5586 = a5584 & ~a5574;
assign a5588 = a5586 & a5572;
assign a5590 = ~a5588 & a2710;
assign a5592 = a5590 & ~l890;
assign a5594 = ~a5592 & ~a5570;
assign a5596 = ~l956 & l890;
assign a5598 = ~a2736 & ~l890;
assign a5600 = ~a5598 & ~a5596;
assign a5602 = ~l958 & l890;
assign a5604 = ~a4140 & ~l890;
assign a5606 = ~a5604 & ~a5602;
assign a5608 = ~l970 & ~l968;
assign a5610 = a5608 & ~l966;
assign a5612 = a5610 & ~l964;
assign a5614 = a5612 & ~l962;
assign a5616 = a5614 & ~l960;
assign a5618 = a5616 & ~a5606;
assign a5620 = a5618 & ~a5600;
assign a5622 = a5620 & ~a5594;
assign a5626 = ~a2512 & l886;
assign a5628 = l928 & l898;
assign a5630 = ~l950 & l890;
assign a5632 = ~a4178 & i226;
assign a5634 = ~a4304 & ~i228;
assign a5636 = a4304 & i228;
assign a5638 = ~a5636 & ~a5634;
assign a5640 = ~a5638 & ~a5632;
assign a5642 = a5638 & a5632;
assign a5644 = ~a5642 & ~a5640;
assign a5646 = ~a4178 & ~i226;
assign a5648 = a4178 & i226;
assign a5650 = ~a5648 & ~a5646;
assign a5652 = ~a5650 & ~a5644;
assign a5654 = ~a4304 & i228;
assign a5656 = ~a5654 & ~a5632;
assign a5658 = a4304 & ~i228;
assign a5660 = ~a5658 & ~a5656;
assign a5662 = ~a4464 & ~i230;
assign a5664 = a4464 & i230;
assign a5666 = ~a5664 & ~a5662;
assign a5668 = ~a5666 & ~a5660;
assign a5670 = a5666 & a5660;
assign a5672 = ~a5670 & ~a5668;
assign a5674 = ~a5672 & a5652;
assign a5676 = ~a4464 & i230;
assign a5678 = ~a5676 & ~a5660;
assign a5680 = a4464 & ~i230;
assign a5682 = ~a5680 & ~a5678;
assign a5684 = ~a4624 & ~i232;
assign a5686 = a4624 & i232;
assign a5688 = ~a5686 & ~a5684;
assign a5690 = ~a5688 & ~a5682;
assign a5692 = a5688 & a5682;
assign a5694 = ~a5692 & ~a5690;
assign a5696 = ~a5694 & a5674;
assign a5698 = ~a4624 & i232;
assign a5700 = ~a5698 & ~a5682;
assign a5702 = a4624 & ~i232;
assign a5704 = ~a5702 & ~a5700;
assign a5706 = ~a4784 & ~i234;
assign a5708 = a4784 & i234;
assign a5710 = ~a5708 & ~a5706;
assign a5712 = ~a5710 & ~a5704;
assign a5714 = a5710 & a5704;
assign a5716 = ~a5714 & ~a5712;
assign a5718 = ~a5716 & a5696;
assign a5720 = ~a4784 & i234;
assign a5722 = ~a5720 & ~a5704;
assign a5724 = a4784 & ~i234;
assign a5726 = ~a5724 & ~a5722;
assign a5728 = ~a5726 & ~a4916;
assign a5730 = a5726 & a4916;
assign a5732 = ~a5730 & ~a5728;
assign a5734 = ~a5732 & a5718;
assign a5736 = a5726 & ~a4916;
assign a5738 = ~a5736 & a4946;
assign a5740 = ~a5738 & a5734;
assign a5742 = a5740 & i92;
assign a5744 = ~a5742 & i224;
assign a5746 = ~a5744 & ~l890;
assign a5748 = ~a5746 & ~a5630;
assign a5750 = ~l1020 & l890;
assign a5752 = a5650 & i92;
assign a5754 = ~a4178 & ~i92;
assign a5756 = ~a5754 & ~a5752;
assign a5758 = ~a5756 & ~l890;
assign a5760 = ~a5758 & ~a5750;
assign a5762 = ~l1036 & l890;
assign a5764 = a5650 & ~a5644;
assign a5766 = ~a5650 & a5644;
assign a5768 = ~a5766 & ~a5764;
assign a5770 = ~a5768 & i92;
assign a5772 = ~a4304 & ~i92;
assign a5774 = ~a5772 & ~a5770;
assign a5776 = ~a5774 & ~l890;
assign a5778 = ~a5776 & ~a5762;
assign a5780 = ~l1040 & l890;
assign a5782 = ~a5672 & ~a5652;
assign a5784 = a5672 & a5652;
assign a5786 = ~a5784 & ~a5782;
assign a5788 = ~a5786 & i92;
assign a5790 = ~a4464 & ~i92;
assign a5792 = ~a5790 & ~a5788;
assign a5794 = ~a5792 & ~l890;
assign a5796 = ~a5794 & ~a5780;
assign a5798 = ~l1044 & l890;
assign a5800 = ~a5694 & ~a5674;
assign a5802 = a5694 & a5674;
assign a5804 = ~a5802 & ~a5800;
assign a5806 = ~a5804 & i92;
assign a5808 = ~a4624 & ~i92;
assign a5810 = ~a5808 & ~a5806;
assign a5812 = ~a5810 & ~l890;
assign a5814 = ~a5812 & ~a5798;
assign a5816 = ~l1048 & l890;
assign a5818 = ~a5716 & ~a5696;
assign a5820 = a5716 & a5696;
assign a5822 = ~a5820 & ~a5818;
assign a5824 = ~a5822 & i92;
assign a5826 = ~a4784 & ~i92;
assign a5828 = ~a5826 & ~a5824;
assign a5830 = ~a5828 & ~l890;
assign a5832 = ~a5830 & ~a5816;
assign a5834 = ~l1052 & l890;
assign a5836 = ~a5732 & ~a5718;
assign a5838 = a5732 & a5718;
assign a5840 = ~a5838 & ~a5836;
assign a5842 = ~a5840 & i92;
assign a5844 = ~a4916 & ~i92;
assign a5846 = ~a5844 & ~a5842;
assign a5848 = ~a5846 & ~l890;
assign a5850 = ~a5848 & ~a5834;
assign a5852 = ~l1056 & l890;
assign a5854 = ~a5738 & ~a5734;
assign a5856 = a5738 & a5734;
assign a5858 = ~a5856 & ~a5854;
assign a5860 = ~a5858 & i92;
assign a5862 = ~a4946 & ~i92;
assign a5864 = ~a5862 & ~a5860;
assign a5866 = ~a5864 & ~l890;
assign a5868 = ~a5866 & ~a5852;
assign a5870 = ~l1080 & l890;
assign a5872 = a5742 & ~l890;
assign a5874 = ~a5872 & ~a5870;
assign a5876 = ~a5874 & l1060;
assign a5878 = a5874 & ~l1060;
assign a5880 = ~a5878 & ~a5876;
assign a5882 = ~a5880 & ~a5868;
assign a5884 = a5880 & l1084;
assign a5886 = ~a5880 & ~l1084;
assign a5888 = ~a5886 & ~a5884;
assign a5890 = ~a5888 & a5868;
assign a5892 = ~a5890 & ~a5882;
assign a5894 = ~a5892 & ~a5850;
assign a5896 = ~a5892 & ~l1086;
assign a5898 = a5888 & ~a5868;
assign a5900 = ~a5880 & a5868;
assign a5902 = ~a5900 & ~a5898;
assign a5904 = a5902 & l1086;
assign a5906 = ~a5904 & ~a5896;
assign a5908 = ~a5906 & a5850;
assign a5910 = ~a5908 & ~a5894;
assign a5912 = ~a5910 & ~a5832;
assign a5914 = ~a5910 & ~l1088;
assign a5916 = a5906 & ~a5850;
assign a5918 = ~a5902 & a5850;
assign a5920 = ~a5918 & ~a5916;
assign a5922 = a5920 & l1088;
assign a5924 = ~a5922 & ~a5914;
assign a5926 = ~a5924 & a5832;
assign a5928 = ~a5926 & ~a5912;
assign a5930 = ~a5928 & ~a5814;
assign a5932 = a5924 & ~a5832;
assign a5934 = ~a5920 & a5832;
assign a5936 = ~a5934 & ~a5932;
assign a5938 = a5936 & l1090;
assign a5940 = ~a5928 & ~l1090;
assign a5942 = ~a5940 & ~a5938;
assign a5944 = ~a5942 & a5814;
assign a5946 = ~a5944 & ~a5930;
assign a5948 = ~a5946 & ~a5796;
assign a5950 = a5942 & ~a5814;
assign a5952 = ~a5936 & a5814;
assign a5954 = ~a5952 & ~a5950;
assign a5956 = a5954 & l1092;
assign a5958 = ~a5946 & ~l1092;
assign a5960 = ~a5958 & ~a5956;
assign a5962 = ~a5960 & a5796;
assign a5964 = ~a5962 & ~a5948;
assign a5966 = a5964 & ~a5778;
assign a5968 = a5960 & ~a5796;
assign a5970 = ~a5954 & a5796;
assign a5972 = ~a5970 & ~a5968;
assign a5974 = ~a5972 & a5778;
assign a5976 = ~a5974 & ~a5966;
assign a5978 = a5976 & l1024;
assign a5980 = ~a5964 & ~l1024;
assign a5982 = ~a5980 & ~a5978;
assign a5984 = a5982 & ~a5760;
assign a5986 = ~a5972 & l1024;
assign a5988 = ~a5976 & ~l1024;
assign a5990 = ~a5988 & ~a5986;
assign a5992 = ~a5990 & a5760;
assign a5994 = ~a5992 & ~a5984;
assign a5996 = a5994 & l972;
assign a5998 = ~a5982 & ~l972;
assign a6000 = ~a5998 & ~a5996;
assign a6002 = ~a6000 & ~a5748;
assign a6004 = ~a5892 & l1086;
assign a6006 = ~a5884 & ~a5868;
assign a6008 = ~a5886 & ~l1084;
assign a6010 = ~a6008 & a5868;
assign a6012 = ~a6010 & ~a6006;
assign a6014 = ~a6012 & ~l1086;
assign a6016 = ~a6014 & ~a6004;
assign a6018 = ~a6016 & ~a5850;
assign a6020 = ~a6008 & ~a5868;
assign a6022 = ~a5880 & l1084;
assign a6024 = ~a6022 & a5868;
assign a6026 = ~a6024 & ~a6020;
assign a6028 = ~a6026 & l1086;
assign a6030 = ~a6028 & ~a5896;
assign a6032 = ~a6030 & a5850;
assign a6034 = ~a6032 & ~a6018;
assign a6036 = ~a6034 & ~a5832;
assign a6038 = ~a6030 & ~a5850;
assign a6040 = ~a6026 & ~l1086;
assign a6042 = ~a6040 & ~a5904;
assign a6044 = ~a6042 & a5850;
assign a6046 = ~a6044 & ~a6038;
assign a6048 = ~a6046 & l1088;
assign a6050 = ~a6034 & ~l1088;
assign a6052 = ~a6050 & ~a6048;
assign a6054 = ~a6052 & a5832;
assign a6056 = ~a6054 & ~a6036;
assign a6058 = ~a6056 & ~a5814;
assign a6060 = ~a6052 & ~a5832;
assign a6062 = ~a6046 & a5832;
assign a6064 = ~a6062 & ~a6060;
assign a6066 = ~a6064 & l1090;
assign a6068 = ~a6056 & ~l1090;
assign a6070 = ~a6068 & ~a6066;
assign a6072 = ~a6070 & a5814;
assign a6074 = ~a6072 & ~a6058;
assign a6076 = ~a6074 & ~a5796;
assign a6078 = ~a6070 & ~a5814;
assign a6080 = ~a6064 & a5814;
assign a6082 = ~a6080 & ~a6078;
assign a6084 = ~a6082 & l1092;
assign a6086 = ~a6074 & ~l1092;
assign a6088 = ~a6086 & ~a6084;
assign a6090 = ~a6088 & a5796;
assign a6092 = ~a6090 & ~a6076;
assign a6094 = ~a6092 & ~a5778;
assign a6096 = ~a6088 & ~a5796;
assign a6098 = ~a6082 & a5796;
assign a6100 = ~a6098 & ~a6096;
assign a6102 = ~a6100 & a5778;
assign a6104 = ~a6102 & ~a6094;
assign a6106 = ~a6104 & l1024;
assign a6108 = ~a6092 & ~l1024;
assign a6110 = ~a6108 & ~a6106;
assign a6112 = ~a6110 & ~a5760;
assign a6114 = ~a5910 & l1088;
assign a6116 = ~a6114 & ~a6050;
assign a6118 = ~a6116 & ~a5832;
assign a6120 = ~a6048 & ~a5914;
assign a6122 = ~a6120 & a5832;
assign a6124 = ~a6122 & ~a6118;
assign a6126 = ~a6124 & l1090;
assign a6128 = ~a6126 & ~a6068;
assign a6130 = ~a6128 & ~a5814;
assign a6132 = ~a6124 & ~l1090;
assign a6134 = ~a6132 & ~a6066;
assign a6136 = ~a6134 & a5814;
assign a6138 = ~a6136 & ~a6130;
assign a6140 = ~a6138 & l1092;
assign a6142 = ~a6140 & ~a6086;
assign a6144 = ~a6142 & ~a5796;
assign a6146 = ~a6138 & ~l1092;
assign a6148 = ~a6146 & ~a6084;
assign a6150 = ~a6148 & a5796;
assign a6152 = ~a6150 & ~a6144;
assign a6154 = ~a6152 & ~a5778;
assign a6156 = ~a6154 & ~a6102;
assign a6158 = ~a6156 & l1024;
assign a6160 = ~a6152 & a5778;
assign a6162 = ~a6160 & ~a6094;
assign a6164 = ~a6162 & ~l1024;
assign a6166 = ~a6164 & ~a6158;
assign a6168 = ~a6166 & a5760;
assign a6170 = ~a6168 & ~a6112;
assign a6172 = ~a6170 & l972;
assign a6174 = ~a6162 & l1024;
assign a6176 = ~a6074 & l1092;
assign a6178 = ~a6056 & l1090;
assign a6180 = ~a6034 & l1088;
assign a6182 = ~a5902 & ~l1086;
assign a6184 = ~a6182 & ~a6004;
assign a6186 = ~a6184 & ~a5850;
assign a6188 = ~a5892 & a5850;
assign a6190 = ~a6188 & ~a6186;
assign a6192 = ~a6190 & ~l1088;
assign a6194 = ~a6192 & ~a6180;
assign a6196 = ~a6194 & ~a5832;
assign a6198 = ~a6116 & a5832;
assign a6200 = ~a6198 & ~a6196;
assign a6202 = ~a6200 & ~l1090;
assign a6204 = ~a6202 & ~a6178;
assign a6206 = ~a6204 & ~a5814;
assign a6208 = ~a6128 & a5814;
assign a6210 = ~a6208 & ~a6206;
assign a6212 = ~a6210 & ~l1092;
assign a6214 = ~a6212 & ~a6176;
assign a6216 = ~a6214 & ~a5796;
assign a6218 = ~a6142 & a5796;
assign a6220 = ~a6218 & ~a6216;
assign a6222 = ~a6220 & ~a5778;
assign a6224 = ~a6092 & a5778;
assign a6226 = ~a6224 & ~a6222;
assign a6228 = ~a6226 & ~l1024;
assign a6230 = ~a6228 & ~a6174;
assign a6232 = ~a6230 & ~a5760;
assign a6234 = ~a6110 & a5760;
assign a6236 = ~a6234 & ~a6232;
assign a6238 = ~a6236 & ~l972;
assign a6240 = ~a6238 & ~a6172;
assign a6242 = ~a6240 & a5748;
assign a6244 = ~a6242 & ~a6002;
assign a6246 = ~a6244 & ~l886;
assign a6248 = ~l1018 & l890;
assign a6250 = a5346 & i134;
assign a6252 = a6250 & ~l890;
assign a6254 = ~a6252 & ~a6248;
assign a6256 = ~l1038 & l890;
assign a6258 = a5346 & i136;
assign a6260 = a6258 & ~l890;
assign a6262 = ~a6260 & ~a6256;
assign a6264 = ~l1042 & l890;
assign a6266 = a5346 & i138;
assign a6268 = a6266 & ~l890;
assign a6270 = ~a6268 & ~a6264;
assign a6272 = ~l1046 & l890;
assign a6274 = a5346 & i140;
assign a6276 = a6274 & ~l890;
assign a6278 = ~a6276 & ~a6272;
assign a6280 = ~l1050 & l890;
assign a6282 = a5346 & i142;
assign a6284 = a6282 & ~l890;
assign a6286 = ~a6284 & ~a6280;
assign a6288 = l1060 & l978;
assign a6290 = ~l1060 & ~l978;
assign a6292 = ~a6290 & ~a6288;
assign a6294 = a6292 & l1058;
assign a6296 = ~a6292 & ~l1058;
assign a6298 = ~a6296 & ~a6294;
assign a6300 = a6298 & l1084;
assign a6302 = ~a6292 & ~l1084;
assign a6304 = ~a6302 & ~a6300;
assign a6306 = a6304 & l1054;
assign a6308 = ~a6292 & l1084;
assign a6310 = ~a6298 & ~l1084;
assign a6312 = ~a6310 & ~a6308;
assign a6314 = ~a6312 & ~l1054;
assign a6316 = ~a6314 & ~a6306;
assign a6318 = a6316 & l1086;
assign a6320 = ~a6304 & ~l1086;
assign a6322 = ~a6320 & ~a6318;
assign a6324 = a6322 & ~a6286;
assign a6326 = ~a6312 & l1086;
assign a6328 = ~a6316 & ~l1086;
assign a6330 = ~a6328 & ~a6326;
assign a6332 = ~a6330 & a6286;
assign a6334 = ~a6332 & ~a6324;
assign a6336 = a6334 & l1088;
assign a6338 = ~a6322 & ~l1088;
assign a6340 = ~a6338 & ~a6336;
assign a6342 = a6340 & ~a6278;
assign a6344 = ~a6330 & l1088;
assign a6346 = ~a6334 & ~l1088;
assign a6348 = ~a6346 & ~a6344;
assign a6350 = ~a6348 & a6278;
assign a6352 = ~a6350 & ~a6342;
assign a6354 = a6352 & l1090;
assign a6356 = ~a6340 & ~l1090;
assign a6358 = ~a6356 & ~a6354;
assign a6360 = a6358 & ~a6270;
assign a6362 = ~a6348 & l1090;
assign a6364 = ~a6352 & ~l1090;
assign a6366 = ~a6364 & ~a6362;
assign a6368 = ~a6366 & a6270;
assign a6370 = ~a6368 & ~a6360;
assign a6372 = a6370 & l1092;
assign a6374 = ~a6358 & ~l1092;
assign a6376 = ~a6374 & ~a6372;
assign a6378 = a6376 & ~a6262;
assign a6380 = ~a6366 & l1092;
assign a6382 = ~a6370 & ~l1092;
assign a6384 = ~a6382 & ~a6380;
assign a6386 = ~a6384 & a6262;
assign a6388 = ~a6386 & ~a6378;
assign a6390 = a6388 & l1024;
assign a6392 = ~a6376 & ~l1024;
assign a6394 = ~a6392 & ~a6390;
assign a6396 = a6394 & ~a6254;
assign a6398 = ~a6384 & l1024;
assign a6400 = ~a6388 & ~l1024;
assign a6402 = ~a6400 & ~a6398;
assign a6404 = ~a6402 & a6254;
assign a6406 = ~a6404 & ~a6396;
assign a6408 = a6406 & l972;
assign a6410 = ~a6394 & ~l972;
assign a6412 = ~a6410 & ~a6408;
assign a6414 = ~a6412 & l886;
assign a6416 = ~a6414 & ~a6246;
assign a6418 = ~a6416 & ~l970;
assign a6420 = ~l1094 & l890;
assign a6422 = a5370 & a4980;
assign a6424 = a6422 & ~l890;
assign a6426 = ~a6424 & ~a6420;
assign a6428 = ~l1106 & l890;
assign a6430 = a5370 & a5028;
assign a6432 = a6430 & ~l890;
assign a6434 = ~a6432 & ~a6428;
assign a6436 = ~l1114 & l890;
assign a6438 = a5370 & a5076;
assign a6440 = a6438 & ~l890;
assign a6442 = ~a6440 & ~a6436;
assign a6444 = ~l1122 & l890;
assign a6446 = a5370 & a5124;
assign a6448 = a6446 & ~l890;
assign a6450 = ~a6448 & ~a6444;
assign a6452 = l1166 & l1164;
assign a6454 = ~a6452 & l1166;
assign a6456 = ~a6454 & ~l1170;
assign a6458 = ~a6452 & l1170;
assign a6460 = ~a6458 & ~a6456;
assign a6462 = a6460 & l1168;
assign a6464 = ~l1166 & ~l1164;
assign a6466 = a6464 & ~l1170;
assign a6468 = ~a6464 & ~l1166;
assign a6470 = a6468 & l1170;
assign a6472 = ~a6470 & ~a6466;
assign a6474 = ~a6472 & ~l1168;
assign a6476 = ~a6474 & ~a6462;
assign a6478 = a6476 & l1162;
assign a6480 = ~a6478 & l1162;
assign a6482 = a6480 & l1160;
assign a6484 = ~a6476 & ~l1162;
assign a6486 = a6484 & ~l1160;
assign a6488 = ~a6486 & ~a6482;
assign a6490 = a6488 & l1148;
assign a6492 = ~a6490 & l1148;
assign a6494 = a6492 & l1146;
assign a6496 = ~a6488 & ~l1148;
assign a6498 = a6496 & ~l1146;
assign a6500 = ~a6498 & ~a6494;
assign a6502 = a6500 & ~l896;
assign a6504 = ~a6468 & ~l1162;
assign a6506 = ~a6504 & ~l1162;
assign a6508 = ~a6506 & l1216;
assign a6510 = ~a6454 & ~l1162;
assign a6512 = ~a6510 & ~l1162;
assign a6514 = ~a6512 & ~l1216;
assign a6516 = ~a6514 & ~a6508;
assign a6518 = ~a6516 & l1200;
assign a6520 = ~a6454 & l1162;
assign a6522 = ~a6520 & l1162;
assign a6524 = ~a6522 & l1216;
assign a6526 = ~a6464 & l1162;
assign a6528 = ~a6526 & l1162;
assign a6530 = ~a6528 & ~l1216;
assign a6532 = ~a6530 & ~a6524;
assign a6534 = ~a6532 & ~l1232;
assign a6536 = a6512 & l1216;
assign a6538 = a6464 & ~l1162;
assign a6540 = a6538 & ~l1216;
assign a6542 = ~a6540 & ~a6536;
assign a6544 = a6542 & l1232;
assign a6546 = ~a6544 & ~a6534;
assign a6548 = ~a6546 & ~l1200;
assign a6550 = ~a6548 & ~a6518;
assign a6552 = ~a6550 & ~l1148;
assign a6554 = ~a6552 & ~l1148;
assign a6556 = ~a6554 & l1176;
assign a6558 = ~a6452 & l1162;
assign a6560 = ~a6558 & l1162;
assign a6562 = ~a6560 & l1216;
assign a6564 = ~a6468 & l1162;
assign a6566 = ~a6564 & l1162;
assign a6568 = ~a6566 & ~l1216;
assign a6570 = ~a6568 & ~a6562;
assign a6572 = ~a6570 & l1232;
assign a6574 = ~a6572 & ~a6534;
assign a6576 = a6574 & l1200;
assign a6578 = ~a6452 & ~l1162;
assign a6580 = ~a6578 & ~l1162;
assign a6582 = ~a6580 & l1216;
assign a6584 = ~a6506 & ~l1216;
assign a6586 = ~a6584 & ~a6582;
assign a6588 = a6586 & l1232;
assign a6590 = ~a6542 & ~l1232;
assign a6592 = ~a6590 & ~a6588;
assign a6594 = ~a6592 & ~l1200;
assign a6596 = ~a6594 & ~a6576;
assign a6598 = a6596 & l1148;
assign a6600 = ~a6598 & l1148;
assign a6602 = ~a6600 & ~l1176;
assign a6604 = ~a6602 & ~a6556;
assign a6606 = ~a6604 & l1172;
assign a6608 = a6500 & ~l1172;
assign a6610 = ~a6608 & ~a6606;
assign a6612 = ~a6610 & l896;
assign a6614 = ~a6612 & ~a6502;
assign a6616 = ~a6614 & ~l898;
assign a6618 = ~a6506 & l1218;
assign a6620 = ~a6512 & ~l1218;
assign a6622 = ~a6620 & ~a6618;
assign a6624 = ~a6622 & l1202;
assign a6626 = ~a6522 & l1218;
assign a6628 = ~a6528 & ~l1218;
assign a6630 = ~a6628 & ~a6626;
assign a6632 = ~a6630 & ~l1234;
assign a6634 = a6512 & l1218;
assign a6636 = a6538 & ~l1218;
assign a6638 = ~a6636 & ~a6634;
assign a6640 = a6638 & l1234;
assign a6642 = ~a6640 & ~a6632;
assign a6644 = ~a6642 & ~l1202;
assign a6646 = ~a6644 & ~a6624;
assign a6648 = ~a6646 & ~l1148;
assign a6650 = ~a6648 & ~l1148;
assign a6652 = ~a6650 & l1178;
assign a6654 = ~a6560 & l1218;
assign a6656 = ~a6566 & ~l1218;
assign a6658 = ~a6656 & ~a6654;
assign a6660 = ~a6658 & l1234;
assign a6662 = ~a6660 & ~a6632;
assign a6664 = a6662 & l1202;
assign a6666 = ~a6580 & l1218;
assign a6668 = ~a6506 & ~l1218;
assign a6670 = ~a6668 & ~a6666;
assign a6672 = a6670 & l1234;
assign a6674 = ~a6638 & ~l1234;
assign a6676 = ~a6674 & ~a6672;
assign a6678 = ~a6676 & ~l1202;
assign a6680 = ~a6678 & ~a6664;
assign a6682 = a6680 & l1148;
assign a6684 = ~a6682 & l1148;
assign a6686 = ~a6684 & ~l1178;
assign a6688 = ~a6686 & ~a6652;
assign a6690 = ~a6688 & ~l1172;
assign a6692 = ~a6690 & ~a6606;
assign a6694 = ~a6692 & l928;
assign a6696 = ~a6614 & ~l928;
assign a6698 = ~a6696 & ~a6694;
assign a6700 = ~a6698 & l898;
assign a6702 = ~a6700 & ~a6616;
assign a6704 = ~a6702 & ~l900;
assign a6706 = ~a6702 & ~l930;
assign a6708 = ~a6470 & ~l1168;
assign a6710 = ~a6708 & ~l1168;
assign a6712 = ~a6710 & ~l1162;
assign a6714 = ~a6712 & ~l1162;
assign a6716 = ~a6714 & l1220;
assign a6718 = ~a6456 & ~l1170;
assign a6720 = ~a6718 & l1168;
assign a6722 = ~a6720 & l1168;
assign a6724 = ~a6722 & ~l1162;
assign a6726 = ~a6724 & ~l1162;
assign a6728 = ~a6726 & ~l1220;
assign a6730 = ~a6728 & ~a6716;
assign a6732 = ~a6730 & ~l1160;
assign a6734 = ~a6732 & ~l1160;
assign a6736 = ~a6734 & l1204;
assign a6738 = ~a6722 & l1162;
assign a6740 = ~a6738 & l1162;
assign a6742 = ~a6740 & l1220;
assign a6744 = a6466 & ~l1168;
assign a6746 = ~a6744 & l1162;
assign a6748 = ~a6746 & l1162;
assign a6750 = ~a6748 & ~l1220;
assign a6752 = ~a6750 & ~a6742;
assign a6754 = ~a6752 & l1160;
assign a6756 = ~a6754 & l1160;
assign a6758 = ~a6756 & ~l1236;
assign a6760 = a6726 & l1220;
assign a6762 = a6744 & ~l1162;
assign a6764 = a6762 & ~l1220;
assign a6766 = ~a6764 & ~a6760;
assign a6768 = ~a6766 & ~l1160;
assign a6770 = ~a6768 & l1236;
assign a6772 = ~a6770 & ~a6758;
assign a6774 = ~a6772 & ~l1204;
assign a6776 = ~a6774 & ~a6736;
assign a6778 = ~a6776 & ~l1148;
assign a6780 = ~a6778 & ~l1148;
assign a6782 = ~a6780 & ~l1146;
assign a6784 = ~a6782 & ~l1146;
assign a6786 = ~a6784 & l1180;
assign a6788 = ~a6458 & l1170;
assign a6790 = ~a6788 & l1168;
assign a6792 = ~a6790 & l1168;
assign a6794 = ~a6792 & l1162;
assign a6796 = ~a6794 & l1162;
assign a6798 = ~a6796 & l1220;
assign a6800 = ~a6710 & l1162;
assign a6802 = ~a6800 & l1162;
assign a6804 = ~a6802 & ~l1220;
assign a6806 = ~a6804 & ~a6798;
assign a6808 = ~a6806 & l1160;
assign a6810 = ~a6808 & l1160;
assign a6812 = ~a6810 & l1236;
assign a6814 = ~a6812 & ~a6758;
assign a6816 = a6814 & l1204;
assign a6818 = ~a6792 & ~l1162;
assign a6820 = ~a6818 & ~l1162;
assign a6822 = ~a6820 & l1220;
assign a6824 = ~a6714 & ~l1220;
assign a6826 = ~a6824 & ~a6822;
assign a6828 = ~a6826 & ~l1160;
assign a6830 = ~a6828 & ~l1160;
assign a6832 = a6830 & l1236;
assign a6834 = a6768 & ~l1236;
assign a6836 = ~a6834 & ~a6832;
assign a6838 = ~a6836 & ~l1204;
assign a6840 = ~a6838 & ~a6816;
assign a6842 = a6840 & l1148;
assign a6844 = ~a6842 & l1148;
assign a6846 = ~a6844 & l1146;
assign a6848 = ~a6846 & l1146;
assign a6850 = ~a6848 & ~l1180;
assign a6852 = ~a6850 & ~a6786;
assign a6854 = ~a6852 & ~l1172;
assign a6856 = ~a6714 & l1216;
assign a6858 = ~a6726 & ~l1216;
assign a6860 = ~a6858 & ~a6856;
assign a6862 = ~a6860 & ~l1160;
assign a6864 = ~a6862 & ~l1160;
assign a6866 = ~a6864 & l1200;
assign a6868 = ~a6740 & l1216;
assign a6870 = ~a6748 & ~l1216;
assign a6872 = ~a6870 & ~a6868;
assign a6874 = ~a6872 & l1160;
assign a6876 = ~a6874 & l1160;
assign a6878 = ~a6876 & ~l1232;
assign a6880 = a6726 & l1216;
assign a6882 = a6762 & ~l1216;
assign a6884 = ~a6882 & ~a6880;
assign a6886 = ~a6884 & ~l1160;
assign a6888 = ~a6886 & l1232;
assign a6890 = ~a6888 & ~a6878;
assign a6892 = ~a6890 & ~l1200;
assign a6894 = ~a6892 & ~a6866;
assign a6896 = ~a6894 & ~l1148;
assign a6898 = ~a6896 & ~l1148;
assign a6900 = ~a6898 & ~l1146;
assign a6902 = ~a6900 & ~l1146;
assign a6904 = ~a6902 & l1176;
assign a6906 = ~a6796 & l1216;
assign a6908 = ~a6802 & ~l1216;
assign a6910 = ~a6908 & ~a6906;
assign a6912 = ~a6910 & l1160;
assign a6914 = ~a6912 & l1160;
assign a6916 = ~a6914 & l1232;
assign a6918 = ~a6916 & ~a6878;
assign a6920 = a6918 & l1200;
assign a6922 = ~a6820 & l1216;
assign a6924 = ~a6714 & ~l1216;
assign a6926 = ~a6924 & ~a6922;
assign a6928 = ~a6926 & ~l1160;
assign a6930 = ~a6928 & ~l1160;
assign a6932 = a6930 & l1232;
assign a6934 = a6886 & ~l1232;
assign a6936 = ~a6934 & ~a6932;
assign a6938 = ~a6936 & ~l1200;
assign a6940 = ~a6938 & ~a6920;
assign a6942 = a6940 & l1148;
assign a6944 = ~a6942 & l1148;
assign a6946 = ~a6944 & l1146;
assign a6948 = ~a6946 & l1146;
assign a6950 = ~a6948 & ~l1176;
assign a6952 = ~a6950 & ~a6904;
assign a6954 = ~a6952 & l1172;
assign a6956 = ~a6954 & ~a6854;
assign a6958 = ~a6956 & ~l896;
assign a6960 = ~a6854 & ~a6606;
assign a6962 = ~a6960 & l896;
assign a6964 = ~a6962 & ~a6958;
assign a6966 = ~a6964 & ~l928;
assign a6968 = ~a6714 & l1218;
assign a6970 = ~a6726 & ~l1218;
assign a6972 = ~a6970 & ~a6968;
assign a6974 = ~a6972 & ~l1160;
assign a6976 = ~a6974 & ~l1160;
assign a6978 = ~a6976 & l1202;
assign a6980 = ~a6740 & l1218;
assign a6982 = ~a6748 & ~l1218;
assign a6984 = ~a6982 & ~a6980;
assign a6986 = ~a6984 & l1160;
assign a6988 = ~a6986 & l1160;
assign a6990 = ~a6988 & ~l1234;
assign a6992 = a6726 & l1218;
assign a6994 = a6762 & ~l1218;
assign a6996 = ~a6994 & ~a6992;
assign a6998 = ~a6996 & ~l1160;
assign a7000 = ~a6998 & l1234;
assign a7002 = ~a7000 & ~a6990;
assign a7004 = ~a7002 & ~l1202;
assign a7006 = ~a7004 & ~a6978;
assign a7008 = ~a7006 & ~l1148;
assign a7010 = ~a7008 & ~l1148;
assign a7012 = ~a7010 & ~l1146;
assign a7014 = ~a7012 & ~l1146;
assign a7016 = ~a7014 & l1178;
assign a7018 = ~a6796 & l1218;
assign a7020 = ~a6802 & ~l1218;
assign a7022 = ~a7020 & ~a7018;
assign a7024 = ~a7022 & l1160;
assign a7026 = ~a7024 & l1160;
assign a7028 = ~a7026 & l1234;
assign a7030 = ~a7028 & ~a6990;
assign a7032 = a7030 & l1202;
assign a7034 = ~a6820 & l1218;
assign a7036 = ~a6714 & ~l1218;
assign a7038 = ~a7036 & ~a7034;
assign a7040 = ~a7038 & ~l1160;
assign a7042 = ~a7040 & ~l1160;
assign a7044 = a7042 & l1234;
assign a7046 = a6998 & ~l1234;
assign a7048 = ~a7046 & ~a7044;
assign a7050 = ~a7048 & ~l1202;
assign a7052 = ~a7050 & ~a7032;
assign a7054 = a7052 & l1148;
assign a7056 = ~a7054 & l1148;
assign a7058 = ~a7056 & l1146;
assign a7060 = ~a7058 & l1146;
assign a7062 = ~a7060 & ~l1178;
assign a7064 = ~a7062 & ~a7016;
assign a7066 = ~a7064 & ~l1172;
assign a7068 = ~a7066 & ~a6954;
assign a7070 = ~a7068 & ~l896;
assign a7072 = ~a7066 & ~a6606;
assign a7074 = ~a7072 & l896;
assign a7076 = ~a7074 & ~a7070;
assign a7078 = ~a7076 & l928;
assign a7080 = ~a7078 & ~a6966;
assign a7082 = ~a7080 & ~l898;
assign a7084 = ~a6966 & ~a6694;
assign a7086 = ~a7084 & l898;
assign a7088 = ~a7086 & ~a7082;
assign a7090 = ~a7088 & l930;
assign a7092 = ~a7090 & ~a6706;
assign a7094 = ~a7092 & l900;
assign a7096 = ~a7094 & ~a6704;
assign a7098 = a7096 & l1060;
assign a7100 = ~a7098 & l1060;
assign a7102 = a7100 & l1082;
assign a7104 = ~a7096 & ~l1060;
assign a7106 = a7104 & ~l1082;
assign a7108 = ~a7106 & ~a7102;
assign a7110 = ~a7108 & l1138;
assign a7112 = ~a7104 & l1082;
assign a7114 = ~a7100 & ~l1082;
assign a7116 = ~a7114 & ~a7112;
assign a7118 = a7116 & l1084;
assign a7120 = ~a7108 & ~l1084;
assign a7122 = ~a7120 & ~a7118;
assign a7124 = ~a7122 & ~l1138;
assign a7126 = ~a7124 & ~a7110;
assign a7128 = ~a7126 & l1130;
assign a7130 = a7122 & l1138;
assign a7132 = ~a7116 & ~l1138;
assign a7134 = ~a7132 & ~a7130;
assign a7136 = a7134 & l1086;
assign a7138 = ~a7126 & ~l1086;
assign a7140 = ~a7138 & ~a7136;
assign a7142 = ~a7140 & ~l1130;
assign a7144 = ~a7142 & ~a7128;
assign a7146 = ~a7144 & ~a6450;
assign a7148 = a7140 & l1130;
assign a7150 = ~a7134 & ~l1130;
assign a7152 = ~a7150 & ~a7148;
assign a7154 = a7152 & l1088;
assign a7156 = ~a7144 & ~l1088;
assign a7158 = ~a7156 & ~a7154;
assign a7160 = ~a7158 & a6450;
assign a7162 = ~a7160 & ~a7146;
assign a7164 = ~a7162 & ~a6442;
assign a7166 = a7158 & ~a6450;
assign a7168 = ~a7152 & a6450;
assign a7170 = ~a7168 & ~a7166;
assign a7172 = a7170 & l1090;
assign a7174 = ~a7162 & ~l1090;
assign a7176 = ~a7174 & ~a7172;
assign a7178 = ~a7176 & a6442;
assign a7180 = ~a7178 & ~a7164;
assign a7182 = ~a7180 & ~a6434;
assign a7184 = a7176 & ~a6442;
assign a7186 = ~a7170 & a6442;
assign a7188 = ~a7186 & ~a7184;
assign a7190 = a7188 & l1092;
assign a7192 = ~a7180 & ~l1092;
assign a7194 = ~a7192 & ~a7190;
assign a7196 = ~a7194 & a6434;
assign a7198 = ~a7196 & ~a7182;
assign a7200 = a7198 & ~a6426;
assign a7202 = a7194 & ~a6434;
assign a7204 = ~a7188 & a6434;
assign a7206 = ~a7204 & ~a7202;
assign a7208 = ~a7206 & a6426;
assign a7210 = ~a7208 & ~a7200;
assign a7212 = a7210 & l1024;
assign a7214 = ~a7198 & ~l1024;
assign a7216 = ~a7214 & ~a7212;
assign a7218 = ~a7216 & l972;
assign a7220 = ~l1022 & l890;
assign a7222 = a5370 & a3976;
assign a7224 = a7222 & ~l890;
assign a7226 = ~a7224 & ~a7220;
assign a7228 = ~a7198 & l1024;
assign a7230 = ~a7180 & l1092;
assign a7232 = ~a7162 & l1090;
assign a7234 = ~a7144 & l1088;
assign a7236 = ~a7126 & l1086;
assign a7238 = a7108 & l1084;
assign a7240 = ~a7116 & ~l1084;
assign a7242 = ~a7240 & ~a7238;
assign a7244 = a7242 & l1138;
assign a7246 = ~a7108 & ~l1138;
assign a7248 = ~a7246 & ~a7244;
assign a7250 = ~a7248 & ~l1086;
assign a7252 = ~a7250 & ~a7236;
assign a7254 = ~a7252 & l1130;
assign a7256 = ~a7126 & ~l1130;
assign a7258 = ~a7256 & ~a7254;
assign a7260 = ~a7258 & ~l1088;
assign a7262 = ~a7260 & ~a7234;
assign a7264 = ~a7262 & ~a6450;
assign a7266 = ~a7144 & a6450;
assign a7268 = ~a7266 & ~a7264;
assign a7270 = ~a7268 & ~l1090;
assign a7272 = ~a7270 & ~a7232;
assign a7274 = ~a7272 & ~a6442;
assign a7276 = ~a7162 & a6442;
assign a7278 = ~a7276 & ~a7274;
assign a7280 = ~a7278 & ~l1092;
assign a7282 = ~a7280 & ~a7230;
assign a7284 = ~a7282 & ~a6434;
assign a7286 = ~a7180 & a6434;
assign a7288 = ~a7286 & ~a7284;
assign a7290 = ~a7288 & ~a6426;
assign a7292 = ~a7198 & a6426;
assign a7294 = ~a7292 & ~a7290;
assign a7296 = ~a7294 & ~l1024;
assign a7298 = ~a7296 & ~a7228;
assign a7300 = ~a7298 & ~a7226;
assign a7302 = a7226 & ~a7216;
assign a7304 = ~a7302 & ~a7300;
assign a7306 = ~a7304 & ~l972;
assign a7308 = ~a7306 & ~a7218;
assign a7310 = ~a7308 & l948;
assign a7312 = ~l1214 & l890;
assign a7314 = ~a2718 & ~l890;
assign a7316 = ~a7314 & ~a7312;
assign a7318 = ~l1230 & l890;
assign a7320 = ~a2728 & ~l890;
assign a7322 = ~a7320 & ~a7318;
assign a7324 = ~l1158 & l890;
assign a7326 = a4140 & ~l890;
assign a7328 = ~a7326 & ~a7324;
assign a7330 = ~a6560 & l1246;
assign a7332 = ~a6522 & ~l1246;
assign a7334 = ~a7332 & ~a7330;
assign a7336 = ~a7334 & ~a7328;
assign a7338 = ~a6566 & l1246;
assign a7340 = ~a6528 & ~l1246;
assign a7342 = ~a7340 & ~a7338;
assign a7344 = ~a7342 & a7328;
assign a7346 = ~a7344 & ~a7336;
assign a7348 = a7346 & ~a7322;
assign a7350 = ~a6580 & l1246;
assign a7352 = ~a6512 & ~l1246;
assign a7354 = ~a7352 & ~a7350;
assign a7356 = a7354 & ~a7328;
assign a7358 = a6506 & l1246;
assign a7360 = a6538 & ~l1246;
assign a7362 = ~a7360 & ~a7358;
assign a7364 = ~a7362 & a7328;
assign a7366 = ~a7364 & ~a7356;
assign a7368 = ~a7366 & a7322;
assign a7370 = ~a7368 & ~a7348;
assign a7372 = a7370 & l1148;
assign a7374 = ~a7372 & l1148;
assign a7376 = a7374 & ~a7316;
assign a7378 = ~a7370 & ~l1148;
assign a7380 = a7378 & a7316;
assign a7382 = ~a7380 & ~a7376;
assign a7384 = ~a7382 & l1060;
assign a7386 = ~a7384 & l1060;
assign a7388 = ~a7386 & ~a5874;
assign a7390 = ~a7382 & ~l1060;
assign a7392 = ~a7390 & ~l1060;
assign a7394 = ~a7392 & a5874;
assign a7396 = ~a7394 & ~a7388;
assign a7398 = ~a7396 & ~a5868;
assign a7400 = ~a7392 & ~a5874;
assign a7402 = ~a7386 & a5874;
assign a7404 = ~a7402 & ~a7400;
assign a7406 = ~a7404 & l1084;
assign a7408 = ~a7396 & ~l1084;
assign a7410 = ~a7408 & ~a7406;
assign a7412 = ~a7410 & a5868;
assign a7414 = ~a7412 & ~a7398;
assign a7416 = ~a7414 & ~a5850;
assign a7418 = ~a7410 & ~a5868;
assign a7420 = ~a7404 & a5868;
assign a7422 = ~a7420 & ~a7418;
assign a7424 = ~a7422 & l1086;
assign a7426 = ~a7414 & ~l1086;
assign a7428 = ~a7426 & ~a7424;
assign a7430 = ~a7428 & a5850;
assign a7432 = ~a7430 & ~a7416;
assign a7434 = ~a7432 & ~a5832;
assign a7436 = ~a7428 & ~a5850;
assign a7438 = ~a7422 & a5850;
assign a7440 = ~a7438 & ~a7436;
assign a7442 = ~a7440 & l1088;
assign a7444 = ~a7432 & ~l1088;
assign a7446 = ~a7444 & ~a7442;
assign a7448 = ~a7446 & a5832;
assign a7450 = ~a7448 & ~a7434;
assign a7452 = ~a7450 & ~a5814;
assign a7454 = ~a7446 & ~a5832;
assign a7456 = ~a7440 & a5832;
assign a7458 = ~a7456 & ~a7454;
assign a7460 = ~a7458 & l1090;
assign a7462 = ~a7450 & ~l1090;
assign a7464 = ~a7462 & ~a7460;
assign a7466 = ~a7464 & a5814;
assign a7468 = ~a7466 & ~a7452;
assign a7470 = ~a7468 & ~a5796;
assign a7472 = ~a7464 & ~a5814;
assign a7474 = ~a7458 & a5814;
assign a7476 = ~a7474 & ~a7472;
assign a7478 = ~a7476 & l1092;
assign a7480 = ~a7468 & ~l1092;
assign a7482 = ~a7480 & ~a7478;
assign a7484 = ~a7482 & a5796;
assign a7486 = ~a7484 & ~a7470;
assign a7488 = ~a7486 & ~a5778;
assign a7490 = ~a7482 & ~a5796;
assign a7492 = ~a7476 & a5796;
assign a7494 = ~a7492 & ~a7490;
assign a7496 = ~a7494 & a5778;
assign a7498 = ~a7496 & ~a7488;
assign a7500 = ~a7498 & l1024;
assign a7502 = ~a7486 & ~l1024;
assign a7504 = ~a7502 & ~a7500;
assign a7506 = ~a7504 & ~a5760;
assign a7508 = ~a7494 & l1024;
assign a7510 = ~a7498 & ~l1024;
assign a7512 = ~a7510 & ~a7508;
assign a7514 = ~a7512 & a5760;
assign a7516 = ~a7514 & ~a7506;
assign a7518 = ~a7516 & l972;
assign a7520 = ~a7504 & ~l972;
assign a7522 = ~a7520 & ~a7518;
assign a7524 = a7522 & ~a5748;
assign a7526 = ~a6538 & l1246;
assign a7528 = ~a6506 & ~l1246;
assign a7530 = ~a7528 & ~a7526;
assign a7532 = ~a7530 & ~a7328;
assign a7534 = ~a7354 & a7328;
assign a7536 = ~a7534 & ~a7532;
assign a7538 = ~a7536 & ~a7322;
assign a7540 = ~a7526 & ~a7340;
assign a7542 = ~a7540 & a7328;
assign a7544 = ~a7542 & ~a7336;
assign a7546 = ~a7544 & a7322;
assign a7548 = ~a7546 & ~a7538;
assign a7550 = ~a7548 & ~l1148;
assign a7552 = ~a7550 & ~l1148;
assign a7554 = ~a7552 & ~a7316;
assign a7556 = ~a7374 & a7316;
assign a7558 = ~a7556 & ~a7554;
assign a7560 = a7558 & l1060;
assign a7562 = ~a7560 & l1060;
assign a7564 = a7562 & ~a5874;
assign a7566 = ~a7558 & ~l1060;
assign a7568 = a7566 & a5874;
assign a7570 = ~a7568 & ~a7564;
assign a7572 = ~a7570 & ~a5868;
assign a7574 = ~a7566 & ~a5874;
assign a7576 = ~a7562 & a5874;
assign a7578 = ~a7576 & ~a7574;
assign a7580 = a7578 & l1084;
assign a7582 = ~a7570 & ~l1084;
assign a7584 = ~a7582 & ~a7580;
assign a7586 = ~a7584 & a5868;
assign a7588 = ~a7586 & ~a7572;
assign a7590 = ~a7588 & l1086;
assign a7592 = ~a7558 & ~l1084;
assign a7594 = ~a7570 & l1084;
assign a7596 = ~a7594 & ~a7592;
assign a7598 = ~a7596 & ~a5868;
assign a7600 = ~a7558 & l1084;
assign a7602 = ~a7600 & ~a7582;
assign a7604 = ~a7602 & a5868;
assign a7606 = ~a7604 & ~a7598;
assign a7608 = ~a7606 & ~l1086;
assign a7610 = ~a7608 & ~a7590;
assign a7612 = ~a7610 & ~a5850;
assign a7614 = ~a7602 & ~a5868;
assign a7616 = ~a7592 & ~a7580;
assign a7618 = ~a7616 & a5868;
assign a7620 = ~a7618 & ~a7614;
assign a7622 = ~a7620 & l1086;
assign a7624 = ~a7588 & ~l1086;
assign a7626 = ~a7624 & ~a7622;
assign a7628 = ~a7626 & a5850;
assign a7630 = ~a7628 & ~a7612;
assign a7632 = ~a7630 & ~a5832;
assign a7634 = ~a7626 & ~a5850;
assign a7636 = a7584 & ~a5868;
assign a7638 = ~a7578 & a5868;
assign a7640 = ~a7638 & ~a7636;
assign a7642 = a7640 & l1086;
assign a7644 = ~a7620 & ~l1086;
assign a7646 = ~a7644 & ~a7642;
assign a7648 = ~a7646 & a5850;
assign a7650 = ~a7648 & ~a7634;
assign a7652 = ~a7650 & l1088;
assign a7654 = ~a7630 & ~l1088;
assign a7656 = ~a7654 & ~a7652;
assign a7658 = ~a7656 & a5832;
assign a7660 = ~a7658 & ~a7632;
assign a7662 = ~a7660 & ~a5814;
assign a7664 = ~a7656 & ~a5832;
assign a7666 = ~a7650 & a5832;
assign a7668 = ~a7666 & ~a7664;
assign a7670 = ~a7668 & l1090;
assign a7672 = ~a7660 & ~l1090;
assign a7674 = ~a7672 & ~a7670;
assign a7676 = ~a7674 & a5814;
assign a7678 = ~a7676 & ~a7662;
assign a7680 = ~a7678 & ~a5796;
assign a7682 = ~a7674 & ~a5814;
assign a7684 = ~a7668 & a5814;
assign a7686 = ~a7684 & ~a7682;
assign a7688 = ~a7686 & l1092;
assign a7690 = ~a7678 & ~l1092;
assign a7692 = ~a7690 & ~a7688;
assign a7694 = ~a7692 & a5796;
assign a7696 = ~a7694 & ~a7680;
assign a7698 = ~a7696 & ~a5778;
assign a7700 = ~a7692 & ~a5796;
assign a7702 = ~a7686 & a5796;
assign a7704 = ~a7702 & ~a7700;
assign a7706 = ~a7704 & a5778;
assign a7708 = ~a7706 & ~a7698;
assign a7710 = ~a7708 & l1024;
assign a7712 = ~a7696 & ~l1024;
assign a7714 = ~a7712 & ~a7710;
assign a7716 = ~a7714 & ~a5760;
assign a7718 = ~a7588 & ~a5850;
assign a7720 = ~a7642 & ~a7624;
assign a7722 = ~a7720 & a5850;
assign a7724 = ~a7722 & ~a7718;
assign a7726 = ~a7724 & l1088;
assign a7728 = ~a7726 & ~a7654;
assign a7730 = ~a7728 & ~a5832;
assign a7732 = ~a7724 & ~l1088;
assign a7734 = ~a7732 & ~a7652;
assign a7736 = ~a7734 & a5832;
assign a7738 = ~a7736 & ~a7730;
assign a7740 = ~a7738 & l1090;
assign a7742 = ~a7740 & ~a7672;
assign a7744 = ~a7742 & ~a5814;
assign a7746 = ~a7738 & ~l1090;
assign a7748 = ~a7746 & ~a7670;
assign a7750 = ~a7748 & a5814;
assign a7752 = ~a7750 & ~a7744;
assign a7754 = ~a7752 & l1092;
assign a7756 = ~a7754 & ~a7690;
assign a7758 = ~a7756 & ~a5796;
assign a7760 = ~a7752 & ~l1092;
assign a7762 = ~a7760 & ~a7688;
assign a7764 = ~a7762 & a5796;
assign a7766 = ~a7764 & ~a7758;
assign a7768 = ~a7766 & ~a5778;
assign a7770 = ~a7768 & ~a7706;
assign a7772 = ~a7770 & l1024;
assign a7774 = ~a7766 & a5778;
assign a7776 = ~a7774 & ~a7698;
assign a7778 = ~a7776 & ~l1024;
assign a7780 = ~a7778 & ~a7772;
assign a7782 = ~a7780 & a5760;
assign a7784 = ~a7782 & ~a7716;
assign a7786 = ~a7784 & l972;
assign a7788 = ~a7776 & l1024;
assign a7790 = ~a7678 & l1092;
assign a7792 = ~a7660 & l1090;
assign a7794 = ~a7630 & l1088;
assign a7796 = a7570 & l1084;
assign a7798 = ~a7578 & ~l1084;
assign a7800 = ~a7798 & ~a7796;
assign a7802 = a7800 & ~a5868;
assign a7804 = ~a7570 & a5868;
assign a7806 = ~a7804 & ~a7802;
assign a7808 = ~a7806 & ~l1086;
assign a7810 = ~a7808 & ~a7590;
assign a7812 = ~a7810 & ~a5850;
assign a7814 = ~a7588 & a5850;
assign a7816 = ~a7814 & ~a7812;
assign a7818 = ~a7816 & ~l1088;
assign a7820 = ~a7818 & ~a7794;
assign a7822 = ~a7820 & ~a5832;
assign a7824 = ~a7728 & a5832;
assign a7826 = ~a7824 & ~a7822;
assign a7828 = ~a7826 & ~l1090;
assign a7830 = ~a7828 & ~a7792;
assign a7832 = ~a7830 & ~a5814;
assign a7834 = ~a7742 & a5814;
assign a7836 = ~a7834 & ~a7832;
assign a7838 = ~a7836 & ~l1092;
assign a7840 = ~a7838 & ~a7790;
assign a7842 = ~a7840 & ~a5796;
assign a7844 = ~a7756 & a5796;
assign a7846 = ~a7844 & ~a7842;
assign a7848 = ~a7846 & ~a5778;
assign a7850 = ~a7696 & a5778;
assign a7852 = ~a7850 & ~a7848;
assign a7854 = ~a7852 & ~l1024;
assign a7856 = ~a7854 & ~a7788;
assign a7858 = ~a7856 & ~a5760;
assign a7860 = ~a7714 & a5760;
assign a7862 = ~a7860 & ~a7858;
assign a7864 = ~a7862 & ~l972;
assign a7866 = ~a7864 & ~a7786;
assign a7868 = ~a7866 & a5748;
assign a7870 = ~a7868 & ~a7524;
assign a7872 = ~a7870 & ~l948;
assign a7874 = ~a7872 & ~a7310;
assign a7876 = ~a7874 & ~l886;
assign a7878 = ~a6506 & l1002;
assign a7880 = ~a6512 & ~l1002;
assign a7882 = ~a7880 & ~a7878;
assign a7884 = ~a7882 & l1004;
assign a7886 = ~a6522 & l1002;
assign a7888 = ~a6528 & ~l1002;
assign a7890 = ~a7888 & ~a7886;
assign a7892 = ~a7890 & ~l1006;
assign a7894 = a6512 & l1002;
assign a7896 = a6538 & ~l1002;
assign a7898 = ~a7896 & ~a7894;
assign a7900 = a7898 & l1006;
assign a7902 = ~a7900 & ~a7892;
assign a7904 = ~a7902 & ~l1004;
assign a7906 = ~a7904 & ~a7884;
assign a7908 = ~a7906 & ~l1148;
assign a7910 = ~a7908 & ~l1148;
assign a7912 = ~a7910 & l880;
assign a7914 = ~a6560 & l1002;
assign a7916 = ~a6566 & ~l1002;
assign a7918 = ~a7916 & ~a7914;
assign a7920 = ~a7918 & l1006;
assign a7922 = ~a7920 & ~a7892;
assign a7924 = a7922 & l1004;
assign a7926 = ~a6580 & l1002;
assign a7928 = ~a6506 & ~l1002;
assign a7930 = ~a7928 & ~a7926;
assign a7932 = a7930 & l1006;
assign a7934 = ~a7898 & ~l1006;
assign a7936 = ~a7934 & ~a7932;
assign a7938 = ~a7936 & ~l1004;
assign a7940 = ~a7938 & ~a7924;
assign a7942 = a7940 & l1148;
assign a7944 = ~a7942 & l1148;
assign a7946 = ~a7944 & ~l880;
assign a7948 = ~a7946 & ~a7912;
assign a7950 = a7948 & l1060;
assign a7952 = ~a7950 & l1060;
assign a7954 = a7952 & l978;
assign a7956 = ~a7948 & ~l1060;
assign a7958 = a7956 & ~l978;
assign a7960 = ~a7958 & ~a7954;
assign a7962 = a7960 & l1058;
assign a7964 = ~a7956 & l978;
assign a7966 = ~a7952 & ~l978;
assign a7968 = ~a7966 & ~a7964;
assign a7970 = ~a7968 & ~l1058;
assign a7972 = ~a7970 & ~a7962;
assign a7974 = a7972 & l1084;
assign a7976 = ~a7960 & ~l1084;
assign a7978 = ~a7976 & ~a7974;
assign a7980 = a7978 & l1054;
assign a7982 = ~a7968 & l1084;
assign a7984 = ~a7972 & ~l1084;
assign a7986 = ~a7984 & ~a7982;
assign a7988 = ~a7986 & ~l1054;
assign a7990 = ~a7988 & ~a7980;
assign a7992 = a7990 & l1086;
assign a7994 = ~a7978 & ~l1086;
assign a7996 = ~a7994 & ~a7992;
assign a7998 = a7996 & ~a6286;
assign a8000 = ~a7986 & l1086;
assign a8002 = ~a7990 & ~l1086;
assign a8004 = ~a8002 & ~a8000;
assign a8006 = ~a8004 & a6286;
assign a8008 = ~a8006 & ~a7998;
assign a8010 = a8008 & l1088;
assign a8012 = ~a7996 & ~l1088;
assign a8014 = ~a8012 & ~a8010;
assign a8016 = a8014 & ~a6278;
assign a8018 = ~a8004 & l1088;
assign a8020 = ~a8008 & ~l1088;
assign a8022 = ~a8020 & ~a8018;
assign a8024 = ~a8022 & a6278;
assign a8026 = ~a8024 & ~a8016;
assign a8028 = a8026 & l1090;
assign a8030 = ~a8014 & ~l1090;
assign a8032 = ~a8030 & ~a8028;
assign a8034 = a8032 & ~a6270;
assign a8036 = ~a8022 & l1090;
assign a8038 = ~a8026 & ~l1090;
assign a8040 = ~a8038 & ~a8036;
assign a8042 = ~a8040 & a6270;
assign a8044 = ~a8042 & ~a8034;
assign a8046 = a8044 & l1092;
assign a8048 = ~a8032 & ~l1092;
assign a8050 = ~a8048 & ~a8046;
assign a8052 = a8050 & ~a6262;
assign a8054 = ~a8040 & l1092;
assign a8056 = ~a8044 & ~l1092;
assign a8058 = ~a8056 & ~a8054;
assign a8060 = ~a8058 & a6262;
assign a8062 = ~a8060 & ~a8052;
assign a8064 = a8062 & l1024;
assign a8066 = ~a8050 & ~l1024;
assign a8068 = ~a8066 & ~a8064;
assign a8070 = a8068 & ~a6254;
assign a8072 = ~a8058 & l1024;
assign a8074 = ~a8062 & ~l1024;
assign a8076 = ~a8074 & ~a8072;
assign a8078 = ~a8076 & a6254;
assign a8080 = ~a8078 & ~a8070;
assign a8082 = a8080 & l972;
assign a8084 = ~a8068 & ~l972;
assign a8086 = ~a8084 & ~a8082;
assign a8088 = ~a8086 & l886;
assign a8090 = ~a8088 & ~a7876;
assign a8092 = ~a8090 & l970;
assign a8094 = ~a8092 & ~a6418;
assign a8096 = ~a8094 & ~l968;
assign a8098 = ~a8090 & l968;
assign a8100 = ~a8098 & ~a8096;
assign a8102 = ~a8100 & ~l966;
assign a8104 = ~a8090 & l966;
assign a8106 = ~a8104 & ~a8102;
assign a8108 = ~a8106 & ~l964;
assign a8110 = ~a8090 & l964;
assign a8112 = ~a8110 & ~a8108;
assign a8114 = ~a8112 & ~l962;
assign a8116 = ~a8090 & l962;
assign a8118 = ~a8116 & ~a8114;
assign a8120 = ~a8118 & ~l960;
assign a8122 = ~a8090 & l960;
assign a8124 = ~a8122 & ~a8120;
assign a8126 = ~a8124 & ~a5606;
assign a8128 = ~a8090 & a5606;
assign a8130 = ~a8128 & ~a8126;
assign a8132 = ~a8130 & ~a5600;
assign a8134 = ~a8090 & a5600;
assign a8136 = ~a8134 & ~a8132;
assign a8138 = ~a8136 & ~a5594;
assign a8140 = ~a8090 & a5594;
assign a8142 = ~a8140 & ~a8138;
assign a8144 = ~a8142 & ~a5568;
assign a8146 = ~a8090 & a5568;
assign a8148 = ~a8146 & ~a8144;
assign a8152 = a8150 & a8148;
assign a8154 = a6702 & l1060;
assign a8156 = ~a8154 & l1060;
assign a8158 = a8156 & l1082;
assign a8160 = ~a6702 & ~l1060;
assign a8162 = a8160 & ~l1082;
assign a8164 = ~a8162 & ~a8158;
assign a8166 = ~a8164 & l1138;
assign a8168 = ~a8160 & l1082;
assign a8170 = ~a8156 & ~l1082;
assign a8172 = ~a8170 & ~a8168;
assign a8174 = a8172 & l1084;
assign a8176 = ~a8164 & ~l1084;
assign a8178 = ~a8176 & ~a8174;
assign a8180 = ~a8178 & ~l1138;
assign a8182 = ~a8180 & ~a8166;
assign a8184 = ~a8182 & l1130;
assign a8186 = a8178 & l1138;
assign a8188 = ~a8172 & ~l1138;
assign a8190 = ~a8188 & ~a8186;
assign a8192 = a8190 & l1086;
assign a8194 = ~a8182 & ~l1086;
assign a8196 = ~a8194 & ~a8192;
assign a8198 = ~a8196 & ~l1130;
assign a8200 = ~a8198 & ~a8184;
assign a8202 = ~a8200 & ~a6450;
assign a8204 = a8196 & l1130;
assign a8206 = ~a8190 & ~l1130;
assign a8208 = ~a8206 & ~a8204;
assign a8210 = a8208 & l1088;
assign a8212 = ~a8200 & ~l1088;
assign a8214 = ~a8212 & ~a8210;
assign a8216 = ~a8214 & a6450;
assign a8218 = ~a8216 & ~a8202;
assign a8220 = ~a8218 & ~a6442;
assign a8222 = a8214 & ~a6450;
assign a8224 = ~a8208 & a6450;
assign a8226 = ~a8224 & ~a8222;
assign a8228 = a8226 & l1090;
assign a8230 = ~a8218 & ~l1090;
assign a8232 = ~a8230 & ~a8228;
assign a8234 = ~a8232 & a6442;
assign a8236 = ~a8234 & ~a8220;
assign a8238 = ~a8236 & ~a6434;
assign a8240 = a8232 & ~a6442;
assign a8242 = ~a8226 & a6442;
assign a8244 = ~a8242 & ~a8240;
assign a8246 = a8244 & l1092;
assign a8248 = ~a8236 & ~l1092;
assign a8250 = ~a8248 & ~a8246;
assign a8252 = ~a8250 & a6434;
assign a8254 = ~a8252 & ~a8238;
assign a8256 = a8254 & ~a6426;
assign a8258 = a8250 & ~a6434;
assign a8260 = ~a8244 & a6434;
assign a8262 = ~a8260 & ~a8258;
assign a8264 = ~a8262 & a6426;
assign a8266 = ~a8264 & ~a8256;
assign a8268 = a8266 & l1024;
assign a8270 = ~a8254 & ~l1024;
assign a8272 = ~a8270 & ~a8268;
assign a8274 = ~a8272 & l972;
assign a8276 = ~a8254 & l1024;
assign a8278 = ~a8236 & l1092;
assign a8280 = ~a8218 & l1090;
assign a8282 = ~a8200 & l1088;
assign a8284 = ~a8182 & l1086;
assign a8286 = a8164 & l1084;
assign a8288 = ~a8172 & ~l1084;
assign a8290 = ~a8288 & ~a8286;
assign a8292 = a8290 & l1138;
assign a8294 = ~a8164 & ~l1138;
assign a8296 = ~a8294 & ~a8292;
assign a8298 = ~a8296 & ~l1086;
assign a8300 = ~a8298 & ~a8284;
assign a8302 = ~a8300 & l1130;
assign a8304 = ~a8182 & ~l1130;
assign a8306 = ~a8304 & ~a8302;
assign a8308 = ~a8306 & ~l1088;
assign a8310 = ~a8308 & ~a8282;
assign a8312 = ~a8310 & ~a6450;
assign a8314 = ~a8200 & a6450;
assign a8316 = ~a8314 & ~a8312;
assign a8318 = ~a8316 & ~l1090;
assign a8320 = ~a8318 & ~a8280;
assign a8322 = ~a8320 & ~a6442;
assign a8324 = ~a8218 & a6442;
assign a8326 = ~a8324 & ~a8322;
assign a8328 = ~a8326 & ~l1092;
assign a8330 = ~a8328 & ~a8278;
assign a8332 = ~a8330 & ~a6434;
assign a8334 = ~a8236 & a6434;
assign a8336 = ~a8334 & ~a8332;
assign a8338 = ~a8336 & ~a6426;
assign a8340 = ~a8254 & a6426;
assign a8342 = ~a8340 & ~a8338;
assign a8344 = ~a8342 & ~l1024;
assign a8346 = ~a8344 & ~a8276;
assign a8348 = ~a8346 & ~a7226;
assign a8350 = ~a8272 & a7226;
assign a8352 = ~a8350 & ~a8348;
assign a8354 = ~a8352 & ~l972;
assign a8356 = ~a8354 & ~a8274;
assign a8358 = ~a8356 & l948;
assign a8360 = ~a8358 & ~a7872;
assign a8362 = ~a8360 & ~l886;
assign a8364 = ~a8362 & ~a8088;
assign a8366 = ~a8364 & l970;
assign a8368 = ~a8366 & ~a6418;
assign a8370 = ~a8368 & ~l968;
assign a8372 = ~a8364 & l968;
assign a8374 = ~a8372 & ~a8370;
assign a8376 = ~a8374 & ~l966;
assign a8378 = ~a8364 & l966;
assign a8380 = ~a8378 & ~a8376;
assign a8382 = ~a8380 & ~l964;
assign a8384 = ~a8364 & l964;
assign a8386 = ~a8384 & ~a8382;
assign a8388 = ~a8386 & ~l962;
assign a8390 = ~a8364 & l962;
assign a8392 = ~a8390 & ~a8388;
assign a8394 = ~a8392 & ~l960;
assign a8396 = ~a8364 & l960;
assign a8398 = ~a8396 & ~a8394;
assign a8400 = ~a8398 & ~a5606;
assign a8402 = ~a8364 & a5606;
assign a8404 = ~a8402 & ~a8400;
assign a8406 = ~a8404 & ~a5600;
assign a8408 = ~a8364 & a5600;
assign a8410 = ~a8408 & ~a8406;
assign a8412 = ~a8410 & ~a5594;
assign a8414 = ~a8364 & a5594;
assign a8416 = ~a8414 & ~a8412;
assign a8418 = ~a8416 & ~a5568;
assign a8420 = ~a8364 & a5568;
assign a8422 = ~a8420 & ~a8418;
assign a8424 = a8422 & a8150;
assign a8426 = ~a8424 & ~a8152;
assign a8428 = a8426 & i326;
assign a8430 = ~a8428 & ~a8152;
assign a8432 = a8430 & l930;
assign a8434 = a8430 & a8150;
assign a8436 = ~a6506 & l1220;
assign a8438 = ~a6512 & ~l1220;
assign a8440 = ~a8438 & ~a8436;
assign a8442 = ~a8440 & l1204;
assign a8444 = ~a6522 & l1220;
assign a8446 = ~a6528 & ~l1220;
assign a8448 = ~a8446 & ~a8444;
assign a8450 = ~a8448 & ~l1236;
assign a8452 = a6512 & l1220;
assign a8454 = a6538 & ~l1220;
assign a8456 = ~a8454 & ~a8452;
assign a8458 = a8456 & l1236;
assign a8460 = ~a8458 & ~a8450;
assign a8462 = ~a8460 & ~l1204;
assign a8464 = ~a8462 & ~a8442;
assign a8466 = ~a8464 & ~l1148;
assign a8468 = ~a8466 & ~l1148;
assign a8470 = ~a8468 & l1180;
assign a8472 = ~a6560 & l1220;
assign a8474 = ~a6566 & ~l1220;
assign a8476 = ~a8474 & ~a8472;
assign a8478 = ~a8476 & l1236;
assign a8480 = ~a8478 & ~a8450;
assign a8482 = a8480 & l1204;
assign a8484 = ~a6580 & l1220;
assign a8486 = ~a6506 & ~l1220;
assign a8488 = ~a8486 & ~a8484;
assign a8490 = a8488 & l1236;
assign a8492 = ~a8456 & ~l1236;
assign a8494 = ~a8492 & ~a8490;
assign a8496 = ~a8494 & ~l1204;
assign a8498 = ~a8496 & ~a8482;
assign a8500 = a8498 & l1148;
assign a8502 = ~a8500 & l1148;
assign a8504 = ~a8502 & ~l1180;
assign a8506 = ~a8504 & ~a8470;
assign a8508 = ~a8506 & ~l1172;
assign a8510 = ~a8508 & ~a6606;
assign a8512 = ~a8510 & ~l928;
assign a8514 = ~a8512 & ~a6694;
assign a8516 = ~a8514 & l930;
assign a8518 = ~a8516 & ~a6706;
assign a8520 = ~a8518 & l900;
assign a8522 = ~a8520 & ~a6704;
assign a8524 = a8522 & l1060;
assign a8526 = ~a8524 & l1060;
assign a8528 = a8526 & l1082;
assign a8530 = ~a8522 & ~l1060;
assign a8532 = a8530 & ~l1082;
assign a8534 = ~a8532 & ~a8528;
assign a8536 = ~a8534 & l1138;
assign a8538 = ~a8530 & l1082;
assign a8540 = ~a8526 & ~l1082;
assign a8542 = ~a8540 & ~a8538;
assign a8544 = a8542 & l1084;
assign a8546 = ~a8534 & ~l1084;
assign a8548 = ~a8546 & ~a8544;
assign a8550 = ~a8548 & ~l1138;
assign a8552 = ~a8550 & ~a8536;
assign a8554 = ~a8552 & l1130;
assign a8556 = a8548 & l1138;
assign a8558 = ~a8542 & ~l1138;
assign a8560 = ~a8558 & ~a8556;
assign a8562 = a8560 & l1086;
assign a8564 = ~a8552 & ~l1086;
assign a8566 = ~a8564 & ~a8562;
assign a8568 = ~a8566 & ~l1130;
assign a8570 = ~a8568 & ~a8554;
assign a8572 = ~a8570 & ~a6450;
assign a8574 = a8566 & l1130;
assign a8576 = ~a8560 & ~l1130;
assign a8578 = ~a8576 & ~a8574;
assign a8580 = a8578 & l1088;
assign a8582 = ~a8570 & ~l1088;
assign a8584 = ~a8582 & ~a8580;
assign a8586 = ~a8584 & a6450;
assign a8588 = ~a8586 & ~a8572;
assign a8590 = ~a8588 & ~a6442;
assign a8592 = a8584 & ~a6450;
assign a8594 = ~a8578 & a6450;
assign a8596 = ~a8594 & ~a8592;
assign a8598 = a8596 & l1090;
assign a8600 = ~a8588 & ~l1090;
assign a8602 = ~a8600 & ~a8598;
assign a8604 = ~a8602 & a6442;
assign a8606 = ~a8604 & ~a8590;
assign a8608 = ~a8606 & ~a6434;
assign a8610 = a8602 & ~a6442;
assign a8612 = ~a8596 & a6442;
assign a8614 = ~a8612 & ~a8610;
assign a8616 = a8614 & l1092;
assign a8618 = ~a8606 & ~l1092;
assign a8620 = ~a8618 & ~a8616;
assign a8622 = ~a8620 & a6434;
assign a8624 = ~a8622 & ~a8608;
assign a8626 = a8624 & ~a6426;
assign a8628 = a8620 & ~a6434;
assign a8630 = ~a8614 & a6434;
assign a8632 = ~a8630 & ~a8628;
assign a8634 = ~a8632 & a6426;
assign a8636 = ~a8634 & ~a8626;
assign a8638 = a8636 & l1024;
assign a8640 = ~a8624 & ~l1024;
assign a8642 = ~a8640 & ~a8638;
assign a8644 = ~a8642 & l972;
assign a8646 = ~a8624 & l1024;
assign a8648 = ~a8606 & l1092;
assign a8650 = ~a8588 & l1090;
assign a8652 = ~a8570 & l1088;
assign a8654 = ~a8552 & l1086;
assign a8656 = a8534 & l1084;
assign a8658 = ~a8542 & ~l1084;
assign a8660 = ~a8658 & ~a8656;
assign a8662 = a8660 & l1138;
assign a8664 = ~a8534 & ~l1138;
assign a8666 = ~a8664 & ~a8662;
assign a8668 = ~a8666 & ~l1086;
assign a8670 = ~a8668 & ~a8654;
assign a8672 = ~a8670 & l1130;
assign a8674 = ~a8552 & ~l1130;
assign a8676 = ~a8674 & ~a8672;
assign a8678 = ~a8676 & ~l1088;
assign a8680 = ~a8678 & ~a8652;
assign a8682 = ~a8680 & ~a6450;
assign a8684 = ~a8570 & a6450;
assign a8686 = ~a8684 & ~a8682;
assign a8688 = ~a8686 & ~l1090;
assign a8690 = ~a8688 & ~a8650;
assign a8692 = ~a8690 & ~a6442;
assign a8694 = ~a8588 & a6442;
assign a8696 = ~a8694 & ~a8692;
assign a8698 = ~a8696 & ~l1092;
assign a8700 = ~a8698 & ~a8648;
assign a8702 = ~a8700 & ~a6434;
assign a8704 = ~a8606 & a6434;
assign a8706 = ~a8704 & ~a8702;
assign a8708 = ~a8706 & ~a6426;
assign a8710 = ~a8624 & a6426;
assign a8712 = ~a8710 & ~a8708;
assign a8714 = ~a8712 & ~l1024;
assign a8716 = ~a8714 & ~a8646;
assign a8718 = ~a8716 & ~a7226;
assign a8720 = ~a8642 & a7226;
assign a8722 = ~a8720 & ~a8718;
assign a8724 = ~a8722 & ~l972;
assign a8726 = ~a8724 & ~a8644;
assign a8728 = ~a8726 & l948;
assign a8730 = ~a8728 & ~a7872;
assign a8732 = ~a8730 & ~l886;
assign a8734 = ~a8732 & ~a8088;
assign a8736 = ~a8734 & l970;
assign a8738 = ~a8736 & ~a6418;
assign a8740 = ~a8738 & ~l968;
assign a8742 = ~a8734 & l968;
assign a8744 = ~a8742 & ~a8740;
assign a8746 = ~a8744 & ~l966;
assign a8748 = ~a8734 & l966;
assign a8750 = ~a8748 & ~a8746;
assign a8752 = ~a8750 & ~l964;
assign a8754 = ~a8734 & l964;
assign a8756 = ~a8754 & ~a8752;
assign a8758 = ~a8756 & ~l962;
assign a8760 = ~a8734 & l962;
assign a8762 = ~a8760 & ~a8758;
assign a8764 = ~a8762 & ~l960;
assign a8766 = ~a8734 & l960;
assign a8768 = ~a8766 & ~a8764;
assign a8770 = ~a8768 & ~a5606;
assign a8772 = ~a8734 & a5606;
assign a8774 = ~a8772 & ~a8770;
assign a8776 = ~a8774 & ~a5600;
assign a8778 = ~a8734 & a5600;
assign a8780 = ~a8778 & ~a8776;
assign a8782 = ~a8780 & ~a5594;
assign a8784 = ~a8734 & a5594;
assign a8786 = ~a8784 & ~a8782;
assign a8788 = ~a8786 & ~a5568;
assign a8790 = ~a8734 & a5568;
assign a8792 = ~a8790 & ~a8788;
assign a8794 = a8792 & a8434;
assign a8796 = a8434 & a8422;
assign a8798 = ~a8796 & ~a8794;
assign a8800 = a8798 & i328;
assign a8802 = ~a8800 & ~a8794;
assign a8804 = a8802 & a8432;
assign a8806 = a8804 & l900;
assign a8808 = ~a8806 & ~a5628;
assign a8810 = l1172 & l896;
assign a8812 = ~a8810 & a8808;
assign a8816 = a8814 & l1218;
assign a8818 = ~a8814 & ~l1172;
assign a8820 = a8818 & l1220;
assign a8822 = ~a8820 & ~a8816;
assign a8824 = l1216 & l1172;
assign a8826 = ~a8824 & a8822;
assign a8828 = a8814 & l1178;
assign a8830 = a8818 & l1180;
assign a8832 = ~a8830 & ~a8828;
assign a8834 = l1176 & l1172;
assign a8836 = ~a8834 & a8832;
assign a8838 = a8814 & l1202;
assign a8840 = a8818 & l1204;
assign a8842 = ~a8840 & ~a8838;
assign a8844 = l1200 & l1172;
assign a8846 = ~a8844 & a8842;
assign a8848 = ~a8846 & ~a8836;
assign a8850 = a8848 & ~a8826;
assign a8852 = a8814 & l1234;
assign a8854 = a8818 & l1236;
assign a8856 = ~a8854 & ~a8852;
assign a8858 = l1232 & l1172;
assign a8860 = ~a8858 & a8856;
assign a8862 = ~a8860 & a8836;
assign a8864 = ~a8862 & ~a8850;
assign a8866 = ~a8864 & ~a8812;
assign a8868 = a8812 & l1170;
assign a8870 = ~a8868 & ~a8866;
assign a8872 = ~a8870 & l948;
assign a8874 = ~a5748 & ~l948;
assign a8876 = a8874 & l1246;
assign a8878 = a7322 & ~a7316;
assign a8880 = a8878 & l1246;
assign a8882 = a8880 & a7328;
assign a8884 = ~a8882 & ~a8874;
assign a8886 = ~a7322 & ~a7316;
assign a8888 = a8886 & ~a7328;
assign a8890 = ~a8888 & l1246;
assign a8892 = a8888 & ~l1246;
assign a8894 = ~a8892 & ~a8890;
assign a8896 = ~a8894 & a8884;
assign a8898 = ~a8896 & ~a8876;
assign a8900 = ~a8898 & ~l948;
assign a8902 = ~a8900 & ~a8872;
assign a8904 = ~a8902 & ~l886;
assign a8906 = ~a8904 & ~a5626;
assign a8908 = ~a2532 & l886;
assign a8910 = a8836 & ~a8826;
assign a8912 = a8848 & a8826;
assign a8914 = ~a8912 & ~a8910;
assign a8916 = a8846 & ~a8826;
assign a8918 = ~a8916 & a8914;
assign a8920 = ~a8918 & ~a8812;
assign a8922 = a8812 & l1168;
assign a8924 = ~a8922 & ~a8920;
assign a8926 = ~a8924 & l948;
assign a8928 = a8874 & ~a7328;
assign a8930 = ~a8886 & ~a7328;
assign a8932 = a8886 & a7328;
assign a8934 = ~a8932 & ~a8930;
assign a8936 = ~a8934 & ~a8874;
assign a8938 = ~a8936 & ~a8928;
assign a8940 = ~a8938 & ~l948;
assign a8942 = ~a8940 & ~a8926;
assign a8944 = ~a8942 & ~l886;
assign a8948 = l886 & ~l880;
assign a8950 = a8836 & ~a8812;
assign a8952 = a8812 & l1146;
assign a8954 = ~a8952 & ~a8950;
assign a8956 = ~a8954 & l948;
assign a8958 = a8874 & ~a7316;
assign a8960 = ~a8874 & a7316;
assign a8962 = ~a8960 & ~a8958;
assign a8964 = ~a8962 & ~l948;
assign a8966 = ~a8964 & ~a8956;
assign a8968 = ~a8966 & ~l886;
assign a8972 = ~a2748 & l886;
assign a8974 = a8846 & ~a8836;
assign a8976 = a8974 & a8860;
assign a8978 = ~a8846 & a8836;
assign a8980 = ~a8978 & ~a8976;
assign a8982 = ~a8980 & ~a8812;
assign a8984 = a8812 & l1160;
assign a8986 = ~a8984 & ~a8982;
assign a8988 = ~a8986 & l948;
assign a8990 = a8874 & ~a7322;
assign a8992 = ~a7322 & a7316;
assign a8994 = ~a8992 & ~a8878;
assign a8996 = ~a8994 & a8884;
assign a8998 = ~a8996 & ~a8990;
assign a9000 = ~a8998 & ~l948;
assign a9002 = ~a9000 & ~a8988;
assign a9004 = ~a9002 & ~l886;
assign a9008 = a9006 & a8970;
assign a9010 = a9008 & a8946;
assign a9012 = a9010 & a8906;
assign a9014 = ~a9012 & ~a5624;
assign a9016 = ~a9010 & ~a8906;
assign a9018 = ~a9016 & ~a9012;
assign a9020 = ~a9018 & a9014;
assign a9022 = a8906 & a5624;
assign a9024 = ~a9022 & ~a9014;
assign a9026 = ~a9024 & ~a9020;
assign a9028 = ~a8870 & l1196;
assign a9030 = ~l916 & l890;
assign a9032 = a5178 & i156;
assign a9034 = a9032 & ~a5370;
assign a9036 = ~a9034 & ~l890;
assign a9038 = ~a9036 & ~a9030;
assign a9040 = ~l1192 & l890;
assign a9042 = ~a9034 & ~l890;
assign a9044 = ~a9042 & ~a9040;
assign a9046 = ~a9044 & ~a9038;
assign a9048 = a9046 & l1250;
assign a9050 = a9048 & l1274;
assign a9052 = a9044 & a9038;
assign a9054 = ~l1256 & l890;
assign a9056 = ~a9034 & ~l890;
assign a9058 = ~a9056 & ~a9054;
assign a9060 = a9058 & a9052;
assign a9062 = a9060 & l1274;
assign a9064 = ~l912 & ~l908;
assign a9066 = ~a9064 & l1276;
assign a9068 = ~l1284 & l890;
assign a9070 = ~a4832 & ~l890;
assign a9072 = ~a9070 & ~a9068;
assign a9074 = ~l1132 & l890;
assign a9076 = a2560 & i2;
assign a9078 = a5178 & a3976;
assign a9080 = a9078 & a4166;
assign a9082 = ~a9078 & ~a4166;
assign a9084 = ~a9082 & ~a9080;
assign a9086 = a5178 & a4980;
assign a9088 = ~a9086 & ~a4278;
assign a9090 = a9086 & a4278;
assign a9092 = ~a9090 & ~a9088;
assign a9094 = ~a9092 & ~a9080;
assign a9096 = a9092 & a9080;
assign a9098 = ~a9096 & ~a9094;
assign a9100 = ~a9090 & ~a9080;
assign a9102 = ~a9100 & ~a9088;
assign a9104 = a5178 & a5028;
assign a9106 = ~a9104 & ~a4430;
assign a9108 = a9104 & a4430;
assign a9110 = ~a9108 & ~a9106;
assign a9112 = ~a9110 & ~a9102;
assign a9114 = a9110 & a9102;
assign a9116 = ~a9114 & ~a9112;
assign a9118 = ~a9108 & ~a9102;
assign a9120 = ~a9118 & ~a9106;
assign a9122 = a5178 & a5076;
assign a9124 = ~a9122 & ~a4590;
assign a9126 = a9122 & a4590;
assign a9128 = ~a9126 & ~a9124;
assign a9130 = ~a9128 & ~a9120;
assign a9132 = a9128 & a9120;
assign a9134 = ~a9132 & ~a9130;
assign a9136 = ~a9126 & ~a9120;
assign a9138 = ~a9136 & ~a9124;
assign a9140 = a5178 & a5124;
assign a9142 = ~a9140 & ~a4750;
assign a9144 = a9140 & a4750;
assign a9146 = ~a9144 & ~a9142;
assign a9148 = ~a9146 & ~a9138;
assign a9150 = a9146 & a9138;
assign a9152 = ~a9150 & ~a9148;
assign a9154 = ~a9144 & ~a9138;
assign a9156 = ~a9154 & ~a9142;
assign a9158 = ~a9156 & ~a4888;
assign a9160 = ~a9158 & a9152;
assign a9162 = a9160 & a9134;
assign a9164 = a9162 & a9116;
assign a9166 = a9164 & a9098;
assign a9168 = a9166 & a9084;
assign a9170 = i262 & i260;
assign a9172 = a9170 & i258;
assign a9174 = a9172 & i256;
assign a9176 = a9174 & i254;
assign a9178 = ~i266 & ~i264;
assign a9180 = ~a9178 & a9176;
assign a9182 = ~a9180 & ~i268;
assign a9184 = i274 & i268;
assign a9186 = a9184 & i272;
assign a9188 = ~a9186 & i270;
assign a9190 = a9186 & ~i270;
assign a9192 = ~a9190 & ~a9188;
assign a9194 = ~a9192 & ~a9180;
assign a9196 = ~a9194 & ~a9084;
assign a9198 = a9186 & i270;
assign a9200 = ~a9198 & i266;
assign a9202 = ~a9200 & ~a9180;
assign a9204 = a9198 & ~i266;
assign a9206 = ~a9204 & a9202;
assign a9208 = a9206 & ~a9084;
assign a9210 = a9198 & i266;
assign a9212 = ~a9210 & i264;
assign a9214 = a9210 & ~i264;
assign a9216 = ~a9214 & ~a9212;
assign a9218 = ~a9216 & ~a9180;
assign a9220 = ~a9218 & ~a9084;
assign a9222 = a9210 & i264;
assign a9224 = ~a9222 & i260;
assign a9226 = ~a9224 & ~a9180;
assign a9228 = a9222 & ~i260;
assign a9230 = ~a9228 & a9226;
assign a9232 = ~a9158 & ~a9084;
assign a9234 = a9230 & ~a9084;
assign a9236 = a9222 & i260;
assign a9238 = ~a9236 & i262;
assign a9240 = ~a9238 & ~a9180;
assign a9242 = a9236 & ~i262;
assign a9244 = ~a9242 & a9240;
assign a9246 = a9232 & a9152;
assign a9248 = a9244 & ~a9084;
assign a9250 = a9236 & i262;
assign a9252 = ~a9250 & i258;
assign a9254 = ~a9252 & ~a9180;
assign a9256 = a9250 & ~i258;
assign a9258 = ~a9256 & a9254;
assign a9260 = a9246 & a9134;
assign a9262 = a9258 & ~a9084;
assign a9264 = a9250 & i258;
assign a9266 = ~a9264 & i256;
assign a9268 = ~a9266 & ~a9180;
assign a9270 = a9264 & ~i256;
assign a9272 = ~a9270 & a9268;
assign a9274 = a9260 & a9116;
assign a9276 = a9272 & ~a9084;
assign a9278 = a9264 & i256;
assign a9280 = a9278 & ~i254;
assign a9282 = ~a9280 & ~i254;
assign a9284 = a9274 & a9098;
assign a9286 = a9282 & ~a9084;
assign a9288 = ~a9286 & a9284;
assign a9290 = ~a9288 & ~a9282;
assign a9292 = ~a9290 & ~a9098;
assign a9294 = ~a9292 & ~a9276;
assign a9296 = a9290 & a9098;
assign a9298 = ~a9296 & ~a9294;
assign a9300 = ~a9298 & a9274;
assign a9302 = ~a9300 & ~a9272;
assign a9304 = ~a9302 & ~a9098;
assign a9306 = ~a9304 & ~a9262;
assign a9308 = a9302 & a9098;
assign a9310 = ~a9308 & ~a9306;
assign a9312 = ~a9158 & ~a9098;
assign a9314 = a9312 & a9152;
assign a9316 = a9314 & a9134;
assign a9318 = a9316 & a9116;
assign a9320 = a9318 & ~a9298;
assign a9322 = ~a9320 & a9290;
assign a9324 = ~a9322 & ~a9116;
assign a9326 = ~a9324 & ~a9310;
assign a9328 = a9322 & a9116;
assign a9330 = ~a9328 & ~a9326;
assign a9332 = ~a9330 & a9260;
assign a9334 = a9332 & a9258;
assign a9336 = ~a9332 & ~a9258;
assign a9338 = ~a9336 & ~a9334;
assign a9340 = a9338 & ~a9098;
assign a9342 = ~a9340 & ~a9248;
assign a9344 = ~a9338 & a9098;
assign a9346 = ~a9344 & ~a9342;
assign a9348 = ~a9330 & a9316;
assign a9350 = a9348 & ~a9302;
assign a9352 = ~a9348 & a9302;
assign a9354 = ~a9352 & ~a9350;
assign a9356 = ~a9354 & ~a9334;
assign a9358 = ~a9356 & ~a9116;
assign a9360 = ~a9358 & ~a9346;
assign a9362 = a9356 & a9116;
assign a9364 = ~a9362 & ~a9360;
assign a9366 = ~a9350 & a9322;
assign a9368 = ~a9158 & ~a9116;
assign a9370 = a9368 & a9152;
assign a9372 = a9370 & a9134;
assign a9374 = a9372 & ~a9330;
assign a9376 = ~a9374 & a9366;
assign a9378 = ~a9376 & ~a9134;
assign a9380 = ~a9378 & ~a9364;
assign a9382 = a9376 & a9134;
assign a9384 = ~a9382 & ~a9380;
assign a9386 = ~a9384 & a9246;
assign a9388 = ~a9386 & ~a9244;
assign a9390 = a9386 & a9244;
assign a9392 = ~a9390 & ~a9388;
assign a9394 = a9392 & ~a9098;
assign a9396 = ~a9394 & ~a9234;
assign a9398 = ~a9392 & a9098;
assign a9400 = ~a9398 & ~a9396;
assign a9402 = ~a9384 & a9314;
assign a9404 = a9402 & a9338;
assign a9406 = ~a9402 & ~a9338;
assign a9408 = ~a9406 & ~a9404;
assign a9410 = ~a9408 & ~a9390;
assign a9412 = a9408 & a9390;
assign a9414 = ~a9412 & ~a9410;
assign a9416 = a9414 & ~a9116;
assign a9418 = ~a9416 & ~a9400;
assign a9420 = ~a9414 & a9116;
assign a9422 = ~a9420 & ~a9418;
assign a9424 = ~a9384 & a9370;
assign a9426 = a9424 & ~a9356;
assign a9428 = ~a9424 & a9356;
assign a9430 = ~a9428 & ~a9426;
assign a9432 = ~a9404 & ~a9390;
assign a9434 = ~a9432 & ~a9406;
assign a9436 = ~a9434 & ~a9430;
assign a9438 = a9434 & a9430;
assign a9440 = ~a9438 & ~a9436;
assign a9442 = a9440 & ~a9134;
assign a9444 = ~a9442 & ~a9422;
assign a9446 = ~a9440 & a9134;
assign a9448 = ~a9446 & ~a9444;
assign a9450 = ~a9158 & ~a9134;
assign a9452 = a9450 & a9152;
assign a9454 = a9452 & ~a9384;
assign a9456 = ~a9454 & a9376;
assign a9458 = ~a9434 & ~a9426;
assign a9460 = ~a9458 & ~a9428;
assign a9462 = ~a9460 & a9456;
assign a9464 = ~a9462 & ~a9152;
assign a9466 = ~a9464 & ~a9448;
assign a9468 = a9462 & a9152;
assign a9470 = ~a9468 & ~a9466;
assign a9472 = ~a9470 & a9232;
assign a9474 = ~a9472 & ~a9230;
assign a9476 = a9472 & a9230;
assign a9478 = ~a9476 & ~a9474;
assign a9480 = a9478 & ~a9098;
assign a9482 = ~a9480 & ~a9220;
assign a9484 = ~a9478 & a9098;
assign a9486 = ~a9484 & ~a9482;
assign a9488 = ~a9470 & a9312;
assign a9490 = a9488 & a9392;
assign a9492 = ~a9488 & ~a9392;
assign a9494 = ~a9492 & ~a9490;
assign a9496 = ~a9494 & ~a9476;
assign a9498 = a9494 & a9476;
assign a9500 = ~a9498 & ~a9496;
assign a9502 = a9500 & ~a9116;
assign a9504 = ~a9502 & ~a9486;
assign a9506 = ~a9500 & a9116;
assign a9508 = ~a9506 & ~a9504;
assign a9510 = ~a9470 & a9368;
assign a9512 = a9510 & a9414;
assign a9514 = ~a9510 & ~a9414;
assign a9516 = ~a9514 & ~a9512;
assign a9518 = ~a9490 & ~a9476;
assign a9520 = ~a9518 & ~a9492;
assign a9522 = ~a9520 & ~a9516;
assign a9524 = a9520 & a9516;
assign a9526 = ~a9524 & ~a9522;
assign a9528 = a9526 & ~a9134;
assign a9530 = ~a9528 & ~a9508;
assign a9532 = ~a9526 & a9134;
assign a9534 = ~a9532 & ~a9530;
assign a9536 = ~a9470 & a9450;
assign a9538 = a9536 & a9440;
assign a9540 = ~a9536 & ~a9440;
assign a9542 = ~a9540 & ~a9538;
assign a9544 = ~a9520 & ~a9512;
assign a9546 = ~a9544 & ~a9514;
assign a9548 = ~a9546 & ~a9542;
assign a9550 = a9546 & a9542;
assign a9552 = ~a9550 & ~a9548;
assign a9554 = a9552 & ~a9152;
assign a9556 = ~a9554 & ~a9534;
assign a9558 = ~a9552 & a9152;
assign a9560 = ~a9558 & ~a9556;
assign a9562 = ~a9158 & ~a9152;
assign a9564 = a9562 & ~a9470;
assign a9566 = ~a9564 & a9462;
assign a9568 = ~a9546 & ~a9538;
assign a9570 = ~a9568 & ~a9540;
assign a9572 = ~a9570 & a9566;
assign a9574 = ~a9572 & a9158;
assign a9576 = ~a9574 & ~a9560;
assign a9578 = a9572 & ~a9158;
assign a9580 = ~a9578 & ~a9576;
assign a9582 = ~a9580 & ~a9084;
assign a9584 = a9582 & ~a9218;
assign a9586 = ~a9582 & a9218;
assign a9588 = ~a9586 & ~a9584;
assign a9590 = a9588 & ~a9098;
assign a9592 = ~a9590 & ~a9208;
assign a9594 = ~a9588 & a9098;
assign a9596 = ~a9594 & ~a9592;
assign a9598 = ~a9580 & ~a9098;
assign a9600 = a9598 & a9478;
assign a9602 = ~a9598 & ~a9478;
assign a9604 = ~a9602 & ~a9600;
assign a9606 = ~a9604 & ~a9584;
assign a9608 = a9604 & a9584;
assign a9610 = ~a9608 & ~a9606;
assign a9612 = a9610 & ~a9116;
assign a9614 = ~a9612 & ~a9596;
assign a9616 = ~a9610 & a9116;
assign a9618 = ~a9616 & ~a9614;
assign a9620 = ~a9580 & ~a9116;
assign a9622 = a9620 & a9500;
assign a9624 = ~a9620 & ~a9500;
assign a9626 = ~a9624 & ~a9622;
assign a9628 = ~a9600 & ~a9584;
assign a9630 = ~a9628 & ~a9602;
assign a9632 = ~a9630 & ~a9626;
assign a9634 = a9630 & a9626;
assign a9636 = ~a9634 & ~a9632;
assign a9638 = a9636 & ~a9134;
assign a9640 = ~a9638 & ~a9618;
assign a9642 = ~a9636 & a9134;
assign a9644 = ~a9642 & ~a9640;
assign a9646 = ~a9580 & ~a9134;
assign a9648 = a9646 & a9526;
assign a9650 = ~a9646 & ~a9526;
assign a9652 = ~a9650 & ~a9648;
assign a9654 = ~a9630 & ~a9622;
assign a9656 = ~a9654 & ~a9624;
assign a9658 = ~a9656 & ~a9652;
assign a9660 = a9656 & a9652;
assign a9662 = ~a9660 & ~a9658;
assign a9664 = a9662 & ~a9152;
assign a9666 = ~a9664 & ~a9644;
assign a9668 = ~a9662 & a9152;
assign a9670 = ~a9668 & ~a9666;
assign a9672 = ~a9580 & ~a9152;
assign a9674 = a9672 & a9552;
assign a9676 = ~a9672 & ~a9552;
assign a9678 = ~a9676 & ~a9674;
assign a9680 = ~a9656 & ~a9648;
assign a9682 = ~a9680 & ~a9650;
assign a9684 = ~a9682 & ~a9678;
assign a9686 = a9682 & a9678;
assign a9688 = ~a9686 & ~a9684;
assign a9690 = a9688 & a9158;
assign a9692 = ~a9690 & ~a9670;
assign a9694 = ~a9688 & ~a9158;
assign a9696 = ~a9694 & ~a9692;
assign a9698 = ~a9580 & a9158;
assign a9700 = ~a9698 & a9572;
assign a9702 = ~a9682 & ~a9674;
assign a9704 = ~a9702 & ~a9676;
assign a9706 = ~a9704 & a9700;
assign a9708 = ~a9706 & a9696;
assign a9710 = ~a9708 & ~a9084;
assign a9712 = a9710 & a9206;
assign a9714 = ~a9710 & ~a9206;
assign a9716 = ~a9714 & ~a9712;
assign a9718 = a9716 & ~a9098;
assign a9720 = ~a9718 & ~a9196;
assign a9722 = ~a9716 & a9098;
assign a9724 = ~a9722 & ~a9720;
assign a9726 = ~a9708 & ~a9098;
assign a9728 = ~a9726 & ~a9588;
assign a9730 = a9726 & a9588;
assign a9732 = ~a9730 & ~a9728;
assign a9734 = ~a9732 & ~a9712;
assign a9736 = a9732 & a9712;
assign a9738 = ~a9736 & ~a9734;
assign a9740 = a9738 & ~a9116;
assign a9742 = ~a9740 & ~a9724;
assign a9744 = ~a9738 & a9116;
assign a9746 = ~a9744 & ~a9742;
assign a9748 = ~a9708 & ~a9116;
assign a9750 = a9748 & a9610;
assign a9752 = ~a9748 & ~a9610;
assign a9754 = ~a9752 & ~a9750;
assign a9756 = ~a9730 & ~a9712;
assign a9758 = ~a9756 & ~a9728;
assign a9760 = ~a9758 & ~a9754;
assign a9762 = a9758 & a9754;
assign a9764 = ~a9762 & ~a9760;
assign a9766 = a9764 & ~a9134;
assign a9768 = ~a9766 & ~a9746;
assign a9770 = ~a9764 & a9134;
assign a9772 = ~a9770 & ~a9768;
assign a9774 = ~a9708 & ~a9134;
assign a9776 = a9774 & a9636;
assign a9778 = ~a9774 & ~a9636;
assign a9780 = ~a9778 & ~a9776;
assign a9782 = ~a9758 & ~a9750;
assign a9784 = ~a9782 & ~a9752;
assign a9786 = ~a9784 & ~a9780;
assign a9788 = a9784 & a9780;
assign a9790 = ~a9788 & ~a9786;
assign a9792 = a9790 & ~a9152;
assign a9794 = ~a9792 & ~a9772;
assign a9796 = ~a9790 & a9152;
assign a9798 = ~a9796 & ~a9794;
assign a9800 = ~a9708 & ~a9152;
assign a9802 = a9800 & a9662;
assign a9804 = ~a9800 & ~a9662;
assign a9806 = ~a9804 & ~a9802;
assign a9808 = ~a9784 & ~a9776;
assign a9810 = ~a9808 & ~a9778;
assign a9812 = ~a9810 & ~a9806;
assign a9814 = a9810 & a9806;
assign a9816 = ~a9814 & ~a9812;
assign a9818 = a9816 & a9158;
assign a9820 = ~a9818 & ~a9798;
assign a9822 = ~a9816 & ~a9158;
assign a9824 = ~a9822 & ~a9820;
assign a9826 = ~a9708 & a9158;
assign a9828 = a9826 & a9688;
assign a9830 = ~a9826 & ~a9688;
assign a9832 = ~a9830 & ~a9828;
assign a9834 = ~a9810 & ~a9802;
assign a9836 = ~a9834 & ~a9804;
assign a9838 = ~a9836 & ~a9832;
assign a9840 = a9836 & a9832;
assign a9842 = ~a9840 & ~a9838;
assign a9844 = a9842 & a9824;
assign a9846 = ~a9844 & ~a9084;
assign a9848 = a9846 & ~a9194;
assign a9850 = ~a9844 & ~a9098;
assign a9852 = ~a9850 & ~a9716;
assign a9854 = a9850 & a9716;
assign a9856 = ~a9854 & ~a9852;
assign a9858 = ~a9856 & ~a9848;
assign a9860 = a9856 & a9848;
assign a9862 = ~a9860 & ~a9858;
assign a9864 = ~a9184 & i272;
assign a9866 = a9184 & ~i272;
assign a9868 = ~a9866 & ~a9864;
assign a9870 = ~a9868 & ~a9180;
assign a9872 = ~a9870 & ~a9084;
assign a9874 = ~a9846 & a9194;
assign a9876 = ~a9874 & ~a9848;
assign a9878 = a9876 & ~a9098;
assign a9880 = ~a9878 & ~a9872;
assign a9882 = ~a9876 & a9098;
assign a9884 = ~a9882 & ~a9880;
assign a9886 = a9862 & ~a9116;
assign a9888 = ~a9886 & ~a9884;
assign a9890 = ~a9862 & a9116;
assign a9892 = ~a9890 & ~a9888;
assign a9894 = ~a9854 & ~a9848;
assign a9896 = ~a9894 & ~a9852;
assign a9898 = ~a9844 & ~a9116;
assign a9900 = ~a9898 & ~a9738;
assign a9902 = a9898 & a9738;
assign a9904 = ~a9902 & ~a9900;
assign a9906 = ~a9904 & ~a9896;
assign a9908 = a9904 & a9896;
assign a9910 = ~a9908 & ~a9906;
assign a9912 = a9910 & ~a9134;
assign a9914 = ~a9912 & ~a9892;
assign a9916 = ~a9910 & a9134;
assign a9918 = ~a9916 & ~a9914;
assign a9920 = ~a9844 & ~a9134;
assign a9922 = a9920 & a9764;
assign a9924 = ~a9920 & ~a9764;
assign a9926 = ~a9924 & ~a9922;
assign a9928 = ~a9902 & ~a9896;
assign a9930 = ~a9928 & ~a9900;
assign a9932 = ~a9930 & ~a9926;
assign a9934 = a9930 & a9926;
assign a9936 = ~a9934 & ~a9932;
assign a9938 = a9936 & ~a9152;
assign a9940 = ~a9938 & ~a9918;
assign a9942 = ~a9936 & a9152;
assign a9944 = ~a9942 & ~a9940;
assign a9946 = ~a9844 & ~a9152;
assign a9948 = a9946 & a9790;
assign a9950 = ~a9946 & ~a9790;
assign a9952 = ~a9950 & ~a9948;
assign a9954 = ~a9930 & ~a9922;
assign a9956 = ~a9954 & ~a9924;
assign a9958 = ~a9956 & ~a9952;
assign a9960 = a9956 & a9952;
assign a9962 = ~a9960 & ~a9958;
assign a9964 = a9962 & a9158;
assign a9966 = ~a9964 & ~a9944;
assign a9968 = ~a9962 & ~a9158;
assign a9970 = ~a9968 & ~a9966;
assign a9972 = ~a9844 & a9158;
assign a9974 = a9972 & a9816;
assign a9976 = ~a9972 & ~a9816;
assign a9978 = ~a9976 & ~a9974;
assign a9980 = ~a9956 & ~a9948;
assign a9982 = ~a9980 & ~a9950;
assign a9984 = ~a9982 & ~a9978;
assign a9986 = a9982 & a9978;
assign a9988 = ~a9986 & ~a9984;
assign a9990 = a9988 & a9970;
assign a9992 = ~a9990 & ~a9116;
assign a9994 = ~a9992 & ~a9862;
assign a9996 = a9992 & a9862;
assign a9998 = ~a9990 & ~a9098;
assign a10000 = ~a9998 & ~a9876;
assign a10002 = ~a9990 & ~a9084;
assign a10004 = a10002 & ~a9870;
assign a10006 = a9998 & a9876;
assign a10008 = ~a10006 & ~a10004;
assign a10010 = ~a10008 & ~a10000;
assign a10012 = ~a10010 & ~a9996;
assign a10014 = ~a10012 & ~a9994;
assign a10016 = ~a9990 & ~a9134;
assign a10018 = ~a10016 & ~a9910;
assign a10020 = a10016 & a9910;
assign a10022 = ~a10020 & ~a10018;
assign a10024 = ~a10022 & ~a10014;
assign a10026 = a10022 & a10014;
assign a10028 = ~a10026 & ~a10024;
assign a10030 = i274 & ~i268;
assign a10032 = ~i274 & i268;
assign a10034 = ~a10032 & ~a10030;
assign a10036 = ~a10034 & ~a9180;
assign a10038 = ~a10036 & ~a9084;
assign a10040 = ~a10002 & a9870;
assign a10042 = ~a10040 & ~a10004;
assign a10044 = a10042 & ~a9098;
assign a10046 = ~a10044 & ~a10038;
assign a10048 = ~a10042 & a9098;
assign a10050 = ~a10048 & ~a10046;
assign a10052 = ~a10006 & ~a10000;
assign a10054 = ~a10052 & ~a10004;
assign a10056 = a10052 & a10004;
assign a10058 = ~a10056 & ~a10054;
assign a10060 = a10058 & ~a9116;
assign a10062 = ~a10060 & ~a10050;
assign a10064 = ~a10058 & a9116;
assign a10066 = ~a10064 & ~a10062;
assign a10068 = ~a9996 & ~a9994;
assign a10070 = ~a10068 & ~a10010;
assign a10072 = a10068 & a10010;
assign a10074 = ~a10072 & ~a10070;
assign a10076 = a10074 & ~a9134;
assign a10078 = ~a10076 & ~a10066;
assign a10080 = ~a10074 & a9134;
assign a10082 = ~a10080 & ~a10078;
assign a10084 = a10028 & ~a9152;
assign a10086 = ~a10084 & ~a10082;
assign a10088 = ~a10028 & a9152;
assign a10090 = ~a10088 & ~a10086;
assign a10092 = ~a9990 & ~a9152;
assign a10094 = a10092 & a9936;
assign a10096 = ~a10092 & ~a9936;
assign a10098 = ~a10096 & ~a10094;
assign a10100 = ~a10020 & ~a10014;
assign a10102 = ~a10100 & ~a10018;
assign a10104 = ~a10102 & ~a10098;
assign a10106 = a10102 & a10098;
assign a10108 = ~a10106 & ~a10104;
assign a10110 = a10108 & a9158;
assign a10112 = ~a10110 & ~a10090;
assign a10114 = ~a10108 & ~a9158;
assign a10116 = ~a10114 & ~a10112;
assign a10118 = ~a9990 & a9158;
assign a10120 = a10118 & a9962;
assign a10122 = ~a10118 & ~a9962;
assign a10124 = ~a10122 & ~a10120;
assign a10126 = ~a10102 & ~a10094;
assign a10128 = ~a10126 & ~a10096;
assign a10130 = ~a10128 & ~a10124;
assign a10132 = a10128 & a10124;
assign a10134 = ~a10132 & ~a10130;
assign a10136 = a10134 & a10116;
assign a10138 = ~a10136 & ~a9152;
assign a10140 = ~a10138 & ~a10028;
assign a10142 = a10138 & a10028;
assign a10144 = ~a10136 & ~a9134;
assign a10146 = ~a10144 & ~a10074;
assign a10148 = a10144 & a10074;
assign a10150 = ~a10136 & ~a9116;
assign a10152 = ~a10150 & ~a10058;
assign a10154 = a10150 & a10058;
assign a10156 = ~a10136 & ~a9098;
assign a10158 = ~a10156 & ~a10042;
assign a10160 = a10156 & a10042;
assign a10162 = ~a10136 & ~a9084;
assign a10164 = a10162 & ~a10036;
assign a10166 = ~a10164 & ~a10160;
assign a10168 = ~a10166 & ~a10158;
assign a10170 = ~a10168 & ~a10154;
assign a10172 = ~a10170 & ~a10152;
assign a10174 = ~a10172 & ~a10148;
assign a10176 = ~a10174 & ~a10146;
assign a10178 = ~a10176 & ~a10142;
assign a10180 = ~a10178 & ~a10140;
assign a10182 = ~a10136 & a9158;
assign a10184 = ~a10182 & ~a10108;
assign a10186 = a10182 & a10108;
assign a10188 = ~a10186 & ~a10184;
assign a10190 = ~a10188 & ~a10180;
assign a10192 = a10188 & a10180;
assign a10194 = ~a10192 & ~a10190;
assign a10196 = ~a9182 & ~a9084;
assign a10198 = ~a10162 & a10036;
assign a10200 = ~a10198 & ~a10164;
assign a10202 = a10200 & ~a9098;
assign a10204 = ~a10202 & ~a10196;
assign a10206 = ~a10200 & a9098;
assign a10208 = ~a10206 & ~a10204;
assign a10210 = ~a10160 & ~a10158;
assign a10212 = ~a10210 & ~a10164;
assign a10214 = a10210 & a10164;
assign a10216 = ~a10214 & ~a10212;
assign a10218 = a10216 & ~a9116;
assign a10220 = ~a10218 & ~a10208;
assign a10222 = ~a10216 & a9116;
assign a10224 = ~a10222 & ~a10220;
assign a10226 = ~a10154 & ~a10152;
assign a10228 = ~a10226 & ~a10168;
assign a10230 = a10226 & a10168;
assign a10232 = ~a10230 & ~a10228;
assign a10234 = a10232 & ~a9134;
assign a10236 = ~a10234 & ~a10224;
assign a10238 = ~a10232 & a9134;
assign a10240 = ~a10238 & ~a10236;
assign a10242 = ~a10148 & ~a10146;
assign a10244 = ~a10242 & ~a10172;
assign a10246 = a10242 & a10172;
assign a10248 = ~a10246 & ~a10244;
assign a10250 = a10248 & ~a9152;
assign a10252 = ~a10250 & ~a10240;
assign a10254 = ~a10248 & a9152;
assign a10256 = ~a10254 & ~a10252;
assign a10258 = ~a10142 & ~a10140;
assign a10260 = ~a10258 & ~a10176;
assign a10262 = a10258 & a10176;
assign a10264 = ~a10262 & ~a10260;
assign a10266 = a10264 & a9158;
assign a10268 = ~a10266 & ~a10256;
assign a10270 = ~a10264 & ~a9158;
assign a10272 = ~a10270 & ~a10268;
assign a10274 = a10272 & a10194;
assign a10276 = ~a10274 & ~a9084;
assign a10278 = a10276 & ~a9182;
assign a10280 = ~a10276 & a9182;
assign a10282 = ~a10280 & ~a10278;
assign a10284 = ~a10274 & ~a9098;
assign a10286 = ~a10284 & ~a10200;
assign a10288 = a10284 & a10200;
assign a10290 = ~a10288 & ~a10286;
assign a10292 = ~a10290 & ~a10278;
assign a10294 = a10290 & a10278;
assign a10296 = ~a10294 & ~a10292;
assign a10298 = ~a10296 & ~a10282;
assign a10300 = ~a10288 & ~a10278;
assign a10302 = ~a10300 & ~a10286;
assign a10304 = ~a10274 & ~a9116;
assign a10306 = ~a10304 & ~a10216;
assign a10308 = a10304 & a10216;
assign a10310 = ~a10308 & ~a10306;
assign a10312 = ~a10310 & ~a10302;
assign a10314 = a10310 & a10302;
assign a10316 = ~a10314 & ~a10312;
assign a10318 = ~a10316 & a10298;
assign a10320 = ~a10308 & ~a10302;
assign a10322 = ~a10320 & ~a10306;
assign a10324 = ~a10274 & ~a9134;
assign a10326 = ~a10324 & ~a10232;
assign a10328 = a10324 & a10232;
assign a10330 = ~a10328 & ~a10326;
assign a10332 = ~a10330 & ~a10322;
assign a10334 = a10330 & a10322;
assign a10336 = ~a10334 & ~a10332;
assign a10338 = ~a10336 & a10318;
assign a10340 = ~a10328 & ~a10322;
assign a10342 = ~a10340 & ~a10326;
assign a10344 = ~a10274 & ~a9152;
assign a10346 = ~a10344 & ~a10248;
assign a10348 = a10344 & a10248;
assign a10350 = ~a10348 & ~a10346;
assign a10352 = ~a10350 & ~a10342;
assign a10354 = a10350 & a10342;
assign a10356 = ~a10354 & ~a10352;
assign a10358 = ~a10356 & a10338;
assign a10360 = ~a10348 & ~a10342;
assign a10362 = ~a10360 & ~a10346;
assign a10364 = ~a10274 & a9158;
assign a10366 = ~a10364 & ~a10264;
assign a10368 = a10364 & a10264;
assign a10370 = ~a10368 & ~a10366;
assign a10372 = ~a10370 & ~a10362;
assign a10374 = a10370 & a10362;
assign a10376 = ~a10374 & ~a10372;
assign a10378 = ~a10376 & ~a10358;
assign a10380 = a10376 & a10358;
assign a10382 = ~a10380 & ~a10378;
assign a10384 = ~a10382 & ~a9168;
assign a10386 = a10384 & ~a9076;
assign a10388 = a10282 & ~a9168;
assign a10390 = a10388 & a3976;
assign a10392 = ~a10296 & a10282;
assign a10394 = a10296 & ~a10282;
assign a10396 = ~a10394 & ~a10392;
assign a10398 = ~a10396 & ~a9168;
assign a10400 = a10398 & a4980;
assign a10402 = ~a10400 & ~a10390;
assign a10404 = ~a10398 & ~a4980;
assign a10406 = ~a10404 & ~a10402;
assign a10408 = ~a10316 & ~a10298;
assign a10410 = a10316 & a10298;
assign a10412 = ~a10410 & ~a10408;
assign a10414 = ~a10412 & ~a9168;
assign a10416 = a10414 & a5028;
assign a10418 = ~a10416 & ~a10406;
assign a10420 = ~a10414 & ~a5028;
assign a10422 = ~a10420 & ~a10418;
assign a10424 = ~a10336 & ~a10318;
assign a10426 = a10336 & a10318;
assign a10428 = ~a10426 & ~a10424;
assign a10430 = ~a10428 & ~a9168;
assign a10432 = a10430 & a5076;
assign a10434 = ~a10432 & ~a10422;
assign a10436 = ~a10430 & ~a5076;
assign a10438 = ~a10436 & ~a10434;
assign a10440 = ~a10356 & ~a10338;
assign a10442 = a10356 & a10338;
assign a10444 = ~a10442 & ~a10440;
assign a10446 = ~a10444 & ~a9168;
assign a10448 = a10446 & a5124;
assign a10450 = ~a10448 & ~a10438;
assign a10452 = ~a10446 & ~a5124;
assign a10454 = ~a10452 & ~a10450;
assign a10456 = ~a10384 & a5172;
assign a10458 = a10384 & ~a5172;
assign a10460 = ~a10458 & ~a10456;
assign a10462 = ~a10460 & ~a10454;
assign a10464 = a10460 & a10454;
assign a10466 = ~a10464 & ~a10462;
assign a10468 = ~a10466 & a5178;
assign a10470 = ~a10468 & ~a5172;
assign a10472 = ~a10470 & a9076;
assign a10474 = ~a10472 & ~a10386;
assign a10476 = ~a10474 & ~l890;
assign a10478 = ~a10476 & ~a9074;
assign a10480 = ~l1288 & l890;
assign a10482 = ~a4690 & ~l890;
assign a10484 = ~a10482 & ~a10480;
assign a10486 = ~l1124 & l890;
assign a10488 = a10446 & ~a9076;
assign a10490 = ~a10446 & a5124;
assign a10492 = a10446 & ~a5124;
assign a10494 = ~a10492 & ~a10490;
assign a10496 = ~a10494 & ~a10438;
assign a10498 = a10494 & a10438;
assign a10500 = ~a10498 & ~a10496;
assign a10502 = ~a10500 & a5178;
assign a10504 = ~a5178 & a5124;
assign a10506 = ~a10504 & ~a10502;
assign a10508 = ~a10506 & a9076;
assign a10510 = ~a10508 & ~a10488;
assign a10512 = ~a10510 & ~l890;
assign a10514 = ~a10512 & ~a10486;
assign a10516 = ~l1292 & l890;
assign a10518 = ~a4530 & ~l890;
assign a10520 = ~a10518 & ~a10516;
assign a10522 = ~l1116 & l890;
assign a10524 = a10430 & ~a9076;
assign a10526 = ~a10430 & a5076;
assign a10528 = a10430 & ~a5076;
assign a10530 = ~a10528 & ~a10526;
assign a10532 = ~a10530 & ~a10422;
assign a10534 = a10530 & a10422;
assign a10536 = ~a10534 & ~a10532;
assign a10538 = ~a10536 & a5178;
assign a10540 = ~a5178 & a5076;
assign a10542 = ~a10540 & ~a10538;
assign a10544 = ~a10542 & a9076;
assign a10546 = ~a10544 & ~a10524;
assign a10548 = ~a10546 & ~l890;
assign a10550 = ~a10548 & ~a10522;
assign a10552 = ~l1296 & l890;
assign a10554 = ~a4370 & ~l890;
assign a10556 = ~a10554 & ~a10552;
assign a10558 = ~l1108 & l890;
assign a10560 = a10414 & ~a9076;
assign a10562 = ~a10414 & a5028;
assign a10564 = a10414 & ~a5028;
assign a10566 = ~a10564 & ~a10562;
assign a10568 = ~a10566 & ~a10406;
assign a10570 = a10566 & a10406;
assign a10572 = ~a10570 & ~a10568;
assign a10574 = ~a10572 & a5178;
assign a10576 = ~a5178 & a5028;
assign a10578 = ~a10576 & ~a10574;
assign a10580 = ~a10578 & a9076;
assign a10582 = ~a10580 & ~a10560;
assign a10584 = ~a10582 & ~l890;
assign a10586 = ~a10584 & ~a10558;
assign a10588 = ~l1300 & l890;
assign a10590 = ~a4224 & ~l890;
assign a10592 = ~a10590 & ~a10588;
assign a10594 = ~l1096 & l890;
assign a10596 = a10398 & ~a9076;
assign a10598 = ~a10398 & a4980;
assign a10600 = a10398 & ~a4980;
assign a10602 = ~a10600 & ~a10598;
assign a10604 = ~a10602 & ~a10390;
assign a10606 = a10602 & a10390;
assign a10608 = ~a10606 & ~a10604;
assign a10610 = ~a10608 & a5178;
assign a10612 = ~a5178 & a4980;
assign a10614 = ~a10612 & ~a10610;
assign a10616 = ~a10614 & a9076;
assign a10618 = ~a10616 & ~a10596;
assign a10620 = ~a10618 & ~l890;
assign a10622 = ~a10620 & ~a10594;
assign a10624 = ~l1014 & l890;
assign a10626 = a10388 & ~a9076;
assign a10628 = ~a10388 & a3976;
assign a10630 = a10388 & ~a3976;
assign a10632 = ~a10630 & ~a10628;
assign a10634 = ~a10632 & a5178;
assign a10636 = ~a5178 & a3976;
assign a10638 = ~a10636 & ~a10634;
assign a10640 = ~a10638 & a9076;
assign a10642 = ~a10640 & ~a10626;
assign a10644 = ~a10642 & ~l890;
assign a10646 = ~a10644 & ~a10624;
assign a10648 = ~l1304 & l890;
assign a10650 = ~a4108 & ~l890;
assign a10652 = ~a10650 & ~a10648;
assign a10654 = a10646 & ~l1306;
assign a10656 = a10654 & a10652;
assign a10658 = ~a10656 & a10646;
assign a10660 = ~a10658 & a10622;
assign a10662 = a10646 & l1306;
assign a10664 = a10662 & ~a10652;
assign a10666 = a10664 & ~a10622;
assign a10668 = ~a10666 & ~a10660;
assign a10670 = ~a10668 & ~l1302;
assign a10672 = a10654 & ~a10652;
assign a10674 = a10672 & ~a10622;
assign a10676 = ~a10674 & ~a10670;
assign a10678 = ~a10676 & a10592;
assign a10680 = ~a10658 & ~a10622;
assign a10682 = ~a10680 & ~a10678;
assign a10684 = a10662 & a10652;
assign a10686 = a10684 & ~a10622;
assign a10688 = a10686 & ~l1302;
assign a10690 = ~a10688 & a10682;
assign a10692 = ~a10690 & a10586;
assign a10694 = ~a10668 & l1302;
assign a10696 = a10684 & a10622;
assign a10698 = ~a10696 & ~a10694;
assign a10700 = ~a10698 & ~a10592;
assign a10702 = a10672 & a10622;
assign a10704 = a10702 & l1302;
assign a10706 = ~a10704 & ~a10700;
assign a10708 = a10664 & a10622;
assign a10710 = ~a10708 & a10706;
assign a10712 = ~a10710 & ~a10586;
assign a10714 = ~a10712 & ~a10692;
assign a10716 = ~a10714 & ~l1298;
assign a10718 = ~a10676 & ~a10592;
assign a10720 = a10702 & ~l1302;
assign a10722 = ~a10720 & ~a10718;
assign a10724 = ~a10722 & ~a10586;
assign a10726 = ~a10724 & ~a10716;
assign a10728 = ~a10726 & a10556;
assign a10730 = ~a10690 & ~a10586;
assign a10732 = ~a10730 & ~a10728;
assign a10734 = ~a10698 & a10592;
assign a10736 = a10686 & l1302;
assign a10738 = ~a10736 & ~a10734;
assign a10740 = ~a10738 & ~a10586;
assign a10742 = a10740 & ~l1298;
assign a10744 = ~a10742 & a10732;
assign a10746 = ~a10744 & a10550;
assign a10748 = ~a10714 & l1298;
assign a10750 = ~a10738 & a10586;
assign a10752 = ~a10750 & ~a10748;
assign a10754 = ~a10752 & ~a10556;
assign a10756 = ~a10722 & a10586;
assign a10758 = a10756 & l1298;
assign a10760 = ~a10758 & ~a10754;
assign a10762 = ~a10710 & a10586;
assign a10764 = ~a10762 & a10760;
assign a10766 = ~a10764 & ~a10550;
assign a10768 = ~a10766 & ~a10746;
assign a10770 = ~a10768 & ~l1294;
assign a10772 = ~a10726 & ~a10556;
assign a10774 = a10756 & ~l1298;
assign a10776 = ~a10774 & ~a10772;
assign a10778 = ~a10776 & ~a10550;
assign a10780 = ~a10778 & ~a10770;
assign a10782 = ~a10780 & a10520;
assign a10784 = ~a10744 & ~a10550;
assign a10786 = ~a10784 & ~a10782;
assign a10788 = ~a10752 & a10556;
assign a10790 = a10740 & l1298;
assign a10792 = ~a10790 & ~a10788;
assign a10794 = ~a10792 & ~a10550;
assign a10796 = a10794 & ~l1294;
assign a10798 = ~a10796 & a10786;
assign a10800 = ~a10798 & a10514;
assign a10802 = ~a10768 & l1294;
assign a10804 = ~a10792 & a10550;
assign a10806 = ~a10804 & ~a10802;
assign a10808 = ~a10806 & ~a10520;
assign a10810 = ~a10776 & a10550;
assign a10812 = a10810 & l1294;
assign a10814 = ~a10812 & ~a10808;
assign a10816 = ~a10764 & a10550;
assign a10818 = ~a10816 & a10814;
assign a10820 = ~a10818 & ~a10514;
assign a10822 = ~a10820 & ~a10800;
assign a10824 = ~a10822 & ~l1290;
assign a10826 = ~a10780 & ~a10520;
assign a10828 = a10810 & ~l1294;
assign a10830 = ~a10828 & ~a10826;
assign a10832 = ~a10830 & ~a10514;
assign a10834 = ~a10832 & ~a10824;
assign a10836 = ~a10834 & a10484;
assign a10838 = ~a10798 & ~a10514;
assign a10840 = ~a10838 & ~a10836;
assign a10842 = ~a10806 & a10520;
assign a10844 = a10794 & l1294;
assign a10846 = ~a10844 & ~a10842;
assign a10848 = ~a10846 & ~a10514;
assign a10850 = a10848 & ~l1290;
assign a10852 = ~a10850 & a10840;
assign a10854 = ~a10852 & a10478;
assign a10856 = ~a10822 & l1290;
assign a10858 = ~a10846 & a10514;
assign a10860 = ~a10858 & ~a10856;
assign a10862 = ~a10860 & ~a10484;
assign a10864 = ~a10830 & a10514;
assign a10866 = a10864 & l1290;
assign a10868 = ~a10866 & ~a10862;
assign a10870 = ~a10818 & a10514;
assign a10872 = ~a10870 & a10868;
assign a10874 = ~a10872 & ~a10478;
assign a10876 = ~a10874 & ~a10854;
assign a10878 = ~a10876 & ~l1286;
assign a10880 = ~a10834 & ~a10484;
assign a10882 = a10864 & ~l1290;
assign a10884 = ~a10882 & ~a10880;
assign a10886 = ~a10884 & ~a10478;
assign a10888 = ~a10886 & ~a10878;
assign a10890 = ~a10888 & a9072;
assign a10892 = ~a10852 & ~a10478;
assign a10894 = ~a10892 & ~a10890;
assign a10896 = ~a10860 & a10484;
assign a10898 = a10848 & l1290;
assign a10900 = ~a10898 & ~a10896;
assign a10902 = ~a10900 & ~a10478;
assign a10904 = a10902 & ~l1286;
assign a10906 = ~a10904 & a10894;
assign a10908 = ~a10906 & ~l1140;
assign a10910 = ~a10876 & l1286;
assign a10912 = ~a10900 & a10478;
assign a10914 = ~a10912 & ~a10910;
assign a10916 = ~a10914 & ~a9072;
assign a10918 = ~a10884 & a10478;
assign a10920 = a10918 & l1286;
assign a10922 = ~a10920 & ~a10916;
assign a10924 = ~a10872 & a10478;
assign a10926 = ~a10924 & a10922;
assign a10928 = ~a10926 & l1140;
assign a10930 = ~a10928 & ~a10908;
assign a10932 = ~a10930 & ~l1282;
assign a10934 = ~a10888 & ~a9072;
assign a10936 = a10918 & ~l1286;
assign a10938 = ~a10936 & ~a10934;
assign a10940 = ~a10938 & l1140;
assign a10942 = ~a10940 & ~a10932;
assign a10944 = ~a10942 & ~l1280;
assign a10946 = ~a10906 & l1140;
assign a10948 = ~a10946 & ~a10944;
assign a10950 = ~a10914 & a9072;
assign a10952 = a10902 & l1286;
assign a10954 = ~a10952 & ~a10950;
assign a10956 = ~a10954 & l1140;
assign a10958 = a10956 & ~l1282;
assign a10960 = ~a10958 & a10948;
assign a10962 = ~a10960 & ~l1194;
assign a10964 = ~a10930 & l1282;
assign a10966 = ~a10954 & ~l1140;
assign a10968 = ~a10966 & ~a10964;
assign a10970 = ~a10968 & ~l1280;
assign a10972 = a10956 & l1282;
assign a10974 = ~a10972 & ~a10970;
assign a10976 = ~a10974 & l1194;
assign a10978 = ~a10976 & ~a10962;
assign a10980 = ~a10978 & ~l1278;
assign a10982 = ~a10978 & l1278;
assign a10984 = ~a10942 & l1280;
assign a10986 = ~a10938 & ~l1140;
assign a10988 = a10986 & ~l1282;
assign a10990 = ~a10988 & ~a10984;
assign a10992 = ~a10990 & ~l1194;
assign a10994 = ~a10968 & l1280;
assign a10996 = a10986 & l1282;
assign a10998 = ~a10996 & ~a10994;
assign a11000 = ~a10926 & ~l1140;
assign a11002 = ~a11000 & a10998;
assign a11004 = ~a11002 & l1194;
assign a11006 = ~a11004 & ~a10992;
assign a11008 = ~a11006 & ~l1278;
assign a11010 = ~a11008 & ~a10982;
assign a11012 = ~a11010 & l992;
assign a11014 = ~a11012 & ~a10980;
assign a11016 = ~a10960 & l1194;
assign a11018 = ~a10974 & ~l1194;
assign a11020 = ~a11018 & ~a11016;
assign a11022 = ~a11020 & ~l1278;
assign a11024 = ~a10990 & l1194;
assign a11026 = ~a11002 & ~l1194;
assign a11028 = ~a11026 & ~a11024;
assign a11030 = ~a11028 & l1278;
assign a11032 = ~a11030 & ~a11022;
assign a11034 = ~a11032 & ~l992;
assign a11036 = ~a11034 & a11014;
assign a11038 = ~a11020 & l1278;
assign a11040 = ~a11038 & a11036;
assign a11042 = ~a11006 & l1278;
assign a11044 = ~a11042 & a11040;
assign a11046 = ~a11028 & ~l1278;
assign a11048 = ~a11046 & a11044;
assign a11050 = ~a11048 & ~l1000;
assign a11052 = a11050 & l1272;
assign a11054 = a11052 & ~l1266;
assign a11056 = ~a11048 & l1000;
assign a11058 = a11056 & l1272;
assign a11060 = a11058 & ~l1266;
assign a11062 = a11060 & l1308;
assign a11064 = ~a11062 & ~a11054;
assign a11066 = ~a11064 & ~l1260;
assign a11068 = ~l1310 & l890;
assign a11070 = ~a2706 & a2564;
assign a11072 = ~a2712 & a2706;
assign a11074 = ~a11072 & ~a11070;
assign a11076 = ~a11074 & ~a4080;
assign a11078 = ~a11076 & ~a2722;
assign a11080 = ~a11078 & ~a2706;
assign a11082 = i74 & ~i50;
assign a11084 = ~a11082 & ~a4864;
assign a11086 = ~i74 & i50;
assign a11088 = ~a11086 & ~a11084;
assign a11090 = a11088 & a4122;
assign a11092 = ~a11080 & ~a4098;
assign a11094 = ~a4104 & a2722;
assign a11096 = a11094 & a4080;
assign a11098 = ~a4108 & ~a4080;
assign a11100 = ~a11098 & ~a11096;
assign a11102 = a11100 & ~a11092;
assign a11104 = ~a11102 & a4138;
assign a11106 = ~a11080 & ~a4212;
assign a11108 = ~a4218 & a2722;
assign a11110 = a11108 & a4080;
assign a11112 = ~a4224 & ~a4080;
assign a11114 = ~a11112 & ~a11110;
assign a11116 = a11114 & ~a11106;
assign a11118 = ~a11116 & a4264;
assign a11120 = ~a11118 & ~a11104;
assign a11122 = a11116 & ~a4264;
assign a11124 = ~a11122 & ~a11120;
assign a11126 = ~a11080 & ~a4358;
assign a11128 = ~a4364 & a2722;
assign a11130 = a11128 & a4080;
assign a11132 = ~a4370 & ~a4080;
assign a11134 = ~a11132 & ~a11130;
assign a11136 = a11134 & ~a11126;
assign a11138 = ~a11136 & a4416;
assign a11140 = ~a11138 & ~a11124;
assign a11142 = a11136 & ~a4416;
assign a11144 = ~a11142 & ~a11140;
assign a11146 = ~a11080 & ~a4518;
assign a11148 = ~a4524 & a2722;
assign a11150 = a11148 & a4080;
assign a11152 = ~a4530 & ~a4080;
assign a11154 = ~a11152 & ~a11150;
assign a11156 = a11154 & ~a11146;
assign a11158 = ~a11156 & a4576;
assign a11160 = ~a11158 & ~a11144;
assign a11162 = a11156 & ~a4576;
assign a11164 = ~a11162 & ~a11160;
assign a11166 = ~a11080 & ~a4678;
assign a11168 = ~a4684 & a2722;
assign a11170 = a11168 & a4080;
assign a11172 = ~a4690 & ~a4080;
assign a11174 = ~a11172 & ~a11170;
assign a11176 = a11174 & ~a11166;
assign a11178 = ~a11176 & a4736;
assign a11180 = ~a11178 & ~a11164;
assign a11182 = a11176 & ~a4736;
assign a11184 = ~a11182 & ~a11180;
assign a11186 = ~a11080 & ~a4820;
assign a11188 = ~a4826 & a2722;
assign a11190 = a11188 & a4080;
assign a11192 = ~a4832 & ~a4080;
assign a11194 = ~a11192 & ~a11190;
assign a11196 = a11194 & ~a11186;
assign a11198 = ~a11196 & a4884;
assign a11200 = ~a11198 & ~a11184;
assign a11202 = a11196 & ~a4884;
assign a11204 = ~a11202 & ~a11200;
assign a11206 = ~a11080 & a4934;
assign a11208 = a4934 & i14;
assign a11210 = a11208 & a4080;
assign a11212 = ~a11210 & ~a11206;
assign a11214 = a11212 & ~a11204;
assign a11216 = ~a11214 & ~a11090;
assign a11218 = ~a11216 & a11080;
assign a11220 = a11218 & i188;
assign a11222 = a11220 & ~a4080;
assign a11224 = ~a11220 & a4080;
assign a11226 = ~a11224 & ~a11222;
assign a11228 = a11220 & a4080;
assign a11230 = ~a11228 & a11226;
assign a11232 = ~a11226 & a4146;
assign a11234 = a11226 & ~a4146;
assign a11236 = ~a11234 & ~a11232;
assign a11238 = ~a11228 & a2736;
assign a11240 = ~a11238 & a11236;
assign a11242 = ~a11240 & ~a2712;
assign a11244 = ~a11242 & ~a4178;
assign a11246 = ~a4178 & i92;
assign a11248 = i190 & ~i92;
assign a11250 = ~a11248 & ~a11246;
assign a11252 = ~a11250 & a4140;
assign a11254 = a11252 & a11226;
assign a11256 = i192 & ~i92;
assign a11258 = ~a11256 & ~a5572;
assign a11260 = a11258 & a5576;
assign a11262 = a11260 & ~a11250;
assign a11264 = ~a11262 & ~a11094;
assign a11266 = ~a11264 & ~a11226;
assign a11268 = ~a11266 & ~a11254;
assign a11270 = ~a11268 & ~a11230;
assign a11272 = ~a11250 & a5588;
assign a11274 = ~a11272 & a4108;
assign a11276 = ~a11274 & a11226;
assign a11278 = a11276 & a11230;
assign a11280 = ~a11278 & ~a11270;
assign a11282 = a11280 & ~a11244;
assign a11284 = i220 & i218;
assign a11286 = a11284 & i216;
assign a11288 = a11286 & i214;
assign a11290 = a11288 & ~i222;
assign a11292 = ~a11290 & i212;
assign a11294 = a11252 & ~a11226;
assign a11296 = ~a11264 & a11226;
assign a11298 = ~a11296 & ~a11294;
assign a11300 = ~a11298 & a11228;
assign a11302 = ~a11274 & ~a11226;
assign a11304 = ~a11302 & ~a11300;
assign a11306 = ~a11304 & a11292;
assign a11308 = a11304 & ~a11292;
assign a11310 = ~a11308 & ~a11306;
assign a11312 = ~a11310 & a2712;
assign a11314 = a11216 & i182;
assign a11316 = a11314 & ~i184;
assign a11318 = a4122 & ~i186;
assign a11320 = ~a11318 & a11316;
assign a11322 = ~a11282 & a4138;
assign a11324 = ~a11242 & ~a4304;
assign a11326 = ~a4304 & i92;
assign a11328 = i200 & ~i92;
assign a11330 = ~a11328 & ~a11326;
assign a11332 = ~a11330 & a4140;
assign a11334 = a11332 & a11226;
assign a11336 = ~a11330 & a11260;
assign a11338 = ~a11336 & ~a11108;
assign a11340 = ~a11338 & ~a11226;
assign a11342 = ~a11340 & ~a11334;
assign a11344 = ~a11342 & ~a11230;
assign a11346 = ~a11330 & a5588;
assign a11348 = ~a11346 & a4224;
assign a11350 = ~a11348 & a11226;
assign a11352 = a11350 & a11230;
assign a11354 = ~a11352 & ~a11344;
assign a11356 = a11354 & ~a11324;
assign a11358 = ~a11356 & a4264;
assign a11360 = ~a11358 & ~a11322;
assign a11362 = a11356 & ~a4264;
assign a11364 = ~a11362 & ~a11360;
assign a11366 = ~a11242 & ~a4464;
assign a11368 = ~a4464 & i92;
assign a11370 = i202 & ~i92;
assign a11372 = ~a11370 & ~a11368;
assign a11374 = ~a11372 & a4140;
assign a11376 = a11374 & a11226;
assign a11378 = ~a11372 & a11260;
assign a11380 = ~a11378 & ~a11128;
assign a11382 = ~a11380 & ~a11226;
assign a11384 = ~a11382 & ~a11376;
assign a11386 = ~a11384 & ~a11230;
assign a11388 = ~a11372 & a5588;
assign a11390 = ~a11388 & a4370;
assign a11392 = ~a11390 & a11226;
assign a11394 = a11392 & a11230;
assign a11396 = ~a11394 & ~a11386;
assign a11398 = a11396 & ~a11366;
assign a11400 = ~a11398 & a4416;
assign a11402 = ~a11400 & ~a11364;
assign a11404 = a11398 & ~a4416;
assign a11406 = ~a11404 & ~a11402;
assign a11408 = ~a11242 & ~a4624;
assign a11410 = ~a4624 & i92;
assign a11412 = i204 & ~i92;
assign a11414 = ~a11412 & ~a11410;
assign a11416 = ~a11414 & a4140;
assign a11418 = a11416 & a11226;
assign a11420 = ~a11414 & a11260;
assign a11422 = ~a11420 & ~a11148;
assign a11424 = ~a11422 & ~a11226;
assign a11426 = ~a11424 & ~a11418;
assign a11428 = ~a11426 & ~a11230;
assign a11430 = ~a11414 & a5588;
assign a11432 = ~a11430 & a4530;
assign a11434 = ~a11432 & a11226;
assign a11436 = a11434 & a11230;
assign a11438 = ~a11436 & ~a11428;
assign a11440 = a11438 & ~a11408;
assign a11442 = ~a11440 & a4576;
assign a11444 = ~a11442 & ~a11406;
assign a11446 = a11440 & ~a4576;
assign a11448 = ~a11446 & ~a11444;
assign a11450 = ~a11242 & ~a4784;
assign a11452 = ~a4784 & i92;
assign a11454 = i206 & ~i92;
assign a11456 = ~a11454 & ~a11452;
assign a11458 = ~a11456 & a4140;
assign a11460 = a11458 & a11226;
assign a11462 = ~a11456 & a11260;
assign a11464 = ~a11462 & ~a11168;
assign a11466 = ~a11464 & ~a11226;
assign a11468 = ~a11466 & ~a11460;
assign a11470 = ~a11468 & ~a11230;
assign a11472 = ~a11456 & a5588;
assign a11474 = ~a11472 & a4690;
assign a11476 = ~a11474 & a11226;
assign a11478 = a11476 & a11230;
assign a11480 = ~a11478 & ~a11470;
assign a11482 = a11480 & ~a11450;
assign a11484 = ~a11482 & a4736;
assign a11486 = ~a11484 & ~a11448;
assign a11488 = a11482 & ~a4736;
assign a11490 = ~a11488 & ~a11486;
assign a11492 = ~a11242 & ~a4916;
assign a11494 = ~a4916 & i92;
assign a11496 = i208 & ~i92;
assign a11498 = ~a11496 & ~a11494;
assign a11500 = ~a11498 & a4140;
assign a11502 = a11500 & a11226;
assign a11504 = ~a11498 & a11260;
assign a11506 = ~a11504 & ~a11188;
assign a11508 = ~a11506 & ~a11226;
assign a11510 = ~a11508 & ~a11502;
assign a11512 = ~a11510 & ~a11230;
assign a11514 = ~a11498 & a5588;
assign a11516 = ~a11514 & a4832;
assign a11518 = ~a11516 & a11226;
assign a11520 = a11518 & a11230;
assign a11522 = ~a11520 & ~a11512;
assign a11524 = a11522 & ~a11492;
assign a11526 = ~a11524 & a4884;
assign a11528 = ~a11526 & ~a11490;
assign a11530 = a11524 & ~a4884;
assign a11532 = ~a11530 & ~a11528;
assign a11534 = ~a11242 & ~a4946;
assign a11536 = ~a4946 & i92;
assign a11538 = i210 & ~i92;
assign a11540 = ~a11538 & ~a11536;
assign a11542 = ~a11540 & a4140;
assign a11544 = a11542 & a11226;
assign a11546 = ~a11540 & a11260;
assign a11548 = ~a11546 & ~a11208;
assign a11550 = ~a11548 & ~a11226;
assign a11552 = ~a11550 & ~a11544;
assign a11554 = ~a11552 & ~a11230;
assign a11556 = ~a11554 & ~a11534;
assign a11558 = ~a11556 & ~a11090;
assign a11560 = ~a11558 & ~a11532;
assign a11562 = a11556 & a11090;
assign a11564 = ~a11562 & ~a11560;
assign a11566 = a11564 & a11318;
assign a11568 = ~a11566 & ~a11320;
assign a11570 = a11292 & ~a4138;
assign a11572 = ~a11292 & a4138;
assign a11574 = ~a11572 & ~a11570;
assign a11576 = ~a11574 & ~a11568;
assign a11578 = a11568 & ~a4138;
assign a11580 = ~a11578 & ~a11576;
assign a11582 = ~a11580 & ~a2712;
assign a11584 = ~a11582 & ~a11312;
assign a11586 = a11584 & ~a11282;
assign a11588 = ~a11304 & ~a11292;
assign a11590 = a11332 & ~a11226;
assign a11592 = ~a11338 & a11226;
assign a11594 = ~a11592 & ~a11590;
assign a11596 = ~a11594 & a11228;
assign a11598 = ~a11348 & ~a11226;
assign a11600 = ~a11598 & ~a11596;
assign a11602 = ~a11600 & i214;
assign a11604 = a11600 & ~i214;
assign a11606 = ~a11604 & ~a11602;
assign a11608 = ~a11606 & ~a11588;
assign a11610 = a11606 & a11588;
assign a11612 = ~a11610 & ~a11608;
assign a11614 = ~a11612 & a2712;
assign a11616 = ~a11292 & ~a4138;
assign a11618 = ~a4264 & i214;
assign a11620 = a4264 & ~i214;
assign a11622 = ~a11620 & ~a11618;
assign a11624 = ~a11622 & ~a11616;
assign a11626 = a11622 & a11616;
assign a11628 = ~a11626 & ~a11624;
assign a11630 = ~a11628 & ~a11568;
assign a11632 = a11568 & ~a4264;
assign a11634 = ~a11632 & ~a11630;
assign a11636 = ~a11634 & ~a2712;
assign a11638 = ~a11636 & ~a11614;
assign a11640 = a11638 & ~a11356;
assign a11642 = ~a11640 & ~a11586;
assign a11644 = ~a11638 & a11356;
assign a11646 = ~a11644 & ~a11642;
assign a11648 = ~a11600 & ~i214;
assign a11650 = ~a11648 & ~a11588;
assign a11652 = a11600 & i214;
assign a11654 = ~a11652 & ~a11650;
assign a11656 = a11374 & ~a11226;
assign a11658 = ~a11380 & a11226;
assign a11660 = ~a11658 & ~a11656;
assign a11662 = ~a11660 & a11228;
assign a11664 = ~a11390 & ~a11226;
assign a11666 = ~a11664 & ~a11662;
assign a11668 = ~a11666 & i216;
assign a11670 = a11666 & ~i216;
assign a11672 = ~a11670 & ~a11668;
assign a11674 = ~a11672 & ~a11654;
assign a11676 = a11672 & a11654;
assign a11678 = ~a11676 & ~a11674;
assign a11680 = ~a11678 & a2712;
assign a11682 = ~a4264 & ~i214;
assign a11684 = ~a11682 & ~a11616;
assign a11686 = a4264 & i214;
assign a11688 = ~a11686 & ~a11684;
assign a11690 = ~a4416 & i216;
assign a11692 = a4416 & ~i216;
assign a11694 = ~a11692 & ~a11690;
assign a11696 = ~a11694 & ~a11688;
assign a11698 = a11694 & a11688;
assign a11700 = ~a11698 & ~a11696;
assign a11702 = ~a11700 & ~a11568;
assign a11704 = a11568 & ~a4416;
assign a11706 = ~a11704 & ~a11702;
assign a11708 = ~a11706 & ~a2712;
assign a11710 = ~a11708 & ~a11680;
assign a11712 = a11710 & ~a11398;
assign a11714 = ~a11712 & ~a11646;
assign a11716 = ~a11710 & a11398;
assign a11718 = ~a11716 & ~a11714;
assign a11720 = ~a11666 & ~i216;
assign a11722 = ~a11720 & ~a11654;
assign a11724 = a11666 & i216;
assign a11726 = ~a11724 & ~a11722;
assign a11728 = a11416 & ~a11226;
assign a11730 = ~a11422 & a11226;
assign a11732 = ~a11730 & ~a11728;
assign a11734 = ~a11732 & a11228;
assign a11736 = ~a11432 & ~a11226;
assign a11738 = ~a11736 & ~a11734;
assign a11740 = ~a11738 & i220;
assign a11742 = a11738 & ~i220;
assign a11744 = ~a11742 & ~a11740;
assign a11746 = ~a11744 & ~a11726;
assign a11748 = a11744 & a11726;
assign a11750 = ~a11748 & ~a11746;
assign a11752 = ~a11750 & a2712;
assign a11754 = ~a4416 & ~i216;
assign a11756 = ~a11754 & ~a11688;
assign a11758 = a4416 & i216;
assign a11760 = ~a11758 & ~a11756;
assign a11762 = ~a4576 & i220;
assign a11764 = a4576 & ~i220;
assign a11766 = ~a11764 & ~a11762;
assign a11768 = ~a11766 & ~a11760;
assign a11770 = a11766 & a11760;
assign a11772 = ~a11770 & ~a11768;
assign a11774 = ~a11772 & ~a11568;
assign a11776 = a11568 & ~a4576;
assign a11778 = ~a11776 & ~a11774;
assign a11780 = ~a11778 & ~a2712;
assign a11782 = ~a11780 & ~a11752;
assign a11784 = a11782 & ~a11440;
assign a11786 = ~a11784 & ~a11718;
assign a11788 = ~a11782 & a11440;
assign a11790 = ~a11788 & ~a11786;
assign a11792 = ~a11738 & ~i220;
assign a11794 = ~a11792 & ~a11726;
assign a11796 = a11738 & i220;
assign a11798 = ~a11796 & ~a11794;
assign a11800 = a11458 & ~a11226;
assign a11802 = ~a11464 & a11226;
assign a11804 = ~a11802 & ~a11800;
assign a11806 = ~a11804 & a11228;
assign a11808 = ~a11474 & ~a11226;
assign a11810 = ~a11808 & ~a11806;
assign a11812 = ~a11810 & i218;
assign a11814 = a11810 & ~i218;
assign a11816 = ~a11814 & ~a11812;
assign a11818 = ~a11816 & ~a11798;
assign a11820 = a11816 & a11798;
assign a11822 = ~a11820 & ~a11818;
assign a11824 = ~a11822 & a2712;
assign a11826 = ~a4576 & ~i220;
assign a11828 = ~a11826 & ~a11760;
assign a11830 = a4576 & i220;
assign a11832 = ~a11830 & ~a11828;
assign a11834 = ~a4736 & i218;
assign a11836 = a4736 & ~i218;
assign a11838 = ~a11836 & ~a11834;
assign a11840 = ~a11838 & ~a11832;
assign a11842 = a11838 & a11832;
assign a11844 = ~a11842 & ~a11840;
assign a11846 = ~a11844 & ~a11568;
assign a11848 = a11568 & ~a4736;
assign a11850 = ~a11848 & ~a11846;
assign a11852 = ~a11850 & ~a2712;
assign a11854 = ~a11852 & ~a11824;
assign a11856 = a11854 & ~a11482;
assign a11858 = ~a11856 & ~a11790;
assign a11860 = ~a11854 & a11482;
assign a11862 = ~a11860 & ~a11858;
assign a11864 = ~a11810 & ~i218;
assign a11866 = ~a11864 & ~a11798;
assign a11868 = a11810 & i218;
assign a11870 = ~a11868 & ~a11866;
assign a11872 = a11500 & ~a11226;
assign a11874 = ~a11506 & a11226;
assign a11876 = ~a11874 & ~a11872;
assign a11878 = ~a11876 & a11228;
assign a11880 = ~a11516 & ~a11226;
assign a11882 = ~a11880 & ~a11878;
assign a11884 = ~a11882 & ~i222;
assign a11886 = a11882 & i222;
assign a11888 = ~a11886 & ~a11884;
assign a11890 = ~a11888 & ~a11870;
assign a11892 = a11888 & a11870;
assign a11894 = ~a11892 & ~a11890;
assign a11896 = ~a11894 & a2712;
assign a11898 = ~a4736 & ~i218;
assign a11900 = ~a11898 & ~a11832;
assign a11902 = a4736 & i218;
assign a11904 = ~a11902 & ~a11900;
assign a11906 = ~a4884 & ~i222;
assign a11908 = a4884 & i222;
assign a11910 = ~a11908 & ~a11906;
assign a11912 = ~a11910 & ~a11904;
assign a11914 = a11910 & a11904;
assign a11916 = ~a11914 & ~a11912;
assign a11918 = ~a11916 & ~a11568;
assign a11920 = a11568 & ~a4884;
assign a11922 = ~a11920 & ~a11918;
assign a11924 = ~a11922 & ~a2712;
assign a11926 = ~a11924 & ~a11896;
assign a11928 = a11926 & ~a11524;
assign a11930 = ~a11928 & ~a11862;
assign a11932 = ~a11926 & a11524;
assign a11934 = ~a11932 & ~a11930;
assign a11936 = ~a4884 & i222;
assign a11938 = ~a11936 & ~a11904;
assign a11940 = a4884 & ~i222;
assign a11942 = ~a11940 & ~a11938;
assign a11944 = ~a11942 & a11090;
assign a11946 = a11942 & ~a11090;
assign a11948 = ~a11946 & ~a11944;
assign a11950 = ~a11948 & ~a11568;
assign a11952 = ~a11950 & ~a11090;
assign a11954 = a11952 & ~a11556;
assign a11956 = ~a11954 & ~a11934;
assign a11958 = ~a11952 & a11556;
assign a11960 = ~a11958 & ~a11956;
assign a11962 = ~a11960 & a11242;
assign a11964 = a11962 & i334;
assign a11966 = a11964 & ~a11230;
assign a11968 = ~a11964 & a11228;
assign a11970 = ~a11968 & ~a11966;
assign a11972 = ~a11970 & ~l890;
assign a11974 = ~a11972 & ~a11068;
assign a11976 = a11060 & ~l1308;
assign a11978 = a11976 & ~l1260;
assign a11980 = a11978 & ~a11974;
assign a11982 = ~a11980 & ~a11066;
assign a11984 = ~a11982 & l1252;
assign a11986 = ~l1312 & l890;
assign a11988 = a11964 & a11226;
assign a11990 = ~a11964 & ~a11226;
assign a11992 = ~a11990 & ~a11988;
assign a11994 = ~a11992 & ~l890;
assign a11996 = ~a11994 & ~a11986;
assign a11998 = a11978 & a11974;
assign a12000 = a11998 & l1252;
assign a12002 = a12000 & a11996;
assign a12004 = ~a12002 & ~a11984;
assign a12006 = a11050 & ~l1272;
assign a12008 = a12006 & ~l1266;
assign a12010 = a12008 & ~l1308;
assign a12012 = a12006 & l1266;
assign a12014 = a11058 & l1266;
assign a12016 = ~a12014 & ~a12012;
assign a12018 = ~a12016 & l1308;
assign a12020 = ~a12018 & ~a12010;
assign a12022 = ~a12020 & ~l1260;
assign a12024 = a12022 & a11974;
assign a12026 = ~a12020 & l1260;
assign a12028 = a11976 & l1260;
assign a12030 = ~a12028 & ~a12026;
assign a12032 = ~a12030 & ~a11974;
assign a12034 = ~a12032 & ~a12024;
assign a12036 = ~a12034 & ~l1252;
assign a12038 = a11998 & ~l1252;
assign a12040 = ~a12038 & ~a12036;
assign a12042 = ~a12040 & a11996;
assign a12044 = ~a12034 & l1252;
assign a12046 = a12044 & ~a11996;
assign a12048 = ~a12046 & ~a12042;
assign a12050 = a12000 & ~a11996;
assign a12052 = ~a12050 & a12048;
assign a12054 = ~a11010 & ~l992;
assign a12056 = ~a12054 & a12052;
assign a12058 = ~a11032 & l992;
assign a12060 = ~a12058 & a12056;
assign a12062 = ~a12040 & ~a11996;
assign a12064 = a12044 & a11996;
assign a12066 = ~a12064 & ~a12062;
assign a12068 = a12022 & ~a11974;
assign a12070 = ~a12068 & a12066;
assign a12072 = ~a12030 & a11974;
assign a12074 = ~a12072 & a12070;
assign a12076 = a12008 & l1308;
assign a12078 = ~a12076 & a12074;
assign a12080 = ~a12016 & ~l1308;
assign a12082 = ~a12080 & a12078;
assign a12084 = ~a11982 & ~l1252;
assign a12086 = ~a12084 & a12082;
assign a12088 = ~a11064 & l1260;
assign a12090 = ~a12088 & a12086;
assign a12092 = a11052 & l1266;
assign a12094 = ~a12092 & a12090;
assign a12096 = a11056 & ~l1272;
assign a12098 = ~a12096 & a12094;
assign a12100 = ~l1492 & l890;
assign a12102 = ~a2710 & ~l890;
assign a12104 = ~a12102 & ~a12100;
assign a12106 = ~l914 & l890;
assign a12108 = a2712 & ~l890;
assign a12110 = ~a12108 & ~a12106;
assign a12112 = a12110 & a5562;
assign a12114 = ~a12112 & ~a12104;
assign a12116 = ~a12114 & ~a12104;
assign a12118 = ~a12116 & ~a12098;
assign a12120 = ~a12118 & a12060;
assign a12122 = a12120 & a12004;
assign a12124 = a12122 & i332;
assign a12126 = l1260 & l1252;
assign a12128 = a12126 & l1266;
assign a12130 = ~a12128 & l1272;
assign a12132 = a12128 & ~l1272;
assign a12134 = ~a12132 & ~a12130;
assign a12136 = ~a12134 & a12124;
assign a12138 = a12124 & ~a12098;
assign a12140 = a12138 & ~a12116;
assign a12142 = ~a12124 & ~a12004;
assign a12144 = a12142 & ~a12116;
assign a12146 = ~a12124 & ~a12060;
assign a12148 = ~a12124 & ~a12098;
assign a12150 = ~a12148 & ~a12146;
assign a12152 = a12150 & ~a12138;
assign a12154 = a12152 & ~a12144;
assign a12156 = a12154 & ~a12140;
assign a12158 = a12156 & i374;
assign a12160 = ~a12158 & ~a12140;
assign a12162 = a12160 & ~a12124;
assign a12164 = a12162 & l1272;
assign a12166 = ~a12164 & ~a12136;
assign a12168 = ~a12166 & a9064;
assign a12170 = ~a12168 & ~a9066;
assign a12172 = ~a12170 & ~a9060;
assign a12174 = ~a12172 & ~a9062;
assign a12176 = ~a12174 & ~l1196;
assign a12178 = ~a12176 & ~a9028;
assign a12180 = ~a12178 & ~a9048;
assign a12182 = ~a12180 & ~a9050;
assign a12184 = ~a12182 & ~l1196;
assign a12186 = ~a12184 & ~a9028;
assign a12188 = ~a12186 & ~l886;
assign a12190 = ~a12188 & ~a5626;
assign a12192 = ~a12190 & a9026;
assign a12194 = a12190 & ~a9026;
assign a12196 = ~a12194 & ~a12192;
assign a12198 = ~a9008 & ~a8946;
assign a12200 = ~a12198 & ~a9010;
assign a12202 = ~a12200 & a9014;
assign a12204 = ~a9014 & ~a8946;
assign a12206 = ~a12204 & ~a12202;
assign a12208 = ~a8924 & l1196;
assign a12210 = a9048 & l1268;
assign a12212 = a9060 & l1268;
assign a12214 = ~a9064 & l1270;
assign a12216 = ~a12126 & l1266;
assign a12218 = a12126 & ~l1266;
assign a12220 = ~a12218 & ~a12216;
assign a12222 = ~a12220 & a12124;
assign a12224 = ~a12124 & l1266;
assign a12226 = ~a12224 & ~a12222;
assign a12228 = ~a12226 & a9064;
assign a12230 = ~a12228 & ~a12214;
assign a12232 = ~a12230 & ~a9060;
assign a12234 = ~a12232 & ~a12212;
assign a12236 = ~a12234 & ~l1196;
assign a12238 = ~a12236 & ~a12208;
assign a12240 = ~a12238 & ~a9048;
assign a12242 = ~a12240 & ~a12210;
assign a12244 = ~a12242 & ~l1196;
assign a12246 = ~a12244 & ~a12208;
assign a12248 = ~a12246 & ~l886;
assign a12250 = ~a12248 & ~a8908;
assign a12252 = a12250 & ~a12206;
assign a12254 = ~a12252 & a12196;
assign a12256 = ~a12250 & a12206;
assign a12258 = ~a12256 & a12254;
assign a12260 = ~a9006 & ~a8970;
assign a12262 = ~a12260 & ~a9008;
assign a12264 = ~a12262 & a9014;
assign a12266 = ~a9014 & ~a9006;
assign a12268 = ~a12266 & ~a12264;
assign a12270 = ~a8986 & l1196;
assign a12272 = a9048 & l1262;
assign a12274 = a9060 & l1262;
assign a12276 = ~a9064 & l1264;
assign a12278 = ~l1260 & l1252;
assign a12280 = l1260 & ~l1252;
assign a12282 = ~a12280 & ~a12278;
assign a12284 = ~a12282 & a12124;
assign a12286 = ~a12124 & l1260;
assign a12288 = ~a12286 & ~a12284;
assign a12290 = ~a12288 & a9064;
assign a12292 = ~a12290 & ~a12276;
assign a12294 = ~a12292 & ~a9060;
assign a12296 = ~a12294 & ~a12274;
assign a12298 = ~a12296 & ~l1196;
assign a12300 = ~a12298 & ~a12270;
assign a12302 = ~a12300 & ~a9048;
assign a12304 = ~a12302 & ~a12272;
assign a12306 = ~a12304 & ~l1196;
assign a12308 = ~a12306 & ~a12270;
assign a12310 = ~a12308 & ~l886;
assign a12312 = ~a12310 & ~a8972;
assign a12314 = a12312 & ~a12268;
assign a12316 = ~a12314 & a12258;
assign a12318 = ~a12312 & a12268;
assign a12320 = ~a12318 & a12316;
assign a12322 = a9014 & a8970;
assign a12324 = a8970 & a5624;
assign a12326 = ~a12324 & ~a9014;
assign a12328 = ~a12326 & ~a12322;
assign a12330 = ~a8954 & l1196;
assign a12332 = a9048 & l1254;
assign a12334 = a9060 & l1254;
assign a12336 = ~a9064 & l1258;
assign a12338 = a12124 & ~l1252;
assign a12340 = a12162 & l1252;
assign a12342 = ~a12340 & ~a12338;
assign a12344 = ~a12342 & a9064;
assign a12346 = ~a12344 & ~a12336;
assign a12348 = ~a12346 & ~a9060;
assign a12350 = ~a12348 & ~a12334;
assign a12352 = ~a12350 & ~l1196;
assign a12354 = ~a12352 & ~a12330;
assign a12356 = ~a12354 & ~a9048;
assign a12358 = ~a12356 & ~a12332;
assign a12360 = ~a12358 & ~l1196;
assign a12362 = ~a12360 & ~a12330;
assign a12364 = ~a12362 & ~l886;
assign a12366 = ~a12364 & ~a8948;
assign a12368 = a12366 & ~a12328;
assign a12370 = ~a12368 & a12320;
assign a12372 = ~a12366 & a12328;
assign a12374 = ~a12372 & a12370;
assign a12376 = ~l942 & l890;
assign a12378 = a4142 & ~l890;
assign a12380 = ~a12378 & ~a12376;
assign a12382 = ~l1502 & l890;
assign a12384 = i376 & i8;
assign a12386 = ~a5178 & i378;
assign a12388 = a12386 & ~i8;
assign a12390 = ~a12388 & ~a12384;
assign a12392 = i380 & i8;
assign a12394 = ~a5178 & i382;
assign a12396 = a12394 & ~i8;
assign a12398 = ~a12396 & ~a12392;
assign a12400 = i384 & i8;
assign a12402 = ~a5178 & i386;
assign a12404 = ~a12402 & ~a9140;
assign a12406 = ~a12404 & ~i8;
assign a12408 = ~a12406 & ~a12400;
assign a12410 = a12408 & a4746;
assign a12412 = ~a12408 & ~a4746;
assign a12414 = ~a12412 & ~a12410;
assign a12416 = i388 & i8;
assign a12418 = ~a5178 & i390;
assign a12420 = ~a12418 & ~a9122;
assign a12422 = ~a12420 & ~i8;
assign a12424 = ~a12422 & ~a12416;
assign a12426 = a12424 & a4586;
assign a12428 = ~a12424 & ~a4586;
assign a12430 = ~a12428 & ~a12426;
assign a12432 = i392 & i8;
assign a12434 = ~a5178 & i394;
assign a12436 = ~a12434 & ~a9104;
assign a12438 = ~a12436 & ~i8;
assign a12440 = ~a12438 & ~a12432;
assign a12442 = a12440 & a4426;
assign a12444 = ~a12440 & ~a4426;
assign a12446 = ~a12444 & ~a12442;
assign a12448 = i396 & i8;
assign a12450 = ~a5178 & i398;
assign a12452 = a12450 & ~i8;
assign a12454 = ~a12452 & ~a12448;
assign a12456 = i400 & i8;
assign a12458 = ~a5178 & i402;
assign a12460 = ~a12458 & ~a9086;
assign a12462 = ~a12460 & ~i8;
assign a12464 = ~a12462 & ~a12456;
assign a12466 = a12464 & a4274;
assign a12468 = i404 & i8;
assign a12470 = ~a5178 & i406;
assign a12472 = ~a12470 & ~a9078;
assign a12474 = ~a12472 & ~i8;
assign a12476 = ~a12474 & ~a12468;
assign a12478 = ~a12476 & ~a4162;
assign a12480 = ~a12464 & ~a4274;
assign a12482 = ~a12480 & ~a12478;
assign a12484 = a12482 & ~a12466;
assign a12486 = a12476 & a4162;
assign a12488 = ~a12486 & a12484;
assign a12490 = a12488 & a12454;
assign a12492 = a12490 & a12446;
assign a12494 = a12492 & a12430;
assign a12496 = a12494 & a12414;
assign a12498 = a12496 & a12398;
assign a12500 = a12498 & a12390;
assign a12502 = a12500 & a5366;
assign a12504 = a11320 & a11226;
assign a12506 = ~a11320 & i408;
assign a12508 = ~a12506 & ~a12504;
assign a12510 = a12508 & a11320;
assign a12512 = ~a12504 & ~a4122;
assign a12514 = a12512 & ~a12510;
assign a12516 = ~a12514 & ~a12502;
assign a12518 = ~a12516 & a11220;
assign a12520 = a12518 & ~a4080;
assign a12522 = ~a12520 & ~a11224;
assign a12524 = ~a12522 & ~l890;
assign a12526 = ~a12524 & ~a12382;
assign a12528 = ~a12526 & l1510;
assign a12530 = a12526 & l1514;
assign a12532 = ~a12530 & ~a12528;
assign a12534 = ~a12532 & l1494;
assign a12536 = ~l1506 & l890;
assign a12538 = a11228 & ~l890;
assign a12540 = ~a12538 & ~a12536;
assign a12542 = ~a12526 & l1542;
assign a12544 = a12526 & l1584;
assign a12546 = ~a12544 & ~a12542;
assign a12548 = ~a12546 & ~a12540;
assign a12550 = ~a12526 & l1586;
assign a12552 = a12526 & l1588;
assign a12554 = ~a12552 & ~a12550;
assign a12556 = ~a12554 & a12540;
assign a12558 = ~a12556 & ~a12548;
assign a12560 = ~a12558 & l1498;
assign a12562 = ~a12526 & l1590;
assign a12564 = a12526 & l1592;
assign a12566 = ~a12564 & ~a12562;
assign a12568 = ~a12566 & ~a12540;
assign a12570 = ~l1594 & l890;
assign a12572 = ~a12510 & ~l890;
assign a12574 = ~a12572 & ~a12570;
assign a12576 = a12574 & ~a12526;
assign a12578 = ~l1596 & l890;
assign a12580 = a12512 & ~l890;
assign a12582 = ~a12580 & ~a12578;
assign a12584 = a12582 & a12526;
assign a12586 = ~a12584 & ~a12576;
assign a12588 = ~a12586 & a12540;
assign a12590 = ~a12588 & ~a12568;
assign a12592 = ~a12590 & ~l1498;
assign a12594 = ~a12592 & ~a12560;
assign a12596 = ~a12594 & ~l1494;
assign a12598 = ~a12596 & ~a12534;
assign a12600 = a12598 & a12380;
assign a12602 = a12600 & a12374;
assign a12604 = a12602 & l998;
assign a12606 = ~l1498 & l1494;
assign a12608 = a12606 & a12540;
assign a12610 = ~a12526 & l1598;
assign a12612 = a12526 & l1600;
assign a12614 = ~a12612 & ~a12610;
assign a12616 = ~a12614 & a12608;
assign a12618 = ~a12526 & l1602;
assign a12620 = a12526 & l1604;
assign a12622 = ~a12620 & ~a12618;
assign a12624 = ~a12622 & ~a12540;
assign a12626 = ~a12526 & l1606;
assign a12628 = a12526 & l1608;
assign a12630 = ~a12628 & ~a12626;
assign a12632 = ~a12630 & a12540;
assign a12634 = ~a12632 & ~a12624;
assign a12636 = ~a12634 & l1498;
assign a12638 = ~a12526 & l1610;
assign a12640 = a12526 & l1612;
assign a12642 = ~a12640 & ~a12638;
assign a12644 = ~a12642 & ~a12540;
assign a12646 = ~a12526 & l1614;
assign a12648 = a12526 & l1616;
assign a12650 = ~a12648 & ~a12646;
assign a12652 = ~a12650 & a12540;
assign a12654 = ~a12652 & ~a12644;
assign a12656 = ~a12654 & ~l1498;
assign a12658 = ~a12656 & ~a12636;
assign a12660 = ~a12658 & ~l1494;
assign a12662 = ~a12660 & ~a12616;
assign a12664 = ~a12662 & ~a12598;
assign a12666 = ~a12526 & l1314;
assign a12668 = a12526 & l1316;
assign a12670 = ~a12668 & ~a12666;
assign a12672 = ~a12670 & a12608;
assign a12674 = ~a12526 & l1318;
assign a12676 = a12526 & l1320;
assign a12678 = ~a12676 & ~a12674;
assign a12680 = ~a12678 & ~a12540;
assign a12682 = ~a12526 & l1322;
assign a12684 = a12526 & l1324;
assign a12686 = ~a12684 & ~a12682;
assign a12688 = ~a12686 & a12540;
assign a12690 = ~a12688 & ~a12680;
assign a12692 = ~a12690 & l1498;
assign a12694 = ~a12526 & l1326;
assign a12696 = a12526 & l1328;
assign a12698 = ~a12696 & ~a12694;
assign a12700 = ~a12698 & ~a12540;
assign a12702 = ~a12526 & l1330;
assign a12704 = a12526 & l1332;
assign a12706 = ~a12704 & ~a12702;
assign a12708 = ~a12706 & a12540;
assign a12710 = ~a12708 & ~a12700;
assign a12712 = ~a12710 & ~l1498;
assign a12714 = ~a12712 & ~a12692;
assign a12716 = ~a12714 & ~l1494;
assign a12718 = ~a12716 & ~a12672;
assign a12720 = ~a12718 & a12598;
assign a12722 = ~a12720 & ~a12664;
assign a12724 = ~a12722 & ~a12602;
assign a12726 = ~a12724 & ~a12604;
assign a12728 = ~a12104 & l1278;
assign a12730 = ~a5624 & ~l886;
assign a12732 = a5868 & l1084;
assign a12734 = ~a12732 & a5880;
assign a12736 = ~a5760 & ~l972;
assign a12738 = ~a5778 & ~l1024;
assign a12740 = ~a12738 & ~a12736;
assign a12742 = a5778 & l1024;
assign a12744 = ~a12742 & ~a12740;
assign a12746 = ~a5796 & ~l1092;
assign a12748 = ~a12746 & ~a12744;
assign a12750 = a5796 & l1092;
assign a12752 = ~a12750 & ~a12748;
assign a12754 = ~a5814 & ~l1090;
assign a12756 = ~a12754 & ~a12752;
assign a12758 = a5814 & l1090;
assign a12760 = ~a12758 & ~a12756;
assign a12762 = ~a5832 & ~l1088;
assign a12764 = ~a12762 & ~a12760;
assign a12766 = a5832 & l1088;
assign a12768 = ~a12766 & ~a12764;
assign a12770 = ~a5850 & ~l1086;
assign a12772 = ~a12770 & ~a12768;
assign a12774 = a5850 & l1086;
assign a12776 = ~a12774 & ~a12772;
assign a12778 = ~a5868 & ~l1084;
assign a12780 = ~a12778 & ~a12776;
assign a12782 = ~a12780 & a12734;
assign a12784 = a5760 & l972;
assign a12786 = ~a12784 & ~a12742;
assign a12788 = ~a12786 & ~a12738;
assign a12790 = ~a12788 & ~a12750;
assign a12792 = ~a12790 & ~a12746;
assign a12794 = ~a12792 & ~a12758;
assign a12796 = ~a12794 & ~a12754;
assign a12798 = ~a12796 & ~a12766;
assign a12800 = ~a12798 & ~a12762;
assign a12802 = ~a12800 & ~a12774;
assign a12804 = ~a12802 & ~a12770;
assign a12806 = ~a12804 & ~a12732;
assign a12808 = ~a12806 & ~a12778;
assign a12810 = a12808 & ~a5880;
assign a12812 = ~a12810 & ~a12782;
assign a12814 = ~a12812 & a12730;
assign a12816 = a12814 & ~l1060;
assign a12818 = ~a12814 & ~a5874;
assign a12820 = ~a12818 & ~a12816;
assign a12822 = ~a12820 & a12104;
assign a12824 = ~a12822 & ~a12728;
assign a12826 = a12824 & ~a12726;
assign a12828 = ~a12824 & a12726;
assign a12830 = ~a12828 & ~a12826;
assign a12832 = ~l1474 & l890;
assign a12834 = a11584 & ~l890;
assign a12836 = ~a12834 & ~a12832;
assign a12838 = a12836 & a12602;
assign a12840 = ~a12526 & l1618;
assign a12842 = a12526 & l1620;
assign a12844 = ~a12842 & ~a12840;
assign a12846 = ~a12844 & a12608;
assign a12848 = ~a12526 & l1622;
assign a12850 = a12526 & l1624;
assign a12852 = ~a12850 & ~a12848;
assign a12854 = ~a12852 & ~a12540;
assign a12856 = ~a12526 & l1626;
assign a12858 = a12526 & l1628;
assign a12860 = ~a12858 & ~a12856;
assign a12862 = ~a12860 & a12540;
assign a12864 = ~a12862 & ~a12854;
assign a12866 = ~a12864 & l1498;
assign a12868 = ~a12526 & l1630;
assign a12870 = a12526 & l1632;
assign a12872 = ~a12870 & ~a12868;
assign a12874 = ~a12872 & ~a12540;
assign a12876 = ~l1634 & l890;
assign a12878 = a11320 & a4138;
assign a12880 = ~a11320 & i428;
assign a12882 = ~a12880 & ~a12878;
assign a12884 = a12882 & a12510;
assign a12886 = a12884 & ~l890;
assign a12888 = ~a12886 & ~a12876;
assign a12890 = ~a12888 & ~a12526;
assign a12892 = ~l1636 & l890;
assign a12894 = a12882 & a12504;
assign a12896 = ~a12504 & a4162;
assign a12898 = ~a12896 & ~a12894;
assign a12900 = ~a12898 & ~l890;
assign a12902 = ~a12900 & ~a12892;
assign a12904 = ~a12902 & a12526;
assign a12906 = ~a12904 & ~a12890;
assign a12908 = ~a12906 & a12540;
assign a12910 = ~a12908 & ~a12874;
assign a12912 = ~a12910 & ~l1498;
assign a12914 = ~a12912 & ~a12866;
assign a12916 = ~a12914 & ~l1494;
assign a12918 = ~a12916 & ~a12846;
assign a12920 = ~a12918 & ~a12598;
assign a12922 = ~a12526 & l1334;
assign a12924 = a12526 & l1336;
assign a12926 = ~a12924 & ~a12922;
assign a12928 = ~a12926 & a12608;
assign a12930 = ~a12526 & l1338;
assign a12932 = a12526 & l1340;
assign a12934 = ~a12932 & ~a12930;
assign a12936 = ~a12934 & ~a12540;
assign a12938 = ~a12526 & l1342;
assign a12940 = a12526 & l1344;
assign a12942 = ~a12940 & ~a12938;
assign a12944 = ~a12942 & a12540;
assign a12946 = ~a12944 & ~a12936;
assign a12948 = ~a12946 & l1498;
assign a12950 = ~l1346 & l890;
assign a12952 = a11252 & ~l890;
assign a12954 = ~a12952 & ~a12950;
assign a12956 = ~a12954 & ~a12526;
assign a12958 = ~l1348 & l890;
assign a12960 = ~a11264 & ~l890;
assign a12962 = ~a12960 & ~a12958;
assign a12964 = ~a12962 & a12526;
assign a12966 = ~a12964 & ~a12956;
assign a12968 = ~a12966 & ~a12540;
assign a12970 = ~l1350 & l890;
assign a12972 = ~a11274 & ~l890;
assign a12974 = ~a12972 & ~a12970;
assign a12976 = ~a12974 & ~a12526;
assign a12978 = a12526 & l1352;
assign a12980 = ~a12978 & ~a12976;
assign a12982 = ~a12980 & a12540;
assign a12984 = ~a12982 & ~a12968;
assign a12986 = ~a12984 & ~l1498;
assign a12988 = ~a12986 & ~a12948;
assign a12990 = ~a12988 & ~l1494;
assign a12992 = ~a12990 & ~a12928;
assign a12994 = ~a12992 & a12598;
assign a12996 = ~a12994 & ~a12920;
assign a12998 = ~a12996 & ~a12602;
assign a13000 = ~a12998 & ~a12838;
assign a13002 = ~a12104 & ~a10652;
assign a13004 = a12814 & l972;
assign a13006 = ~a12814 & ~a5760;
assign a13008 = ~a13006 & ~a13004;
assign a13010 = ~a13008 & a12104;
assign a13012 = ~a13010 & ~a13002;
assign a13014 = ~a13012 & a13000;
assign a13016 = ~l1476 & l890;
assign a13018 = a11638 & ~l890;
assign a13020 = ~a13018 & ~a13016;
assign a13022 = a13020 & a12602;
assign a13024 = ~a12526 & l1638;
assign a13026 = a12526 & l1640;
assign a13028 = ~a13026 & ~a13024;
assign a13030 = ~a13028 & a12608;
assign a13032 = ~a12526 & l1642;
assign a13034 = a12526 & l1644;
assign a13036 = ~a13034 & ~a13032;
assign a13038 = ~a13036 & ~a12540;
assign a13040 = ~a12526 & l1646;
assign a13042 = a12526 & l1648;
assign a13044 = ~a13042 & ~a13040;
assign a13046 = ~a13044 & a12540;
assign a13048 = ~a13046 & ~a13038;
assign a13050 = ~a13048 & l1498;
assign a13052 = ~a12526 & l1650;
assign a13054 = a12526 & l1652;
assign a13056 = ~a13054 & ~a13052;
assign a13058 = ~a13056 & ~a12540;
assign a13060 = ~l1654 & l890;
assign a13062 = a11320 & a4264;
assign a13064 = ~a11320 & i432;
assign a13066 = ~a13064 & ~a13062;
assign a13068 = a13066 & a12510;
assign a13070 = a13068 & ~l890;
assign a13072 = ~a13070 & ~a13060;
assign a13074 = ~a13072 & ~a12526;
assign a13076 = ~l1656 & l890;
assign a13078 = a13066 & a12504;
assign a13080 = ~a12504 & a4274;
assign a13082 = ~a13080 & ~a13078;
assign a13084 = ~a13082 & ~l890;
assign a13086 = ~a13084 & ~a13076;
assign a13088 = ~a13086 & a12526;
assign a13090 = ~a13088 & ~a13074;
assign a13092 = ~a13090 & a12540;
assign a13094 = ~a13092 & ~a13058;
assign a13096 = ~a13094 & ~l1498;
assign a13098 = ~a13096 & ~a13050;
assign a13100 = ~a13098 & ~l1494;
assign a13102 = ~a13100 & ~a13030;
assign a13104 = ~a13102 & ~a12598;
assign a13106 = ~a12526 & l1354;
assign a13108 = a12526 & l1356;
assign a13110 = ~a13108 & ~a13106;
assign a13112 = ~a13110 & a12608;
assign a13114 = ~a12526 & l1358;
assign a13116 = a12526 & l1360;
assign a13118 = ~a13116 & ~a13114;
assign a13120 = ~a13118 & ~a12540;
assign a13122 = ~a12526 & l1362;
assign a13124 = a12526 & l1364;
assign a13126 = ~a13124 & ~a13122;
assign a13128 = ~a13126 & a12540;
assign a13130 = ~a13128 & ~a13120;
assign a13132 = ~a13130 & l1498;
assign a13134 = ~l1366 & l890;
assign a13136 = a11332 & ~l890;
assign a13138 = ~a13136 & ~a13134;
assign a13140 = ~a13138 & ~a12526;
assign a13142 = ~l1368 & l890;
assign a13144 = ~a11338 & ~l890;
assign a13146 = ~a13144 & ~a13142;
assign a13148 = ~a13146 & a12526;
assign a13150 = ~a13148 & ~a13140;
assign a13152 = ~a13150 & ~a12540;
assign a13154 = ~l1370 & l890;
assign a13156 = ~a11348 & ~l890;
assign a13158 = ~a13156 & ~a13154;
assign a13160 = ~a13158 & ~a12526;
assign a13162 = a12526 & l1372;
assign a13164 = ~a13162 & ~a13160;
assign a13166 = ~a13164 & a12540;
assign a13168 = ~a13166 & ~a13152;
assign a13170 = ~a13168 & ~l1498;
assign a13172 = ~a13170 & ~a13132;
assign a13174 = ~a13172 & ~l1494;
assign a13176 = ~a13174 & ~a13112;
assign a13178 = ~a13176 & a12598;
assign a13180 = ~a13178 & ~a13104;
assign a13182 = ~a13180 & ~a12602;
assign a13184 = ~a13182 & ~a13022;
assign a13186 = ~a12104 & ~a10592;
assign a13188 = a12814 & l1024;
assign a13190 = ~a12814 & ~a5778;
assign a13192 = ~a13190 & ~a13188;
assign a13194 = ~a13192 & a12104;
assign a13196 = ~a13194 & ~a13186;
assign a13198 = ~a13196 & a13184;
assign a13200 = ~a13198 & ~a13014;
assign a13202 = a13196 & ~a13184;
assign a13204 = ~a13202 & ~a13200;
assign a13206 = ~l1478 & l890;
assign a13208 = a11710 & ~l890;
assign a13210 = ~a13208 & ~a13206;
assign a13212 = a13210 & a12602;
assign a13214 = ~a12526 & l1658;
assign a13216 = a12526 & l1660;
assign a13218 = ~a13216 & ~a13214;
assign a13220 = ~a13218 & a12608;
assign a13222 = ~a12526 & l1662;
assign a13224 = a12526 & l1664;
assign a13226 = ~a13224 & ~a13222;
assign a13228 = ~a13226 & ~a12540;
assign a13230 = ~a12526 & l1666;
assign a13232 = a12526 & l1668;
assign a13234 = ~a13232 & ~a13230;
assign a13236 = ~a13234 & a12540;
assign a13238 = ~a13236 & ~a13228;
assign a13240 = ~a13238 & l1498;
assign a13242 = ~a12526 & l1670;
assign a13244 = a12526 & l1672;
assign a13246 = ~a13244 & ~a13242;
assign a13248 = ~a13246 & ~a12540;
assign a13250 = ~l1674 & l890;
assign a13252 = a11320 & a4416;
assign a13254 = ~a11320 & i436;
assign a13256 = ~a13254 & ~a13252;
assign a13258 = a13256 & a12510;
assign a13260 = a13258 & ~l890;
assign a13262 = ~a13260 & ~a13250;
assign a13264 = ~a13262 & ~a12526;
assign a13266 = ~l1676 & l890;
assign a13268 = a13256 & a12504;
assign a13270 = ~a12504 & a4426;
assign a13272 = ~a13270 & ~a13268;
assign a13274 = ~a13272 & ~l890;
assign a13276 = ~a13274 & ~a13266;
assign a13278 = ~a13276 & a12526;
assign a13280 = ~a13278 & ~a13264;
assign a13282 = ~a13280 & a12540;
assign a13284 = ~a13282 & ~a13248;
assign a13286 = ~a13284 & ~l1498;
assign a13288 = ~a13286 & ~a13240;
assign a13290 = ~a13288 & ~l1494;
assign a13292 = ~a13290 & ~a13220;
assign a13294 = ~a13292 & ~a12598;
assign a13296 = ~a12526 & l1374;
assign a13298 = a12526 & l1376;
assign a13300 = ~a13298 & ~a13296;
assign a13302 = ~a13300 & a12608;
assign a13304 = ~a12526 & l1378;
assign a13306 = a12526 & l1380;
assign a13308 = ~a13306 & ~a13304;
assign a13310 = ~a13308 & ~a12540;
assign a13312 = ~a12526 & l1382;
assign a13314 = a12526 & l1384;
assign a13316 = ~a13314 & ~a13312;
assign a13318 = ~a13316 & a12540;
assign a13320 = ~a13318 & ~a13310;
assign a13322 = ~a13320 & l1498;
assign a13324 = ~l1386 & l890;
assign a13326 = a11374 & ~l890;
assign a13328 = ~a13326 & ~a13324;
assign a13330 = ~a13328 & ~a12526;
assign a13332 = ~l1388 & l890;
assign a13334 = ~a11380 & ~l890;
assign a13336 = ~a13334 & ~a13332;
assign a13338 = ~a13336 & a12526;
assign a13340 = ~a13338 & ~a13330;
assign a13342 = ~a13340 & ~a12540;
assign a13344 = ~l1390 & l890;
assign a13346 = ~a11390 & ~l890;
assign a13348 = ~a13346 & ~a13344;
assign a13350 = ~a13348 & ~a12526;
assign a13352 = a12526 & l1392;
assign a13354 = ~a13352 & ~a13350;
assign a13356 = ~a13354 & a12540;
assign a13358 = ~a13356 & ~a13342;
assign a13360 = ~a13358 & ~l1498;
assign a13362 = ~a13360 & ~a13322;
assign a13364 = ~a13362 & ~l1494;
assign a13366 = ~a13364 & ~a13302;
assign a13368 = ~a13366 & a12598;
assign a13370 = ~a13368 & ~a13294;
assign a13372 = ~a13370 & ~a12602;
assign a13374 = ~a13372 & ~a13212;
assign a13376 = ~a12104 & ~a10556;
assign a13378 = a12814 & l1092;
assign a13380 = ~a12814 & ~a5796;
assign a13382 = ~a13380 & ~a13378;
assign a13384 = ~a13382 & a12104;
assign a13386 = ~a13384 & ~a13376;
assign a13388 = ~a13386 & a13374;
assign a13390 = ~a13388 & ~a13204;
assign a13392 = a13386 & ~a13374;
assign a13394 = ~a13392 & ~a13390;
assign a13396 = ~l1480 & l890;
assign a13398 = a11782 & ~l890;
assign a13400 = ~a13398 & ~a13396;
assign a13402 = a13400 & a12602;
assign a13404 = ~a12526 & l1678;
assign a13406 = a12526 & l1680;
assign a13408 = ~a13406 & ~a13404;
assign a13410 = ~a13408 & a12608;
assign a13412 = ~a12526 & l1682;
assign a13414 = a12526 & l1684;
assign a13416 = ~a13414 & ~a13412;
assign a13418 = ~a13416 & ~a12540;
assign a13420 = ~a12526 & l1686;
assign a13422 = a12526 & l1688;
assign a13424 = ~a13422 & ~a13420;
assign a13426 = ~a13424 & a12540;
assign a13428 = ~a13426 & ~a13418;
assign a13430 = ~a13428 & l1498;
assign a13432 = ~a12526 & l1690;
assign a13434 = a12526 & l1692;
assign a13436 = ~a13434 & ~a13432;
assign a13438 = ~a13436 & ~a12540;
assign a13440 = ~l1694 & l890;
assign a13442 = a11320 & a4576;
assign a13444 = ~a11320 & i440;
assign a13446 = ~a13444 & ~a13442;
assign a13448 = a13446 & a12510;
assign a13450 = a13448 & ~l890;
assign a13452 = ~a13450 & ~a13440;
assign a13454 = ~a13452 & ~a12526;
assign a13456 = ~l1696 & l890;
assign a13458 = a13446 & a12504;
assign a13460 = ~a12504 & a4586;
assign a13462 = ~a13460 & ~a13458;
assign a13464 = ~a13462 & ~l890;
assign a13466 = ~a13464 & ~a13456;
assign a13468 = ~a13466 & a12526;
assign a13470 = ~a13468 & ~a13454;
assign a13472 = ~a13470 & a12540;
assign a13474 = ~a13472 & ~a13438;
assign a13476 = ~a13474 & ~l1498;
assign a13478 = ~a13476 & ~a13430;
assign a13480 = ~a13478 & ~l1494;
assign a13482 = ~a13480 & ~a13410;
assign a13484 = ~a13482 & ~a12598;
assign a13486 = ~a12526 & l1394;
assign a13488 = a12526 & l1396;
assign a13490 = ~a13488 & ~a13486;
assign a13492 = ~a13490 & a12608;
assign a13494 = ~a12526 & l1398;
assign a13496 = a12526 & l1400;
assign a13498 = ~a13496 & ~a13494;
assign a13500 = ~a13498 & ~a12540;
assign a13502 = ~a12526 & l1402;
assign a13504 = a12526 & l1404;
assign a13506 = ~a13504 & ~a13502;
assign a13508 = ~a13506 & a12540;
assign a13510 = ~a13508 & ~a13500;
assign a13512 = ~a13510 & l1498;
assign a13514 = ~l1406 & l890;
assign a13516 = a11416 & ~l890;
assign a13518 = ~a13516 & ~a13514;
assign a13520 = ~a13518 & ~a12526;
assign a13522 = ~l1408 & l890;
assign a13524 = ~a11422 & ~l890;
assign a13526 = ~a13524 & ~a13522;
assign a13528 = ~a13526 & a12526;
assign a13530 = ~a13528 & ~a13520;
assign a13532 = ~a13530 & ~a12540;
assign a13534 = ~l1410 & l890;
assign a13536 = ~a11432 & ~l890;
assign a13538 = ~a13536 & ~a13534;
assign a13540 = ~a13538 & ~a12526;
assign a13542 = a12526 & l1412;
assign a13544 = ~a13542 & ~a13540;
assign a13546 = ~a13544 & a12540;
assign a13548 = ~a13546 & ~a13532;
assign a13550 = ~a13548 & ~l1498;
assign a13552 = ~a13550 & ~a13512;
assign a13554 = ~a13552 & ~l1494;
assign a13556 = ~a13554 & ~a13492;
assign a13558 = ~a13556 & a12598;
assign a13560 = ~a13558 & ~a13484;
assign a13562 = ~a13560 & ~a12602;
assign a13564 = ~a13562 & ~a13402;
assign a13566 = ~a12104 & ~a10520;
assign a13568 = a12814 & l1090;
assign a13570 = ~a12814 & ~a5814;
assign a13572 = ~a13570 & ~a13568;
assign a13574 = ~a13572 & a12104;
assign a13576 = ~a13574 & ~a13566;
assign a13578 = ~a13576 & a13564;
assign a13580 = ~a13578 & ~a13394;
assign a13582 = a13576 & ~a13564;
assign a13584 = ~a13582 & ~a13580;
assign a13586 = ~l1482 & l890;
assign a13588 = a11854 & ~l890;
assign a13590 = ~a13588 & ~a13586;
assign a13592 = a13590 & a12602;
assign a13594 = ~a12526 & l1698;
assign a13596 = a12526 & l1700;
assign a13598 = ~a13596 & ~a13594;
assign a13600 = ~a13598 & a12608;
assign a13602 = ~a12526 & l1702;
assign a13604 = a12526 & l1704;
assign a13606 = ~a13604 & ~a13602;
assign a13608 = ~a13606 & ~a12540;
assign a13610 = ~a12526 & l1706;
assign a13612 = a12526 & l1708;
assign a13614 = ~a13612 & ~a13610;
assign a13616 = ~a13614 & a12540;
assign a13618 = ~a13616 & ~a13608;
assign a13620 = ~a13618 & l1498;
assign a13622 = ~a12526 & l1710;
assign a13624 = a12526 & l1712;
assign a13626 = ~a13624 & ~a13622;
assign a13628 = ~a13626 & ~a12540;
assign a13630 = ~l1714 & l890;
assign a13632 = a11320 & a4736;
assign a13634 = ~a11320 & i444;
assign a13636 = ~a13634 & ~a13632;
assign a13638 = a13636 & a12510;
assign a13640 = a13638 & ~l890;
assign a13642 = ~a13640 & ~a13630;
assign a13644 = ~a13642 & ~a12526;
assign a13646 = ~l1716 & l890;
assign a13648 = a13636 & a12504;
assign a13650 = ~a12504 & a4746;
assign a13652 = ~a13650 & ~a13648;
assign a13654 = ~a13652 & ~l890;
assign a13656 = ~a13654 & ~a13646;
assign a13658 = ~a13656 & a12526;
assign a13660 = ~a13658 & ~a13644;
assign a13662 = ~a13660 & a12540;
assign a13664 = ~a13662 & ~a13628;
assign a13666 = ~a13664 & ~l1498;
assign a13668 = ~a13666 & ~a13620;
assign a13670 = ~a13668 & ~l1494;
assign a13672 = ~a13670 & ~a13600;
assign a13674 = ~a13672 & ~a12598;
assign a13676 = ~a12526 & l1414;
assign a13678 = a12526 & l1416;
assign a13680 = ~a13678 & ~a13676;
assign a13682 = ~a13680 & a12608;
assign a13684 = ~a12526 & l1418;
assign a13686 = a12526 & l1420;
assign a13688 = ~a13686 & ~a13684;
assign a13690 = ~a13688 & ~a12540;
assign a13692 = ~a12526 & l1422;
assign a13694 = a12526 & l1424;
assign a13696 = ~a13694 & ~a13692;
assign a13698 = ~a13696 & a12540;
assign a13700 = ~a13698 & ~a13690;
assign a13702 = ~a13700 & l1498;
assign a13704 = ~l1426 & l890;
assign a13706 = a11458 & ~l890;
assign a13708 = ~a13706 & ~a13704;
assign a13710 = ~a13708 & ~a12526;
assign a13712 = ~l1428 & l890;
assign a13714 = ~a11464 & ~l890;
assign a13716 = ~a13714 & ~a13712;
assign a13718 = ~a13716 & a12526;
assign a13720 = ~a13718 & ~a13710;
assign a13722 = ~a13720 & ~a12540;
assign a13724 = ~l1430 & l890;
assign a13726 = ~a11474 & ~l890;
assign a13728 = ~a13726 & ~a13724;
assign a13730 = ~a13728 & ~a12526;
assign a13732 = a12526 & l1432;
assign a13734 = ~a13732 & ~a13730;
assign a13736 = ~a13734 & a12540;
assign a13738 = ~a13736 & ~a13722;
assign a13740 = ~a13738 & ~l1498;
assign a13742 = ~a13740 & ~a13702;
assign a13744 = ~a13742 & ~l1494;
assign a13746 = ~a13744 & ~a13682;
assign a13748 = ~a13746 & a12598;
assign a13750 = ~a13748 & ~a13674;
assign a13752 = ~a13750 & ~a12602;
assign a13754 = ~a13752 & ~a13592;
assign a13756 = ~a12104 & ~a10484;
assign a13758 = a12814 & l1088;
assign a13760 = ~a12814 & ~a5832;
assign a13762 = ~a13760 & ~a13758;
assign a13764 = ~a13762 & a12104;
assign a13766 = ~a13764 & ~a13756;
assign a13768 = ~a13766 & a13754;
assign a13770 = ~a13768 & ~a13584;
assign a13772 = a13766 & ~a13754;
assign a13774 = ~a13772 & ~a13770;
assign a13776 = ~l1484 & l890;
assign a13778 = a11926 & ~l890;
assign a13780 = ~a13778 & ~a13776;
assign a13782 = a13780 & a12602;
assign a13784 = ~a12526 & l1718;
assign a13786 = a12526 & l1720;
assign a13788 = ~a13786 & ~a13784;
assign a13790 = ~a13788 & a12608;
assign a13792 = ~a12526 & l1722;
assign a13794 = a12526 & l1724;
assign a13796 = ~a13794 & ~a13792;
assign a13798 = ~a13796 & ~a12540;
assign a13800 = ~a12526 & l1726;
assign a13802 = a12526 & l1728;
assign a13804 = ~a13802 & ~a13800;
assign a13806 = ~a13804 & a12540;
assign a13808 = ~a13806 & ~a13798;
assign a13810 = ~a13808 & l1498;
assign a13812 = ~a12526 & l1730;
assign a13814 = a12526 & l1732;
assign a13816 = ~a13814 & ~a13812;
assign a13818 = ~a13816 & ~a12540;
assign a13820 = ~l1734 & l890;
assign a13822 = a11320 & a4884;
assign a13824 = ~a11320 & i448;
assign a13826 = ~a13824 & ~a13822;
assign a13828 = a13826 & a12510;
assign a13830 = a13828 & ~l890;
assign a13832 = ~a13830 & ~a13820;
assign a13834 = ~a13832 & ~a12526;
assign a13836 = a12526 & l1736;
assign a13838 = ~a13836 & ~a13834;
assign a13840 = ~a13838 & a12540;
assign a13842 = ~a13840 & ~a13818;
assign a13844 = ~a13842 & ~l1498;
assign a13846 = ~a13844 & ~a13810;
assign a13848 = ~a13846 & ~l1494;
assign a13850 = ~a13848 & ~a13790;
assign a13852 = ~a13850 & ~a12598;
assign a13854 = ~a12526 & l1434;
assign a13856 = a12526 & l1436;
assign a13858 = ~a13856 & ~a13854;
assign a13860 = ~a13858 & a12608;
assign a13862 = ~a12526 & l1438;
assign a13864 = a12526 & l1440;
assign a13866 = ~a13864 & ~a13862;
assign a13868 = ~a13866 & ~a12540;
assign a13870 = ~a12526 & l1442;
assign a13872 = a12526 & l1444;
assign a13874 = ~a13872 & ~a13870;
assign a13876 = ~a13874 & a12540;
assign a13878 = ~a13876 & ~a13868;
assign a13880 = ~a13878 & l1498;
assign a13882 = ~l1446 & l890;
assign a13884 = a11500 & ~l890;
assign a13886 = ~a13884 & ~a13882;
assign a13888 = ~a13886 & ~a12526;
assign a13890 = ~l1448 & l890;
assign a13892 = ~a11506 & ~l890;
assign a13894 = ~a13892 & ~a13890;
assign a13896 = ~a13894 & a12526;
assign a13898 = ~a13896 & ~a13888;
assign a13900 = ~a13898 & ~a12540;
assign a13902 = ~l1450 & l890;
assign a13904 = ~a11516 & ~l890;
assign a13906 = ~a13904 & ~a13902;
assign a13908 = ~a13906 & ~a12526;
assign a13910 = a12526 & l1452;
assign a13912 = ~a13910 & ~a13908;
assign a13914 = ~a13912 & a12540;
assign a13916 = ~a13914 & ~a13900;
assign a13918 = ~a13916 & ~l1498;
assign a13920 = ~a13918 & ~a13880;
assign a13922 = ~a13920 & ~l1494;
assign a13924 = ~a13922 & ~a13860;
assign a13926 = ~a13924 & a12598;
assign a13928 = ~a13926 & ~a13852;
assign a13930 = ~a13928 & ~a12602;
assign a13932 = ~a13930 & ~a13782;
assign a13934 = ~a12104 & ~a9072;
assign a13936 = a12814 & l1086;
assign a13938 = ~a12814 & ~a5850;
assign a13940 = ~a13938 & ~a13936;
assign a13942 = ~a13940 & a12104;
assign a13944 = ~a13942 & ~a13934;
assign a13946 = ~a13944 & a13932;
assign a13948 = ~a13946 & ~a13774;
assign a13950 = a13944 & ~a13932;
assign a13952 = ~a13950 & ~a13948;
assign a13954 = ~l940 & l890;
assign a13956 = ~a11952 & ~l890;
assign a13958 = ~a13956 & ~a13954;
assign a13960 = ~a13958 & a12602;
assign a13962 = ~a12526 & l1738;
assign a13964 = a12526 & l1740;
assign a13966 = ~a13964 & ~a13962;
assign a13968 = ~a13966 & a12608;
assign a13970 = ~a12526 & l1742;
assign a13972 = a12526 & l1744;
assign a13974 = ~a13972 & ~a13970;
assign a13976 = ~a13974 & ~a12540;
assign a13978 = ~a12526 & l1746;
assign a13980 = a12526 & l1748;
assign a13982 = ~a13980 & ~a13978;
assign a13984 = ~a13982 & a12540;
assign a13986 = ~a13984 & ~a13976;
assign a13988 = ~a13986 & l1498;
assign a13990 = ~a12526 & l1750;
assign a13992 = a12526 & l1752;
assign a13994 = ~a13992 & ~a13990;
assign a13996 = ~a13994 & ~a12540;
assign a13998 = ~a12526 & l1754;
assign a14000 = a12526 & l1756;
assign a14002 = ~a14000 & ~a13998;
assign a14004 = ~a14002 & a12540;
assign a14006 = ~a14004 & ~a13996;
assign a14008 = ~a14006 & ~l1498;
assign a14010 = ~a14008 & ~a13988;
assign a14012 = ~a14010 & ~l1494;
assign a14014 = ~a14012 & ~a13968;
assign a14016 = ~a14014 & ~a12598;
assign a14018 = ~a12526 & l1454;
assign a14020 = a12526 & l1456;
assign a14022 = ~a14020 & ~a14018;
assign a14024 = ~a14022 & a12608;
assign a14026 = ~a12526 & l1458;
assign a14028 = a12526 & l1460;
assign a14030 = ~a14028 & ~a14026;
assign a14032 = ~a14030 & ~a12540;
assign a14034 = ~a12526 & l1462;
assign a14036 = a12526 & l1464;
assign a14038 = ~a14036 & ~a14034;
assign a14040 = ~a14038 & a12540;
assign a14042 = ~a14040 & ~a14032;
assign a14044 = ~a14042 & l1498;
assign a14046 = ~l1466 & l890;
assign a14048 = a11542 & ~l890;
assign a14050 = ~a14048 & ~a14046;
assign a14052 = ~a14050 & ~a12526;
assign a14054 = ~l1468 & l890;
assign a14056 = ~a11548 & ~l890;
assign a14058 = ~a14056 & ~a14054;
assign a14060 = ~a14058 & a12526;
assign a14062 = ~a14060 & ~a14052;
assign a14064 = ~a14062 & ~a12540;
assign a14066 = ~a12526 & l1470;
assign a14068 = a12526 & l1472;
assign a14070 = ~a14068 & ~a14066;
assign a14072 = ~a14070 & a12540;
assign a14074 = ~a14072 & ~a14064;
assign a14076 = ~a14074 & ~l1498;
assign a14078 = ~a14076 & ~a14044;
assign a14080 = ~a14078 & ~l1494;
assign a14082 = ~a14080 & ~a14024;
assign a14084 = ~a14082 & a12598;
assign a14086 = ~a14084 & ~a14016;
assign a14088 = ~a14086 & ~a12602;
assign a14090 = ~a14088 & ~a13960;
assign a14092 = ~a12104 & l1280;
assign a14094 = a12814 & l1084;
assign a14096 = ~a12814 & ~a5868;
assign a14098 = ~a14096 & ~a14094;
assign a14100 = ~a14098 & a12104;
assign a14102 = ~a14100 & ~a14092;
assign a14104 = ~a14102 & a14090;
assign a14106 = ~a14104 & ~a13952;
assign a14108 = a14102 & ~a14090;
assign a14110 = ~a14108 & ~a14106;
assign a14112 = a14110 & a12830;
assign a14114 = ~a14110 & ~a12830;
assign a14116 = ~a14114 & ~a14112;
assign a14118 = ~a14116 & ~a12726;
assign a14120 = a13196 & a13012;
assign a14122 = a14120 & a13386;
assign a14124 = a14122 & a13576;
assign a14126 = a14124 & a13766;
assign a14128 = a14126 & a13944;
assign a14130 = a14128 & a14102;
assign a14132 = ~a14130 & ~a12824;
assign a14134 = a14130 & a12824;
assign a14136 = ~a14134 & ~a14132;
assign a14138 = ~a14136 & a14116;
assign a14140 = ~a14138 & ~a14118;
assign a14142 = a14140 & l992;
assign a14144 = ~a14140 & ~l992;
assign a14146 = ~a14144 & ~a14142;
assign a14148 = a14116 & a13012;
assign a14150 = ~a14148 & ~a10646;
assign a14152 = ~a14116 & ~a13000;
assign a14154 = ~a14152 & a14150;
assign a14156 = ~a14116 & ~a13184;
assign a14158 = ~a13196 & ~a13012;
assign a14160 = ~a14158 & ~a14120;
assign a14162 = ~a14160 & a14116;
assign a14164 = ~a14162 & ~a14156;
assign a14166 = a14164 & ~a10622;
assign a14168 = ~a14166 & ~a14154;
assign a14170 = ~a14164 & a10622;
assign a14172 = ~a14170 & ~a14168;
assign a14174 = ~a14116 & ~a13374;
assign a14176 = ~a14120 & ~a13386;
assign a14178 = ~a14176 & ~a14122;
assign a14180 = ~a14178 & a14116;
assign a14182 = ~a14180 & ~a14174;
assign a14184 = a14182 & ~a10586;
assign a14186 = ~a14184 & ~a14172;
assign a14188 = ~a14182 & a10586;
assign a14190 = ~a14188 & ~a14186;
assign a14192 = ~a14116 & ~a13564;
assign a14194 = ~a14122 & ~a13576;
assign a14196 = ~a14194 & ~a14124;
assign a14198 = ~a14196 & a14116;
assign a14200 = ~a14198 & ~a14192;
assign a14202 = a14200 & ~a10550;
assign a14204 = ~a14202 & ~a14190;
assign a14206 = ~a14200 & a10550;
assign a14208 = ~a14206 & ~a14204;
assign a14210 = ~a14116 & ~a13754;
assign a14212 = ~a14124 & ~a13766;
assign a14214 = ~a14212 & ~a14126;
assign a14216 = ~a14214 & a14116;
assign a14218 = ~a14216 & ~a14210;
assign a14220 = a14218 & ~a10514;
assign a14222 = ~a14220 & ~a14208;
assign a14224 = ~a14218 & a10514;
assign a14226 = ~a14224 & ~a14222;
assign a14228 = ~a14116 & ~a13932;
assign a14230 = ~a14126 & ~a13944;
assign a14232 = ~a14230 & ~a14128;
assign a14234 = ~a14232 & a14116;
assign a14236 = ~a14234 & ~a14228;
assign a14238 = a14236 & ~a10478;
assign a14240 = ~a14238 & ~a14226;
assign a14242 = ~a14236 & a10478;
assign a14244 = ~a14242 & ~a14240;
assign a14246 = ~a14116 & ~a14090;
assign a14248 = ~a14128 & ~a14102;
assign a14250 = ~a14248 & ~a14130;
assign a14252 = ~a14250 & a14116;
assign a14254 = ~a14252 & ~a14246;
assign a14256 = a14254 & l1140;
assign a14258 = ~a14256 & ~a14244;
assign a14260 = ~a14254 & ~l1140;
assign a14262 = ~a14260 & ~a14258;
assign a14264 = ~a14262 & a14146;
assign a14266 = a14262 & ~a14146;
assign a14268 = ~a14266 & ~a14264;
assign a14270 = ~a14268 & ~l908;
assign a14272 = ~l994 & l992;
assign a14274 = l994 & ~l992;
assign a14276 = ~a14274 & ~a14272;
assign a14278 = l1142 & ~l1140;
assign a14280 = ~a14278 & a14276;
assign a14282 = ~l1142 & l1140;
assign a14284 = ~a14282 & a14280;
assign a14286 = a10478 & l1134;
assign a14288 = ~a14286 & a14284;
assign a14290 = ~a10478 & ~l1134;
assign a14292 = ~a14290 & a14288;
assign a14294 = ~l1126 & l890;
assign a14296 = a9140 & ~l890;
assign a14298 = ~a14296 & ~a14294;
assign a14300 = ~a14298 & a10514;
assign a14302 = ~a14300 & a14292;
assign a14304 = a14298 & ~a10514;
assign a14306 = ~a14304 & a14302;
assign a14308 = ~l1118 & l890;
assign a14310 = a9122 & ~l890;
assign a14312 = ~a14310 & ~a14308;
assign a14314 = ~a14312 & a10550;
assign a14316 = ~a14314 & a14306;
assign a14318 = a14312 & ~a10550;
assign a14320 = ~a14318 & a14316;
assign a14322 = ~l1110 & l890;
assign a14324 = a9104 & ~l890;
assign a14326 = ~a14324 & ~a14322;
assign a14328 = ~a14326 & a10586;
assign a14330 = ~a14328 & a14320;
assign a14332 = a14326 & ~a10586;
assign a14334 = ~a14332 & a14330;
assign a14336 = ~l1098 & l890;
assign a14338 = a9086 & ~l890;
assign a14340 = ~a14338 & ~a14336;
assign a14342 = ~a14340 & a10622;
assign a14344 = ~a14342 & a14334;
assign a14346 = a14340 & ~a10622;
assign a14348 = ~a14346 & a14344;
assign a14350 = ~l1016 & l890;
assign a14352 = a9078 & ~l890;
assign a14354 = ~a14352 & ~a14350;
assign a14356 = ~a14354 & a10646;
assign a14358 = ~a14356 & a14348;
assign a14360 = a14354 & ~a10646;
assign a14362 = ~a14360 & a14358;
assign a14364 = ~l1758 & l890;
assign a14366 = a5178 & ~l890;
assign a14368 = ~a14366 & ~a14364;
assign a14370 = ~a14368 & a14362;
assign a14372 = ~a14370 & a14270;
assign a14374 = a14372 & a5562;
assign a14376 = a14374 & a5408;
assign a14378 = a14376 & a5404;
assign a14380 = a14378 & a5594;
assign a14382 = a14378 & l992;
assign a14384 = ~a14378 & i452;
assign a14386 = ~a14384 & ~a14382;
assign a14388 = ~a14386 & ~i252;
assign a14390 = i454 & i252;
assign a14392 = ~a14390 & ~a14388;
assign a14394 = ~a14392 & ~l1614;
assign a14396 = a14392 & l1614;
assign a14398 = ~a14396 & ~a14394;
assign a14400 = a14378 & ~a10646;
assign a14402 = ~a14378 & i456;
assign a14404 = ~a14402 & ~a14400;
assign a14406 = ~a14404 & ~i252;
assign a14408 = i458 & i252;
assign a14410 = ~a14408 & ~a14406;
assign a14412 = ~a14410 & a12888;
assign a14414 = a14378 & ~a10622;
assign a14416 = ~a14378 & i460;
assign a14418 = ~a14416 & ~a14414;
assign a14420 = ~a14418 & ~i252;
assign a14422 = i462 & i252;
assign a14424 = ~a14422 & ~a14420;
assign a14426 = ~a14424 & a13072;
assign a14428 = ~a14426 & ~a14412;
assign a14430 = a14424 & ~a13072;
assign a14432 = ~a14430 & ~a14428;
assign a14434 = a14378 & ~a10586;
assign a14436 = ~a14378 & i464;
assign a14438 = ~a14436 & ~a14434;
assign a14440 = ~a14438 & ~i252;
assign a14442 = i466 & i252;
assign a14444 = ~a14442 & ~a14440;
assign a14446 = ~a14444 & a13262;
assign a14448 = ~a14446 & ~a14432;
assign a14450 = a14444 & ~a13262;
assign a14452 = ~a14450 & ~a14448;
assign a14454 = a14378 & ~a10550;
assign a14456 = ~a14378 & i468;
assign a14458 = ~a14456 & ~a14454;
assign a14460 = ~a14458 & ~i252;
assign a14462 = i470 & i252;
assign a14464 = ~a14462 & ~a14460;
assign a14466 = ~a14464 & a13452;
assign a14468 = ~a14466 & ~a14452;
assign a14470 = a14464 & ~a13452;
assign a14472 = ~a14470 & ~a14468;
assign a14474 = a14378 & ~a10514;
assign a14476 = ~a14378 & i472;
assign a14478 = ~a14476 & ~a14474;
assign a14480 = ~a14478 & ~i252;
assign a14482 = i474 & i252;
assign a14484 = ~a14482 & ~a14480;
assign a14486 = ~a14484 & a13642;
assign a14488 = ~a14486 & ~a14472;
assign a14490 = a14484 & ~a13642;
assign a14492 = ~a14490 & ~a14488;
assign a14494 = a14378 & ~a10478;
assign a14496 = ~a14378 & i476;
assign a14498 = ~a14496 & ~a14494;
assign a14500 = ~a14498 & ~i252;
assign a14502 = i478 & i252;
assign a14504 = ~a14502 & ~a14500;
assign a14506 = ~a14504 & a13832;
assign a14508 = ~a14506 & ~a14492;
assign a14510 = a14504 & ~a13832;
assign a14512 = ~a14510 & ~a14508;
assign a14514 = a14378 & l1140;
assign a14516 = ~a14378 & i480;
assign a14518 = ~a14516 & ~a14514;
assign a14520 = ~a14518 & ~i252;
assign a14522 = i482 & i252;
assign a14524 = ~a14522 & ~a14520;
assign a14526 = ~a14524 & ~l1754;
assign a14528 = ~a14526 & ~a14512;
assign a14530 = a14524 & l1754;
assign a14532 = ~a14530 & ~a14528;
assign a14534 = ~a14532 & a14398;
assign a14536 = a14532 & ~a14398;
assign a14538 = ~a14536 & ~a14534;
assign a14540 = ~a14538 & a14380;
assign a14542 = ~l1562 & l890;
assign a14544 = a2764 & ~l890;
assign a14546 = ~a14544 & ~a14542;
assign a14548 = ~l1568 & l890;
assign a14550 = a2736 & ~l890;
assign a14552 = ~a14550 & ~a14548;
assign a14554 = ~l1566 & ~l1558;
assign a14556 = a14554 & a14552;
assign a14558 = a14556 & ~a14546;
assign a14560 = ~a14558 & ~a14540;
assign a14562 = ~a14392 & ~l1330;
assign a14564 = a14392 & l1330;
assign a14566 = ~a14564 & ~a14562;
assign a14568 = a14410 & ~a12974;
assign a14570 = a14424 & ~a13158;
assign a14572 = ~a14570 & ~a14568;
assign a14574 = ~a14424 & a13158;
assign a14576 = ~a14574 & ~a14572;
assign a14578 = a14444 & ~a13348;
assign a14580 = ~a14578 & ~a14576;
assign a14582 = ~a14444 & a13348;
assign a14584 = ~a14582 & ~a14580;
assign a14586 = a14464 & ~a13538;
assign a14588 = ~a14586 & ~a14584;
assign a14590 = ~a14464 & a13538;
assign a14592 = ~a14590 & ~a14588;
assign a14594 = a14484 & ~a13728;
assign a14596 = ~a14594 & ~a14592;
assign a14598 = ~a14484 & a13728;
assign a14600 = ~a14598 & ~a14596;
assign a14602 = a14504 & ~a13906;
assign a14604 = ~a14602 & ~a14600;
assign a14606 = ~a14504 & a13906;
assign a14608 = ~a14606 & ~a14604;
assign a14610 = a14524 & l1470;
assign a14612 = ~a14610 & ~a14608;
assign a14614 = ~a14524 & ~l1470;
assign a14616 = ~a14614 & ~a14612;
assign a14618 = ~a14616 & a14566;
assign a14620 = ~a14410 & a12974;
assign a14622 = ~a14620 & ~a14574;
assign a14624 = ~a14622 & ~a14570;
assign a14626 = ~a14624 & ~a14582;
assign a14628 = ~a14626 & ~a14578;
assign a14630 = ~a14628 & ~a14590;
assign a14632 = ~a14630 & ~a14586;
assign a14634 = ~a14632 & ~a14598;
assign a14636 = ~a14634 & ~a14594;
assign a14638 = ~a14636 & ~a14606;
assign a14640 = ~a14638 & ~a14602;
assign a14642 = ~a14640 & ~a14614;
assign a14644 = ~a14642 & ~a14610;
assign a14646 = ~a14644 & ~a14566;
assign a14648 = ~a14646 & ~a14618;
assign a14650 = ~a14648 & ~a14560;
assign a14652 = a14650 & a12574;
assign a14654 = a14652 & a14380;
assign a14656 = ~a14654 & ~l886;
assign a14658 = a14378 & a5600;
assign a14660 = ~a14392 & ~l1612;
assign a14662 = a14392 & l1612;
assign a14664 = ~a14662 & ~a14660;
assign a14666 = ~a14410 & ~l1632;
assign a14668 = ~a14424 & ~l1652;
assign a14670 = ~a14668 & ~a14666;
assign a14672 = a14424 & l1652;
assign a14674 = ~a14672 & ~a14670;
assign a14676 = ~a14444 & ~l1672;
assign a14678 = ~a14676 & ~a14674;
assign a14680 = a14444 & l1672;
assign a14682 = ~a14680 & ~a14678;
assign a14684 = ~a14464 & ~l1692;
assign a14686 = ~a14684 & ~a14682;
assign a14688 = a14464 & l1692;
assign a14690 = ~a14688 & ~a14686;
assign a14692 = ~a14484 & ~l1712;
assign a14694 = ~a14692 & ~a14690;
assign a14696 = a14484 & l1712;
assign a14698 = ~a14696 & ~a14694;
assign a14700 = ~a14504 & ~l1732;
assign a14702 = ~a14700 & ~a14698;
assign a14704 = a14504 & l1732;
assign a14706 = ~a14704 & ~a14702;
assign a14708 = ~a14524 & ~l1752;
assign a14710 = ~a14708 & ~a14706;
assign a14712 = a14524 & l1752;
assign a14714 = ~a14712 & ~a14710;
assign a14716 = ~a14714 & a14664;
assign a14718 = a14714 & ~a14664;
assign a14720 = ~a14718 & ~a14716;
assign a14722 = ~a14720 & a14658;
assign a14724 = ~a14552 & ~l1558;
assign a14726 = a14724 & a14546;
assign a14728 = a14726 & ~l1566;
assign a14730 = ~a14728 & ~a14722;
assign a14732 = ~a14392 & ~l1328;
assign a14734 = a14392 & l1328;
assign a14736 = ~a14734 & ~a14732;
assign a14738 = a14410 & ~a12962;
assign a14740 = a14424 & ~a13146;
assign a14742 = ~a14740 & ~a14738;
assign a14744 = ~a14424 & a13146;
assign a14746 = ~a14744 & ~a14742;
assign a14748 = a14444 & ~a13336;
assign a14750 = ~a14748 & ~a14746;
assign a14752 = ~a14444 & a13336;
assign a14754 = ~a14752 & ~a14750;
assign a14756 = a14464 & ~a13526;
assign a14758 = ~a14756 & ~a14754;
assign a14760 = ~a14464 & a13526;
assign a14762 = ~a14760 & ~a14758;
assign a14764 = a14484 & ~a13716;
assign a14766 = ~a14764 & ~a14762;
assign a14768 = ~a14484 & a13716;
assign a14770 = ~a14768 & ~a14766;
assign a14772 = a14504 & ~a13894;
assign a14774 = ~a14772 & ~a14770;
assign a14776 = ~a14504 & a13894;
assign a14778 = ~a14776 & ~a14774;
assign a14780 = a14524 & ~a14058;
assign a14782 = ~a14780 & ~a14778;
assign a14784 = ~a14524 & a14058;
assign a14786 = ~a14784 & ~a14782;
assign a14788 = ~a14786 & a14736;
assign a14790 = ~a14410 & a12962;
assign a14792 = ~a14790 & ~a14744;
assign a14794 = ~a14792 & ~a14740;
assign a14796 = ~a14794 & ~a14752;
assign a14798 = ~a14796 & ~a14748;
assign a14800 = ~a14798 & ~a14760;
assign a14802 = ~a14800 & ~a14756;
assign a14804 = ~a14802 & ~a14768;
assign a14806 = ~a14804 & ~a14764;
assign a14808 = ~a14806 & ~a14776;
assign a14810 = ~a14808 & ~a14772;
assign a14812 = ~a14810 & ~a14784;
assign a14814 = ~a14812 & ~a14780;
assign a14816 = ~a14814 & ~a14736;
assign a14818 = ~a14816 & ~a14788;
assign a14820 = ~a14818 & ~a14730;
assign a14822 = a14820 & l1592;
assign a14824 = a14822 & a14658;
assign a14826 = ~a14824 & ~l886;
assign a14828 = a14378 & a5606;
assign a14830 = ~a14392 & ~l1610;
assign a14832 = a14392 & l1610;
assign a14834 = ~a14832 & ~a14830;
assign a14836 = ~a14410 & ~l1630;
assign a14838 = ~a14424 & ~l1650;
assign a14840 = ~a14838 & ~a14836;
assign a14842 = a14424 & l1650;
assign a14844 = ~a14842 & ~a14840;
assign a14846 = ~a14444 & ~l1670;
assign a14848 = ~a14846 & ~a14844;
assign a14850 = a14444 & l1670;
assign a14852 = ~a14850 & ~a14848;
assign a14854 = ~a14464 & ~l1690;
assign a14856 = ~a14854 & ~a14852;
assign a14858 = a14464 & l1690;
assign a14860 = ~a14858 & ~a14856;
assign a14862 = ~a14484 & ~l1710;
assign a14864 = ~a14862 & ~a14860;
assign a14866 = a14484 & l1710;
assign a14868 = ~a14866 & ~a14864;
assign a14870 = ~a14504 & ~l1730;
assign a14872 = ~a14870 & ~a14868;
assign a14874 = a14504 & l1730;
assign a14876 = ~a14874 & ~a14872;
assign a14878 = ~a14524 & ~l1750;
assign a14880 = ~a14878 & ~a14876;
assign a14882 = a14524 & l1750;
assign a14884 = ~a14882 & ~a14880;
assign a14886 = ~a14884 & a14834;
assign a14888 = a14884 & ~a14834;
assign a14890 = ~a14888 & ~a14886;
assign a14892 = ~a14890 & a14828;
assign a14894 = a14724 & ~a14546;
assign a14896 = a14894 & ~l1566;
assign a14898 = ~a14896 & ~a14892;
assign a14900 = ~a14392 & ~l1326;
assign a14902 = a14392 & l1326;
assign a14904 = ~a14902 & ~a14900;
assign a14906 = a14410 & ~a12954;
assign a14908 = a14424 & ~a13138;
assign a14910 = ~a14908 & ~a14906;
assign a14912 = ~a14424 & a13138;
assign a14914 = ~a14912 & ~a14910;
assign a14916 = a14444 & ~a13328;
assign a14918 = ~a14916 & ~a14914;
assign a14920 = ~a14444 & a13328;
assign a14922 = ~a14920 & ~a14918;
assign a14924 = a14464 & ~a13518;
assign a14926 = ~a14924 & ~a14922;
assign a14928 = ~a14464 & a13518;
assign a14930 = ~a14928 & ~a14926;
assign a14932 = a14484 & ~a13708;
assign a14934 = ~a14932 & ~a14930;
assign a14936 = ~a14484 & a13708;
assign a14938 = ~a14936 & ~a14934;
assign a14940 = a14504 & ~a13886;
assign a14942 = ~a14940 & ~a14938;
assign a14944 = ~a14504 & a13886;
assign a14946 = ~a14944 & ~a14942;
assign a14948 = a14524 & ~a14050;
assign a14950 = ~a14948 & ~a14946;
assign a14952 = ~a14524 & a14050;
assign a14954 = ~a14952 & ~a14950;
assign a14956 = ~a14954 & a14904;
assign a14958 = ~a14410 & a12954;
assign a14960 = ~a14958 & ~a14912;
assign a14962 = ~a14960 & ~a14908;
assign a14964 = ~a14962 & ~a14920;
assign a14966 = ~a14964 & ~a14916;
assign a14968 = ~a14966 & ~a14928;
assign a14970 = ~a14968 & ~a14924;
assign a14972 = ~a14970 & ~a14936;
assign a14974 = ~a14972 & ~a14932;
assign a14976 = ~a14974 & ~a14944;
assign a14978 = ~a14976 & ~a14940;
assign a14980 = ~a14978 & ~a14952;
assign a14982 = ~a14980 & ~a14948;
assign a14984 = ~a14982 & ~a14904;
assign a14986 = ~a14984 & ~a14956;
assign a14988 = ~a14986 & ~a14898;
assign a14990 = a14988 & l1590;
assign a14992 = a14990 & a14828;
assign a14994 = ~a14992 & ~l886;
assign a14996 = a14378 & l960;
assign a14998 = ~a14392 & ~l1608;
assign a15000 = a14392 & l1608;
assign a15002 = ~a15000 & ~a14998;
assign a15004 = ~a14410 & ~l1628;
assign a15006 = ~a14424 & ~l1648;
assign a15008 = ~a15006 & ~a15004;
assign a15010 = a14424 & l1648;
assign a15012 = ~a15010 & ~a15008;
assign a15014 = ~a14444 & ~l1668;
assign a15016 = ~a15014 & ~a15012;
assign a15018 = a14444 & l1668;
assign a15020 = ~a15018 & ~a15016;
assign a15022 = ~a14464 & ~l1688;
assign a15024 = ~a15022 & ~a15020;
assign a15026 = a14464 & l1688;
assign a15028 = ~a15026 & ~a15024;
assign a15030 = ~a14484 & ~l1708;
assign a15032 = ~a15030 & ~a15028;
assign a15034 = a14484 & l1708;
assign a15036 = ~a15034 & ~a15032;
assign a15038 = ~a14504 & ~l1728;
assign a15040 = ~a15038 & ~a15036;
assign a15042 = a14504 & l1728;
assign a15044 = ~a15042 & ~a15040;
assign a15046 = ~a14524 & ~l1748;
assign a15048 = ~a15046 & ~a15044;
assign a15050 = a14524 & l1748;
assign a15052 = ~a15050 & ~a15048;
assign a15054 = ~a15052 & a15002;
assign a15056 = a15052 & ~a15002;
assign a15058 = ~a15056 & ~a15054;
assign a15060 = ~a15058 & a14996;
assign a15062 = l1566 & ~l1558;
assign a15064 = a15062 & a14552;
assign a15066 = a15064 & a14546;
assign a15068 = ~a15066 & ~a15060;
assign a15070 = ~a14392 & ~l1324;
assign a15072 = a14392 & l1324;
assign a15074 = ~a15072 & ~a15070;
assign a15076 = a14410 & l1344;
assign a15078 = a14424 & l1364;
assign a15080 = ~a15078 & ~a15076;
assign a15082 = ~a14424 & ~l1364;
assign a15084 = ~a15082 & ~a15080;
assign a15086 = a14444 & l1384;
assign a15088 = ~a15086 & ~a15084;
assign a15090 = ~a14444 & ~l1384;
assign a15092 = ~a15090 & ~a15088;
assign a15094 = a14464 & l1404;
assign a15096 = ~a15094 & ~a15092;
assign a15098 = ~a14464 & ~l1404;
assign a15100 = ~a15098 & ~a15096;
assign a15102 = a14484 & l1424;
assign a15104 = ~a15102 & ~a15100;
assign a15106 = ~a14484 & ~l1424;
assign a15108 = ~a15106 & ~a15104;
assign a15110 = a14504 & l1444;
assign a15112 = ~a15110 & ~a15108;
assign a15114 = ~a14504 & ~l1444;
assign a15116 = ~a15114 & ~a15112;
assign a15118 = a14524 & l1464;
assign a15120 = ~a15118 & ~a15116;
assign a15122 = ~a14524 & ~l1464;
assign a15124 = ~a15122 & ~a15120;
assign a15126 = ~a15124 & a15074;
assign a15128 = ~a14410 & ~l1344;
assign a15130 = ~a15128 & ~a15082;
assign a15132 = ~a15130 & ~a15078;
assign a15134 = ~a15132 & ~a15090;
assign a15136 = ~a15134 & ~a15086;
assign a15138 = ~a15136 & ~a15098;
assign a15140 = ~a15138 & ~a15094;
assign a15142 = ~a15140 & ~a15106;
assign a15144 = ~a15142 & ~a15102;
assign a15146 = ~a15144 & ~a15114;
assign a15148 = ~a15146 & ~a15110;
assign a15150 = ~a15148 & ~a15122;
assign a15152 = ~a15150 & ~a15118;
assign a15154 = ~a15152 & ~a15074;
assign a15156 = ~a15154 & ~a15126;
assign a15158 = ~a15156 & ~a15068;
assign a15160 = a15158 & l1588;
assign a15162 = a15160 & a14996;
assign a15164 = ~a15162 & ~l886;
assign a15166 = a14378 & l962;
assign a15168 = ~a14392 & ~l1606;
assign a15170 = a14392 & l1606;
assign a15172 = ~a15170 & ~a15168;
assign a15174 = ~a14410 & ~l1626;
assign a15176 = ~a14424 & ~l1646;
assign a15178 = ~a15176 & ~a15174;
assign a15180 = a14424 & l1646;
assign a15182 = ~a15180 & ~a15178;
assign a15184 = ~a14444 & ~l1666;
assign a15186 = ~a15184 & ~a15182;
assign a15188 = a14444 & l1666;
assign a15190 = ~a15188 & ~a15186;
assign a15192 = ~a14464 & ~l1686;
assign a15194 = ~a15192 & ~a15190;
assign a15196 = a14464 & l1686;
assign a15198 = ~a15196 & ~a15194;
assign a15200 = ~a14484 & ~l1706;
assign a15202 = ~a15200 & ~a15198;
assign a15204 = a14484 & l1706;
assign a15206 = ~a15204 & ~a15202;
assign a15208 = ~a14504 & ~l1726;
assign a15210 = ~a15208 & ~a15206;
assign a15212 = a14504 & l1726;
assign a15214 = ~a15212 & ~a15210;
assign a15216 = ~a14524 & ~l1746;
assign a15218 = ~a15216 & ~a15214;
assign a15220 = a14524 & l1746;
assign a15222 = ~a15220 & ~a15218;
assign a15224 = ~a15222 & a15172;
assign a15226 = a15222 & ~a15172;
assign a15228 = ~a15226 & ~a15224;
assign a15230 = ~a15228 & a15166;
assign a15232 = a15064 & ~a14546;
assign a15234 = ~a15232 & ~a15230;
assign a15236 = ~a14392 & ~l1322;
assign a15238 = a14392 & l1322;
assign a15240 = ~a15238 & ~a15236;
assign a15242 = a14410 & l1342;
assign a15244 = a14424 & l1362;
assign a15246 = ~a15244 & ~a15242;
assign a15248 = ~a14424 & ~l1362;
assign a15250 = ~a15248 & ~a15246;
assign a15252 = a14444 & l1382;
assign a15254 = ~a15252 & ~a15250;
assign a15256 = ~a14444 & ~l1382;
assign a15258 = ~a15256 & ~a15254;
assign a15260 = a14464 & l1402;
assign a15262 = ~a15260 & ~a15258;
assign a15264 = ~a14464 & ~l1402;
assign a15266 = ~a15264 & ~a15262;
assign a15268 = a14484 & l1422;
assign a15270 = ~a15268 & ~a15266;
assign a15272 = ~a14484 & ~l1422;
assign a15274 = ~a15272 & ~a15270;
assign a15276 = a14504 & l1442;
assign a15278 = ~a15276 & ~a15274;
assign a15280 = ~a14504 & ~l1442;
assign a15282 = ~a15280 & ~a15278;
assign a15284 = a14524 & l1462;
assign a15286 = ~a15284 & ~a15282;
assign a15288 = ~a14524 & ~l1462;
assign a15290 = ~a15288 & ~a15286;
assign a15292 = ~a15290 & a15240;
assign a15294 = ~a14410 & ~l1342;
assign a15296 = ~a15294 & ~a15248;
assign a15298 = ~a15296 & ~a15244;
assign a15300 = ~a15298 & ~a15256;
assign a15302 = ~a15300 & ~a15252;
assign a15304 = ~a15302 & ~a15264;
assign a15306 = ~a15304 & ~a15260;
assign a15308 = ~a15306 & ~a15272;
assign a15310 = ~a15308 & ~a15268;
assign a15312 = ~a15310 & ~a15280;
assign a15314 = ~a15312 & ~a15276;
assign a15316 = ~a15314 & ~a15288;
assign a15318 = ~a15316 & ~a15284;
assign a15320 = ~a15318 & ~a15240;
assign a15322 = ~a15320 & ~a15292;
assign a15324 = ~a15322 & ~a15234;
assign a15326 = a15324 & l1586;
assign a15328 = a15326 & a15166;
assign a15330 = ~a15328 & ~l886;
assign a15332 = a14378 & l964;
assign a15334 = ~a14392 & ~l1604;
assign a15336 = a14392 & l1604;
assign a15338 = ~a15336 & ~a15334;
assign a15340 = ~a14410 & ~l1624;
assign a15342 = ~a14424 & ~l1644;
assign a15344 = ~a15342 & ~a15340;
assign a15346 = a14424 & l1644;
assign a15348 = ~a15346 & ~a15344;
assign a15350 = ~a14444 & ~l1664;
assign a15352 = ~a15350 & ~a15348;
assign a15354 = a14444 & l1664;
assign a15356 = ~a15354 & ~a15352;
assign a15358 = ~a14464 & ~l1684;
assign a15360 = ~a15358 & ~a15356;
assign a15362 = a14464 & l1684;
assign a15364 = ~a15362 & ~a15360;
assign a15366 = ~a14484 & ~l1704;
assign a15368 = ~a15366 & ~a15364;
assign a15370 = a14484 & l1704;
assign a15372 = ~a15370 & ~a15368;
assign a15374 = ~a14504 & ~l1724;
assign a15376 = ~a15374 & ~a15372;
assign a15378 = a14504 & l1724;
assign a15380 = ~a15378 & ~a15376;
assign a15382 = ~a14524 & ~l1744;
assign a15384 = ~a15382 & ~a15380;
assign a15386 = a14524 & l1744;
assign a15388 = ~a15386 & ~a15384;
assign a15390 = ~a15388 & a15338;
assign a15392 = a15388 & ~a15338;
assign a15394 = ~a15392 & ~a15390;
assign a15396 = ~a15394 & a15332;
assign a15398 = a14726 & l1566;
assign a15400 = ~a15398 & ~a15396;
assign a15402 = ~a14392 & ~l1320;
assign a15404 = a14392 & l1320;
assign a15406 = ~a15404 & ~a15402;
assign a15408 = a14410 & l1340;
assign a15410 = a14424 & l1360;
assign a15412 = ~a15410 & ~a15408;
assign a15414 = ~a14424 & ~l1360;
assign a15416 = ~a15414 & ~a15412;
assign a15418 = a14444 & l1380;
assign a15420 = ~a15418 & ~a15416;
assign a15422 = ~a14444 & ~l1380;
assign a15424 = ~a15422 & ~a15420;
assign a15426 = a14464 & l1400;
assign a15428 = ~a15426 & ~a15424;
assign a15430 = ~a14464 & ~l1400;
assign a15432 = ~a15430 & ~a15428;
assign a15434 = a14484 & l1420;
assign a15436 = ~a15434 & ~a15432;
assign a15438 = ~a14484 & ~l1420;
assign a15440 = ~a15438 & ~a15436;
assign a15442 = a14504 & l1440;
assign a15444 = ~a15442 & ~a15440;
assign a15446 = ~a14504 & ~l1440;
assign a15448 = ~a15446 & ~a15444;
assign a15450 = a14524 & l1460;
assign a15452 = ~a15450 & ~a15448;
assign a15454 = ~a14524 & ~l1460;
assign a15456 = ~a15454 & ~a15452;
assign a15458 = ~a15456 & a15406;
assign a15460 = ~a14410 & ~l1340;
assign a15462 = ~a15460 & ~a15414;
assign a15464 = ~a15462 & ~a15410;
assign a15466 = ~a15464 & ~a15422;
assign a15468 = ~a15466 & ~a15418;
assign a15470 = ~a15468 & ~a15430;
assign a15472 = ~a15470 & ~a15426;
assign a15474 = ~a15472 & ~a15438;
assign a15476 = ~a15474 & ~a15434;
assign a15478 = ~a15476 & ~a15446;
assign a15480 = ~a15478 & ~a15442;
assign a15482 = ~a15480 & ~a15454;
assign a15484 = ~a15482 & ~a15450;
assign a15486 = ~a15484 & ~a15406;
assign a15488 = ~a15486 & ~a15458;
assign a15490 = ~a15488 & ~a15400;
assign a15492 = a15490 & l1584;
assign a15494 = a15492 & a15332;
assign a15496 = ~a15494 & ~l886;
assign a15498 = a14378 & l966;
assign a15500 = ~a14392 & ~l1602;
assign a15502 = a14392 & l1602;
assign a15504 = ~a15502 & ~a15500;
assign a15506 = ~a14410 & ~l1622;
assign a15508 = ~a14424 & ~l1642;
assign a15510 = ~a15508 & ~a15506;
assign a15512 = a14424 & l1642;
assign a15514 = ~a15512 & ~a15510;
assign a15516 = ~a14444 & ~l1662;
assign a15518 = ~a15516 & ~a15514;
assign a15520 = a14444 & l1662;
assign a15522 = ~a15520 & ~a15518;
assign a15524 = ~a14464 & ~l1682;
assign a15526 = ~a15524 & ~a15522;
assign a15528 = a14464 & l1682;
assign a15530 = ~a15528 & ~a15526;
assign a15532 = ~a14484 & ~l1702;
assign a15534 = ~a15532 & ~a15530;
assign a15536 = a14484 & l1702;
assign a15538 = ~a15536 & ~a15534;
assign a15540 = ~a14504 & ~l1722;
assign a15542 = ~a15540 & ~a15538;
assign a15544 = a14504 & l1722;
assign a15546 = ~a15544 & ~a15542;
assign a15548 = ~a14524 & ~l1742;
assign a15550 = ~a15548 & ~a15546;
assign a15552 = a14524 & l1742;
assign a15554 = ~a15552 & ~a15550;
assign a15556 = ~a15554 & a15504;
assign a15558 = a15554 & ~a15504;
assign a15560 = ~a15558 & ~a15556;
assign a15562 = ~a15560 & a15498;
assign a15564 = a14894 & l1566;
assign a15566 = ~a15564 & ~a15562;
assign a15568 = ~a14392 & ~l1318;
assign a15570 = a14392 & l1318;
assign a15572 = ~a15570 & ~a15568;
assign a15574 = a14410 & l1338;
assign a15576 = a14424 & l1358;
assign a15578 = ~a15576 & ~a15574;
assign a15580 = ~a14424 & ~l1358;
assign a15582 = ~a15580 & ~a15578;
assign a15584 = a14444 & l1378;
assign a15586 = ~a15584 & ~a15582;
assign a15588 = ~a14444 & ~l1378;
assign a15590 = ~a15588 & ~a15586;
assign a15592 = a14464 & l1398;
assign a15594 = ~a15592 & ~a15590;
assign a15596 = ~a14464 & ~l1398;
assign a15598 = ~a15596 & ~a15594;
assign a15600 = a14484 & l1418;
assign a15602 = ~a15600 & ~a15598;
assign a15604 = ~a14484 & ~l1418;
assign a15606 = ~a15604 & ~a15602;
assign a15608 = a14504 & l1438;
assign a15610 = ~a15608 & ~a15606;
assign a15612 = ~a14504 & ~l1438;
assign a15614 = ~a15612 & ~a15610;
assign a15616 = a14524 & l1458;
assign a15618 = ~a15616 & ~a15614;
assign a15620 = ~a14524 & ~l1458;
assign a15622 = ~a15620 & ~a15618;
assign a15624 = ~a15622 & a15572;
assign a15626 = ~a14410 & ~l1338;
assign a15628 = ~a15626 & ~a15580;
assign a15630 = ~a15628 & ~a15576;
assign a15632 = ~a15630 & ~a15588;
assign a15634 = ~a15632 & ~a15584;
assign a15636 = ~a15634 & ~a15596;
assign a15638 = ~a15636 & ~a15592;
assign a15640 = ~a15638 & ~a15604;
assign a15642 = ~a15640 & ~a15600;
assign a15644 = ~a15642 & ~a15612;
assign a15646 = ~a15644 & ~a15608;
assign a15648 = ~a15646 & ~a15620;
assign a15650 = ~a15648 & ~a15616;
assign a15652 = ~a15650 & ~a15572;
assign a15654 = ~a15652 & ~a15624;
assign a15656 = ~a15654 & ~a15566;
assign a15658 = a15656 & l1542;
assign a15660 = a15658 & a15498;
assign a15662 = ~a15660 & ~l886;
assign a15664 = a14378 & l970;
assign a15666 = ~a14392 & ~l1600;
assign a15668 = a14392 & l1600;
assign a15670 = ~a15668 & ~a15666;
assign a15672 = ~a14410 & ~l1620;
assign a15674 = ~a14424 & ~l1640;
assign a15676 = ~a15674 & ~a15672;
assign a15678 = a14424 & l1640;
assign a15680 = ~a15678 & ~a15676;
assign a15682 = ~a14444 & ~l1660;
assign a15684 = ~a15682 & ~a15680;
assign a15686 = a14444 & l1660;
assign a15688 = ~a15686 & ~a15684;
assign a15690 = ~a14464 & ~l1680;
assign a15692 = ~a15690 & ~a15688;
assign a15694 = a14464 & l1680;
assign a15696 = ~a15694 & ~a15692;
assign a15698 = ~a14484 & ~l1700;
assign a15700 = ~a15698 & ~a15696;
assign a15702 = a14484 & l1700;
assign a15704 = ~a15702 & ~a15700;
assign a15706 = ~a14504 & ~l1720;
assign a15708 = ~a15706 & ~a15704;
assign a15710 = a14504 & l1720;
assign a15712 = ~a15710 & ~a15708;
assign a15714 = ~a14524 & ~l1740;
assign a15716 = ~a15714 & ~a15712;
assign a15718 = a14524 & l1740;
assign a15720 = ~a15718 & ~a15716;
assign a15722 = ~a15720 & a15670;
assign a15724 = a15720 & ~a15670;
assign a15726 = ~a15724 & ~a15722;
assign a15728 = ~a15726 & a15664;
assign a15730 = ~l1566 & l1558;
assign a15732 = a15730 & a14552;
assign a15734 = a15732 & a14546;
assign a15736 = ~a15734 & ~a15728;
assign a15738 = ~a14392 & ~l1316;
assign a15740 = a14392 & l1316;
assign a15742 = ~a15740 & ~a15738;
assign a15744 = a14410 & l1336;
assign a15746 = a14424 & l1356;
assign a15748 = ~a15746 & ~a15744;
assign a15750 = ~a14424 & ~l1356;
assign a15752 = ~a15750 & ~a15748;
assign a15754 = a14444 & l1376;
assign a15756 = ~a15754 & ~a15752;
assign a15758 = ~a14444 & ~l1376;
assign a15760 = ~a15758 & ~a15756;
assign a15762 = a14464 & l1396;
assign a15764 = ~a15762 & ~a15760;
assign a15766 = ~a14464 & ~l1396;
assign a15768 = ~a15766 & ~a15764;
assign a15770 = a14484 & l1416;
assign a15772 = ~a15770 & ~a15768;
assign a15774 = ~a14484 & ~l1416;
assign a15776 = ~a15774 & ~a15772;
assign a15778 = a14504 & l1436;
assign a15780 = ~a15778 & ~a15776;
assign a15782 = ~a14504 & ~l1436;
assign a15784 = ~a15782 & ~a15780;
assign a15786 = a14524 & l1456;
assign a15788 = ~a15786 & ~a15784;
assign a15790 = ~a14524 & ~l1456;
assign a15792 = ~a15790 & ~a15788;
assign a15794 = ~a15792 & a15742;
assign a15796 = ~a14410 & ~l1336;
assign a15798 = ~a15796 & ~a15750;
assign a15800 = ~a15798 & ~a15746;
assign a15802 = ~a15800 & ~a15758;
assign a15804 = ~a15802 & ~a15754;
assign a15806 = ~a15804 & ~a15766;
assign a15808 = ~a15806 & ~a15762;
assign a15810 = ~a15808 & ~a15774;
assign a15812 = ~a15810 & ~a15770;
assign a15814 = ~a15812 & ~a15782;
assign a15816 = ~a15814 & ~a15778;
assign a15818 = ~a15816 & ~a15790;
assign a15820 = ~a15818 & ~a15786;
assign a15822 = ~a15820 & ~a15742;
assign a15824 = ~a15822 & ~a15794;
assign a15826 = ~a15824 & ~a15736;
assign a15828 = a15826 & l1514;
assign a15830 = a15828 & a15664;
assign a15832 = ~a15830 & ~l886;
assign a15834 = a14378 & l1510;
assign a15836 = ~a14392 & ~l1598;
assign a15838 = a14392 & l1598;
assign a15840 = ~a15838 & ~a15836;
assign a15842 = ~a14410 & ~l1618;
assign a15844 = ~a14424 & ~l1638;
assign a15846 = ~a15844 & ~a15842;
assign a15848 = a14424 & l1638;
assign a15850 = ~a15848 & ~a15846;
assign a15852 = ~a14444 & ~l1658;
assign a15854 = ~a15852 & ~a15850;
assign a15856 = a14444 & l1658;
assign a15858 = ~a15856 & ~a15854;
assign a15860 = ~a14464 & ~l1678;
assign a15862 = ~a15860 & ~a15858;
assign a15864 = a14464 & l1678;
assign a15866 = ~a15864 & ~a15862;
assign a15868 = ~a14484 & ~l1698;
assign a15870 = ~a15868 & ~a15866;
assign a15872 = a14484 & l1698;
assign a15874 = ~a15872 & ~a15870;
assign a15876 = ~a14504 & ~l1718;
assign a15878 = ~a15876 & ~a15874;
assign a15880 = a14504 & l1718;
assign a15882 = ~a15880 & ~a15878;
assign a15884 = ~a14524 & ~l1738;
assign a15886 = ~a15884 & ~a15882;
assign a15888 = a14524 & l1738;
assign a15890 = ~a15888 & ~a15886;
assign a15892 = ~a15890 & a15840;
assign a15894 = a15890 & ~a15840;
assign a15896 = ~a15894 & ~a15892;
assign a15898 = ~a15896 & l968;
assign a15900 = a15898 & a14378;
assign a15902 = a15732 & ~a14546;
assign a15904 = ~a15902 & ~a15900;
assign a15906 = ~a14392 & ~l1314;
assign a15908 = a14392 & l1314;
assign a15910 = ~a15908 & ~a15906;
assign a15912 = a14410 & l1334;
assign a15914 = a14424 & l1354;
assign a15916 = ~a15914 & ~a15912;
assign a15918 = ~a14424 & ~l1354;
assign a15920 = ~a15918 & ~a15916;
assign a15922 = a14444 & l1374;
assign a15924 = ~a15922 & ~a15920;
assign a15926 = ~a14444 & ~l1374;
assign a15928 = ~a15926 & ~a15924;
assign a15930 = a14464 & l1394;
assign a15932 = ~a15930 & ~a15928;
assign a15934 = ~a14464 & ~l1394;
assign a15936 = ~a15934 & ~a15932;
assign a15938 = a14484 & l1414;
assign a15940 = ~a15938 & ~a15936;
assign a15942 = ~a14484 & ~l1414;
assign a15944 = ~a15942 & ~a15940;
assign a15946 = a14504 & l1434;
assign a15948 = ~a15946 & ~a15944;
assign a15950 = ~a14504 & ~l1434;
assign a15952 = ~a15950 & ~a15948;
assign a15954 = a14524 & l1454;
assign a15956 = ~a15954 & ~a15952;
assign a15958 = ~a14524 & ~l1454;
assign a15960 = ~a15958 & ~a15956;
assign a15962 = ~a15960 & a15910;
assign a15964 = ~a14410 & ~l1334;
assign a15966 = ~a15964 & ~a15918;
assign a15968 = ~a15966 & ~a15914;
assign a15970 = ~a15968 & ~a15926;
assign a15972 = ~a15970 & ~a15922;
assign a15974 = ~a15972 & ~a15934;
assign a15976 = ~a15974 & ~a15930;
assign a15978 = ~a15976 & ~a15942;
assign a15980 = ~a15978 & ~a15938;
assign a15982 = ~a15980 & ~a15950;
assign a15984 = ~a15982 & ~a15946;
assign a15986 = ~a15984 & ~a15958;
assign a15988 = ~a15986 & ~a15954;
assign a15990 = ~a15988 & ~a15910;
assign a15992 = ~a15990 & ~a15962;
assign a15994 = ~a15992 & ~a15904;
assign a15996 = a15994 & l968;
assign a15998 = a15996 & a15834;
assign a16000 = ~a15998 & ~l886;
assign a16002 = a14378 & a5568;
assign a16004 = ~a14392 & ~l1616;
assign a16006 = a14392 & l1616;
assign a16008 = ~a16006 & ~a16004;
assign a16010 = ~a14410 & a12902;
assign a16012 = ~a14424 & a13086;
assign a16014 = ~a16012 & ~a16010;
assign a16016 = a14424 & ~a13086;
assign a16018 = ~a16016 & ~a16014;
assign a16020 = ~a14444 & a13276;
assign a16022 = ~a16020 & ~a16018;
assign a16024 = a14444 & ~a13276;
assign a16026 = ~a16024 & ~a16022;
assign a16028 = ~a14464 & a13466;
assign a16030 = ~a16028 & ~a16026;
assign a16032 = a14464 & ~a13466;
assign a16034 = ~a16032 & ~a16030;
assign a16036 = ~a14484 & a13656;
assign a16038 = ~a16036 & ~a16034;
assign a16040 = a14484 & ~a13656;
assign a16042 = ~a16040 & ~a16038;
assign a16044 = ~a14504 & ~l1736;
assign a16046 = ~a16044 & ~a16042;
assign a16048 = a14504 & l1736;
assign a16050 = ~a16048 & ~a16046;
assign a16052 = ~a14524 & ~l1756;
assign a16054 = ~a16052 & ~a16050;
assign a16056 = a14524 & l1756;
assign a16058 = ~a16056 & ~a16054;
assign a16060 = ~a16058 & a16008;
assign a16062 = a16058 & ~a16008;
assign a16064 = ~a16062 & ~a16060;
assign a16066 = ~a16064 & a16002;
assign a16068 = a14556 & a14546;
assign a16070 = ~a16068 & ~a16066;
assign a16072 = ~a14392 & ~l1332;
assign a16074 = a14392 & l1332;
assign a16076 = ~a16074 & ~a16072;
assign a16078 = a14410 & l1352;
assign a16080 = a14424 & l1372;
assign a16082 = ~a16080 & ~a16078;
assign a16084 = ~a14424 & ~l1372;
assign a16086 = ~a16084 & ~a16082;
assign a16088 = a14444 & l1392;
assign a16090 = ~a16088 & ~a16086;
assign a16092 = ~a14444 & ~l1392;
assign a16094 = ~a16092 & ~a16090;
assign a16096 = a14464 & l1412;
assign a16098 = ~a16096 & ~a16094;
assign a16100 = ~a14464 & ~l1412;
assign a16102 = ~a16100 & ~a16098;
assign a16104 = a14484 & l1432;
assign a16106 = ~a16104 & ~a16102;
assign a16108 = ~a14484 & ~l1432;
assign a16110 = ~a16108 & ~a16106;
assign a16112 = a14504 & l1452;
assign a16114 = ~a16112 & ~a16110;
assign a16116 = ~a14504 & ~l1452;
assign a16118 = ~a16116 & ~a16114;
assign a16120 = a14524 & l1472;
assign a16122 = ~a16120 & ~a16118;
assign a16124 = ~a14524 & ~l1472;
assign a16126 = ~a16124 & ~a16122;
assign a16128 = ~a16126 & a16076;
assign a16130 = ~a14410 & ~l1352;
assign a16132 = ~a16130 & ~a16084;
assign a16134 = ~a16132 & ~a16080;
assign a16136 = ~a16134 & ~a16092;
assign a16138 = ~a16136 & ~a16088;
assign a16140 = ~a16138 & ~a16100;
assign a16142 = ~a16140 & ~a16096;
assign a16144 = ~a16142 & ~a16108;
assign a16146 = ~a16144 & ~a16104;
assign a16148 = ~a16146 & ~a16116;
assign a16150 = ~a16148 & ~a16112;
assign a16152 = ~a16150 & ~a16124;
assign a16154 = ~a16152 & ~a16120;
assign a16156 = ~a16154 & ~a16076;
assign a16158 = ~a16156 & ~a16128;
assign a16160 = ~a16158 & ~a16070;
assign a16162 = a16160 & a12582;
assign a16164 = a16162 & a16002;
assign a16166 = ~a16164 & ~l886;
assign a16168 = a16166 & a16000;
assign a16170 = a16168 & a15832;
assign a16172 = a16170 & a15662;
assign a16174 = a16172 & a15496;
assign a16176 = a16174 & a15330;
assign a16178 = a16176 & a15164;
assign a16180 = a16178 & a14994;
assign a16182 = a16180 & a14826;
assign a16184 = a16182 & a14656;
assign a16188 = ~a9058 & ~l1250;
assign a16190 = a16188 & a9046;
assign a16192 = a16190 & a5394;
assign a16194 = a16192 & i484;
assign a16198 = ~a16196 & a5394;
assign a16200 = ~l984 & l890;
assign a16202 = a5178 & i248;
assign a16204 = a16202 & ~a5370;
assign a16206 = a16204 & ~l890;
assign a16208 = ~a16206 & ~a16200;
assign a16210 = ~l988 & l890;
assign a16212 = a16204 & ~l890;
assign a16214 = ~a16212 & ~a16210;
assign a16216 = a16214 & ~l986;
assign a16218 = a16216 & a16208;
assign a16220 = a16218 & ~l990;
assign a16222 = a16220 & ~l910;
assign a16224 = ~l982 & ~l980;
assign a16226 = a16224 & ~a5352;
assign a16228 = ~l886 & i244;
assign a16230 = ~l1012 & l890;
assign a16232 = a16204 & a3976;
assign a16234 = a16232 & ~l890;
assign a16236 = ~a16234 & ~a16230;
assign a16238 = ~a16236 & ~a16222;
assign a16240 = a16196 & ~a10646;
assign a16242 = ~a14354 & a9060;
assign a16244 = ~a9060 & ~a7226;
assign a16246 = ~a16244 & ~a16242;
assign a16248 = ~a16246 & ~a16196;
assign a16252 = ~a16196 & a16192;
assign a16254 = a16252 & ~l1764;
assign a16256 = ~a16254 & ~a16250;
assign a16258 = a16254 & ~a10646;
assign a16260 = ~a16258 & ~a16256;
assign a16262 = ~a16260 & a16222;
assign a16264 = ~a16262 & ~a16238;
assign a16266 = ~a16222 & l996;
assign a16268 = a16196 & l992;
assign a16270 = a9060 & l994;
assign a16272 = ~a9060 & l1082;
assign a16274 = ~a16272 & ~a16270;
assign a16276 = ~a16274 & ~a16196;
assign a16278 = ~a16276 & ~a16268;
assign a16280 = ~a16278 & ~a16254;
assign a16282 = a16254 & l992;
assign a16284 = ~a16282 & ~a16280;
assign a16286 = ~a16284 & a16222;
assign a16288 = ~a16286 & ~a16266;
assign a16290 = ~a12366 & ~a12312;
assign a16292 = a16290 & ~a12250;
assign a16294 = ~a16292 & ~a12190;
assign a16296 = a16292 & a12190;
assign a16298 = ~a16296 & ~a16294;
assign a16300 = ~a16290 & ~a12250;
assign a16302 = a16290 & a12250;
assign a16304 = ~a16302 & ~a16300;
assign a16306 = ~a12366 & a12312;
assign a16308 = a12366 & ~a12312;
assign a16310 = ~a16308 & ~a16306;
assign a16312 = a12366 & l1318;
assign a16314 = ~a12366 & l1320;
assign a16316 = ~a16314 & ~a16312;
assign a16318 = ~a16316 & ~a16310;
assign a16320 = a12366 & l1322;
assign a16322 = ~a12366 & l1324;
assign a16324 = ~a16322 & ~a16320;
assign a16326 = ~a16324 & a16310;
assign a16328 = ~a16326 & ~a16318;
assign a16330 = ~a16328 & ~a16304;
assign a16332 = a12366 & l1326;
assign a16334 = ~a12366 & l1328;
assign a16336 = ~a16334 & ~a16332;
assign a16338 = ~a16336 & ~a16310;
assign a16340 = a12366 & l1330;
assign a16342 = ~a12366 & l1332;
assign a16344 = ~a16342 & ~a16340;
assign a16346 = ~a16344 & a16310;
assign a16348 = ~a16346 & ~a16338;
assign a16350 = ~a16348 & a16304;
assign a16352 = ~a16350 & ~a16330;
assign a16354 = ~a16352 & a16298;
assign a16356 = a12250 & ~a12190;
assign a16358 = a16356 & a16306;
assign a16360 = a16358 & l1332;
assign a16362 = ~a16360 & ~a16354;
assign a16364 = a16304 & ~a16298;
assign a16366 = a16364 & a16310;
assign a16368 = a12366 & l1314;
assign a16370 = ~a12366 & l1316;
assign a16372 = ~a16370 & ~a16368;
assign a16374 = ~a16372 & a16366;
assign a16376 = ~a16374 & a16362;
assign a16378 = ~l948 & ~l924;
assign a16380 = a16378 & ~l1512;
assign a16382 = a12366 & l968;
assign a16384 = ~a12366 & l970;
assign a16386 = ~a16384 & ~a16382;
assign a16388 = ~a16386 & ~a16298;
assign a16390 = a12366 & l966;
assign a16392 = ~a12366 & l964;
assign a16394 = ~a16392 & ~a16390;
assign a16396 = ~a16394 & ~a16310;
assign a16398 = a12366 & l962;
assign a16400 = ~a12366 & l960;
assign a16402 = ~a16400 & ~a16398;
assign a16404 = ~a16402 & a16310;
assign a16406 = ~a16404 & ~a16396;
assign a16408 = ~a16406 & ~a16304;
assign a16410 = a12366 & a5606;
assign a16412 = ~a12366 & a5600;
assign a16414 = ~a16412 & ~a16410;
assign a16416 = ~a16414 & ~a16310;
assign a16418 = a12366 & a5594;
assign a16420 = ~a12366 & a5568;
assign a16422 = ~a16420 & ~a16418;
assign a16424 = ~a16422 & a16310;
assign a16426 = ~a16424 & ~a16416;
assign a16428 = ~a16426 & a16304;
assign a16430 = ~a16428 & ~a16408;
assign a16432 = ~a16430 & a16298;
assign a16434 = ~a16432 & ~a16388;
assign a16436 = ~a16434 & ~a16358;
assign a16438 = a16358 & a5568;
assign a16442 = ~a16440 & ~a12374;
assign a16444 = a16442 & a16380;
assign a16446 = a16444 & ~a16376;
assign a16448 = ~a16444 & ~a12820;
assign a16450 = ~a16448 & ~a16446;
assign a16452 = ~a16450 & a16288;
assign a16454 = a16450 & ~a16288;
assign a16456 = ~a16454 & ~a16452;
assign a16458 = a12366 & l1338;
assign a16460 = ~a12366 & l1340;
assign a16462 = ~a16460 & ~a16458;
assign a16464 = ~a16462 & ~a16310;
assign a16466 = a12366 & l1342;
assign a16468 = ~a12366 & l1344;
assign a16470 = ~a16468 & ~a16466;
assign a16472 = ~a16470 & a16310;
assign a16474 = ~a16472 & ~a16464;
assign a16476 = ~a16474 & ~a16304;
assign a16478 = ~a12954 & a12366;
assign a16480 = ~a12962 & ~a12366;
assign a16482 = ~a16480 & ~a16478;
assign a16484 = ~a16482 & ~a16310;
assign a16486 = ~a12974 & a12366;
assign a16488 = ~a12366 & l1352;
assign a16490 = ~a16488 & ~a16486;
assign a16492 = ~a16490 & a16310;
assign a16494 = ~a16492 & ~a16484;
assign a16496 = ~a16494 & a16304;
assign a16498 = ~a16496 & ~a16476;
assign a16500 = ~a16498 & a16298;
assign a16502 = a16358 & l1352;
assign a16504 = ~a16502 & ~a16500;
assign a16506 = a12366 & l1334;
assign a16508 = ~a12366 & l1336;
assign a16510 = ~a16508 & ~a16506;
assign a16512 = ~a16510 & a16366;
assign a16516 = ~a16514 & a16444;
assign a16518 = ~a16444 & ~a13008;
assign a16520 = ~a16518 & ~a16516;
assign a16522 = a16520 & ~a16264;
assign a16524 = a12366 & l1358;
assign a16526 = ~a12366 & l1360;
assign a16528 = ~a16526 & ~a16524;
assign a16530 = ~a16528 & ~a16310;
assign a16532 = a12366 & l1362;
assign a16534 = ~a12366 & l1364;
assign a16536 = ~a16534 & ~a16532;
assign a16538 = ~a16536 & a16310;
assign a16540 = ~a16538 & ~a16530;
assign a16542 = ~a16540 & ~a16304;
assign a16544 = ~a13138 & a12366;
assign a16546 = ~a13146 & ~a12366;
assign a16548 = ~a16546 & ~a16544;
assign a16550 = ~a16548 & ~a16310;
assign a16552 = ~a13158 & a12366;
assign a16554 = ~a12366 & l1372;
assign a16556 = ~a16554 & ~a16552;
assign a16558 = ~a16556 & a16310;
assign a16560 = ~a16558 & ~a16550;
assign a16562 = ~a16560 & a16304;
assign a16564 = ~a16562 & ~a16542;
assign a16566 = ~a16564 & a16298;
assign a16568 = a16358 & l1372;
assign a16570 = ~a16568 & ~a16566;
assign a16572 = a12366 & l1354;
assign a16574 = ~a12366 & l1356;
assign a16576 = ~a16574 & ~a16572;
assign a16578 = ~a16576 & a16366;
assign a16582 = ~a16580 & a16444;
assign a16584 = ~a16444 & ~a13192;
assign a16586 = ~a16584 & ~a16582;
assign a16588 = ~l1104 & l890;
assign a16590 = a16204 & a4980;
assign a16592 = a16590 & ~l890;
assign a16594 = ~a16592 & ~a16588;
assign a16596 = ~a16594 & ~a16222;
assign a16598 = a16196 & ~a10622;
assign a16600 = ~a14340 & a9060;
assign a16602 = ~a9060 & ~a6426;
assign a16604 = ~a16602 & ~a16600;
assign a16606 = ~a16604 & ~a16196;
assign a16610 = ~a16608 & ~a16254;
assign a16612 = a16254 & ~a10622;
assign a16614 = ~a16612 & ~a16610;
assign a16616 = ~a16614 & a16222;
assign a16618 = ~a16616 & ~a16596;
assign a16620 = ~a16618 & a16586;
assign a16622 = ~a16620 & ~a16522;
assign a16624 = a16618 & ~a16586;
assign a16626 = ~a16624 & ~a16622;
assign a16628 = a12366 & l1378;
assign a16630 = ~a12366 & l1380;
assign a16632 = ~a16630 & ~a16628;
assign a16634 = ~a16632 & ~a16310;
assign a16636 = a12366 & l1382;
assign a16638 = ~a12366 & l1384;
assign a16640 = ~a16638 & ~a16636;
assign a16642 = ~a16640 & a16310;
assign a16644 = ~a16642 & ~a16634;
assign a16646 = ~a16644 & ~a16304;
assign a16648 = ~a13328 & a12366;
assign a16650 = ~a13336 & ~a12366;
assign a16652 = ~a16650 & ~a16648;
assign a16654 = ~a16652 & ~a16310;
assign a16656 = ~a13348 & a12366;
assign a16658 = ~a12366 & l1392;
assign a16660 = ~a16658 & ~a16656;
assign a16662 = ~a16660 & a16310;
assign a16664 = ~a16662 & ~a16654;
assign a16666 = ~a16664 & a16304;
assign a16668 = ~a16666 & ~a16646;
assign a16670 = ~a16668 & a16298;
assign a16672 = a16358 & l1392;
assign a16674 = ~a16672 & ~a16670;
assign a16676 = a12366 & l1374;
assign a16678 = ~a12366 & l1376;
assign a16680 = ~a16678 & ~a16676;
assign a16682 = ~a16680 & a16366;
assign a16686 = ~a16684 & a16444;
assign a16688 = ~a16444 & ~a13382;
assign a16690 = ~a16688 & ~a16686;
assign a16692 = ~l1112 & l890;
assign a16694 = a16204 & a5028;
assign a16696 = a16694 & ~l890;
assign a16698 = ~a16696 & ~a16692;
assign a16700 = ~a16698 & ~a16222;
assign a16702 = a16196 & ~a10586;
assign a16704 = ~a14326 & a9060;
assign a16706 = ~a9060 & ~a6434;
assign a16708 = ~a16706 & ~a16704;
assign a16710 = ~a16708 & ~a16196;
assign a16714 = ~a16712 & ~a16254;
assign a16716 = a16254 & ~a10586;
assign a16718 = ~a16716 & ~a16714;
assign a16720 = ~a16718 & a16222;
assign a16722 = ~a16720 & ~a16700;
assign a16724 = ~a16722 & a16690;
assign a16726 = ~a16724 & ~a16626;
assign a16728 = a16722 & ~a16690;
assign a16730 = ~a16728 & ~a16726;
assign a16732 = a12366 & l1398;
assign a16734 = ~a12366 & l1400;
assign a16736 = ~a16734 & ~a16732;
assign a16738 = ~a16736 & ~a16310;
assign a16740 = a12366 & l1402;
assign a16742 = ~a12366 & l1404;
assign a16744 = ~a16742 & ~a16740;
assign a16746 = ~a16744 & a16310;
assign a16748 = ~a16746 & ~a16738;
assign a16750 = ~a16748 & ~a16304;
assign a16752 = ~a13518 & a12366;
assign a16754 = ~a13526 & ~a12366;
assign a16756 = ~a16754 & ~a16752;
assign a16758 = ~a16756 & ~a16310;
assign a16760 = ~a13538 & a12366;
assign a16762 = ~a12366 & l1412;
assign a16764 = ~a16762 & ~a16760;
assign a16766 = ~a16764 & a16310;
assign a16768 = ~a16766 & ~a16758;
assign a16770 = ~a16768 & a16304;
assign a16772 = ~a16770 & ~a16750;
assign a16774 = ~a16772 & a16298;
assign a16776 = a16358 & l1412;
assign a16778 = ~a16776 & ~a16774;
assign a16780 = a12366 & l1394;
assign a16782 = ~a12366 & l1396;
assign a16784 = ~a16782 & ~a16780;
assign a16786 = ~a16784 & a16366;
assign a16790 = ~a16788 & a16444;
assign a16792 = ~a16444 & ~a13572;
assign a16794 = ~a16792 & ~a16790;
assign a16796 = ~l1120 & l890;
assign a16798 = a16204 & a5076;
assign a16800 = a16798 & ~l890;
assign a16802 = ~a16800 & ~a16796;
assign a16804 = ~a16802 & ~a16222;
assign a16806 = a16196 & ~a10550;
assign a16808 = ~a14312 & a9060;
assign a16810 = ~a9060 & ~a6442;
assign a16812 = ~a16810 & ~a16808;
assign a16814 = ~a16812 & ~a16196;
assign a16818 = ~a16816 & ~a16254;
assign a16820 = a16254 & ~a10550;
assign a16822 = ~a16820 & ~a16818;
assign a16824 = ~a16822 & a16222;
assign a16826 = ~a16824 & ~a16804;
assign a16828 = ~a16826 & a16794;
assign a16830 = ~a16828 & ~a16730;
assign a16832 = a16826 & ~a16794;
assign a16834 = ~a16832 & ~a16830;
assign a16836 = a12366 & l1418;
assign a16838 = ~a12366 & l1420;
assign a16840 = ~a16838 & ~a16836;
assign a16842 = ~a16840 & ~a16310;
assign a16844 = a12366 & l1422;
assign a16846 = ~a12366 & l1424;
assign a16848 = ~a16846 & ~a16844;
assign a16850 = ~a16848 & a16310;
assign a16852 = ~a16850 & ~a16842;
assign a16854 = ~a16852 & ~a16304;
assign a16856 = ~a13708 & a12366;
assign a16858 = ~a13716 & ~a12366;
assign a16860 = ~a16858 & ~a16856;
assign a16862 = ~a16860 & ~a16310;
assign a16864 = ~a13728 & a12366;
assign a16866 = ~a12366 & l1432;
assign a16868 = ~a16866 & ~a16864;
assign a16870 = ~a16868 & a16310;
assign a16872 = ~a16870 & ~a16862;
assign a16874 = ~a16872 & a16304;
assign a16876 = ~a16874 & ~a16854;
assign a16878 = ~a16876 & a16298;
assign a16880 = a16358 & l1432;
assign a16882 = ~a16880 & ~a16878;
assign a16884 = a12366 & l1414;
assign a16886 = ~a12366 & l1416;
assign a16888 = ~a16886 & ~a16884;
assign a16890 = ~a16888 & a16366;
assign a16894 = ~a16892 & a16444;
assign a16896 = ~a16444 & ~a13762;
assign a16898 = ~a16896 & ~a16894;
assign a16900 = ~l1128 & l890;
assign a16902 = a16204 & a5124;
assign a16904 = a16902 & ~l890;
assign a16906 = ~a16904 & ~a16900;
assign a16908 = ~a16906 & ~a16222;
assign a16910 = a16196 & ~a10514;
assign a16912 = ~a14298 & a9060;
assign a16914 = ~a9060 & ~a6450;
assign a16916 = ~a16914 & ~a16912;
assign a16918 = ~a16916 & ~a16196;
assign a16922 = ~a16920 & ~a16254;
assign a16924 = a16254 & ~a10514;
assign a16926 = ~a16924 & ~a16922;
assign a16928 = ~a16926 & a16222;
assign a16930 = ~a16928 & ~a16908;
assign a16932 = ~a16930 & a16898;
assign a16934 = ~a16932 & ~a16834;
assign a16936 = a16930 & ~a16898;
assign a16938 = ~a16936 & ~a16934;
assign a16940 = a12366 & l1438;
assign a16942 = ~a12366 & l1440;
assign a16944 = ~a16942 & ~a16940;
assign a16946 = ~a16944 & ~a16310;
assign a16948 = a12366 & l1442;
assign a16950 = ~a12366 & l1444;
assign a16952 = ~a16950 & ~a16948;
assign a16954 = ~a16952 & a16310;
assign a16956 = ~a16954 & ~a16946;
assign a16958 = ~a16956 & ~a16304;
assign a16960 = ~a13886 & a12366;
assign a16962 = ~a13894 & ~a12366;
assign a16964 = ~a16962 & ~a16960;
assign a16966 = ~a16964 & ~a16310;
assign a16968 = ~a13906 & a12366;
assign a16970 = ~a12366 & l1452;
assign a16972 = ~a16970 & ~a16968;
assign a16974 = ~a16972 & a16310;
assign a16976 = ~a16974 & ~a16966;
assign a16978 = ~a16976 & a16304;
assign a16980 = ~a16978 & ~a16958;
assign a16982 = ~a16980 & a16298;
assign a16984 = a16358 & l1452;
assign a16986 = ~a16984 & ~a16982;
assign a16988 = a12366 & l1434;
assign a16990 = ~a12366 & l1436;
assign a16992 = ~a16990 & ~a16988;
assign a16994 = ~a16992 & a16366;
assign a16998 = ~a16996 & a16444;
assign a17000 = ~a16444 & ~a13940;
assign a17002 = ~a17000 & ~a16998;
assign a17004 = ~a16222 & l1136;
assign a17006 = a16196 & ~a10478;
assign a17008 = a9060 & l1134;
assign a17010 = ~a9060 & l1130;
assign a17012 = ~a17010 & ~a17008;
assign a17014 = ~a17012 & ~a16196;
assign a17016 = ~a17014 & ~a17006;
assign a17018 = ~a17016 & ~a16254;
assign a17020 = a16254 & ~a10478;
assign a17022 = ~a17020 & ~a17018;
assign a17024 = ~a17022 & a16222;
assign a17026 = ~a17024 & ~a17004;
assign a17028 = ~a17026 & a17002;
assign a17030 = ~a17028 & ~a16938;
assign a17032 = a17026 & ~a17002;
assign a17034 = ~a17032 & ~a17030;
assign a17036 = a12366 & l1458;
assign a17038 = ~a12366 & l1460;
assign a17040 = ~a17038 & ~a17036;
assign a17042 = ~a17040 & ~a16310;
assign a17044 = a12366 & l1462;
assign a17046 = ~a12366 & l1464;
assign a17048 = ~a17046 & ~a17044;
assign a17050 = ~a17048 & a16310;
assign a17052 = ~a17050 & ~a17042;
assign a17054 = ~a17052 & ~a16304;
assign a17056 = ~a14050 & a12366;
assign a17058 = ~a14058 & ~a12366;
assign a17060 = ~a17058 & ~a17056;
assign a17062 = ~a17060 & ~a16310;
assign a17064 = a12366 & l1470;
assign a17066 = ~a12366 & l1472;
assign a17068 = ~a17066 & ~a17064;
assign a17070 = ~a17068 & a16310;
assign a17072 = ~a17070 & ~a17062;
assign a17074 = ~a17072 & a16304;
assign a17076 = ~a17074 & ~a17054;
assign a17078 = ~a17076 & a16298;
assign a17080 = a16358 & l1472;
assign a17082 = ~a17080 & ~a17078;
assign a17084 = a12366 & l1454;
assign a17086 = ~a12366 & l1456;
assign a17088 = ~a17086 & ~a17084;
assign a17090 = ~a17088 & a16366;
assign a17092 = ~a17090 & a17082;
assign a17094 = ~a17092 & a16444;
assign a17096 = ~a16444 & ~a14098;
assign a17098 = ~a17096 & ~a17094;
assign a17100 = ~a16222 & l1144;
assign a17102 = a16196 & l1140;
assign a17104 = a9060 & l1142;
assign a17106 = ~a9060 & l1138;
assign a17108 = ~a17106 & ~a17104;
assign a17110 = ~a17108 & ~a16196;
assign a17112 = ~a17110 & ~a17102;
assign a17114 = ~a17112 & ~a16254;
assign a17116 = a16254 & l1140;
assign a17118 = ~a17116 & ~a17114;
assign a17120 = ~a17118 & a16222;
assign a17122 = ~a17120 & ~a17100;
assign a17124 = ~a17122 & a17098;
assign a17126 = ~a17124 & ~a17034;
assign a17128 = a17122 & ~a17098;
assign a17130 = ~a17128 & ~a17126;
assign a17132 = ~a17130 & a16456;
assign a17134 = ~a16520 & a16264;
assign a17136 = ~a17134 & ~a16624;
assign a17138 = ~a17136 & ~a16620;
assign a17140 = ~a17138 & ~a16728;
assign a17142 = ~a17140 & ~a16724;
assign a17144 = ~a17142 & ~a16832;
assign a17146 = ~a17144 & ~a16828;
assign a17148 = ~a17146 & ~a16936;
assign a17150 = ~a17148 & ~a16932;
assign a17152 = ~a17150 & ~a17032;
assign a17154 = ~a17152 & ~a17028;
assign a17156 = ~a17154 & ~a17128;
assign a17158 = ~a17156 & ~a17124;
assign a17160 = ~a17158 & ~a16456;
assign a17162 = ~a17160 & ~a17132;
assign a17164 = ~a17162 & ~a16264;
assign a17166 = a17162 & ~a16520;
assign a17168 = ~a17166 & ~a17164;
assign a17170 = ~a17168 & ~i246;
assign a17172 = ~a17162 & ~a16618;
assign a17174 = a17162 & ~a16586;
assign a17176 = ~a17174 & ~a17172;
assign a17178 = ~a17176 & ~i286;
assign a17180 = ~a17178 & ~a17170;
assign a17182 = a17176 & i286;
assign a17184 = ~a17182 & ~a17180;
assign a17186 = ~a17162 & ~a16722;
assign a17188 = a17162 & ~a16690;
assign a17190 = ~a17188 & ~a17186;
assign a17192 = ~a17190 & ~i288;
assign a17194 = ~a17192 & ~a17184;
assign a17196 = a17190 & i288;
assign a17198 = ~a17196 & ~a17194;
assign a17200 = ~a17162 & ~a16826;
assign a17202 = a17162 & ~a16794;
assign a17204 = ~a17202 & ~a17200;
assign a17206 = ~a17204 & ~i290;
assign a17208 = ~a17206 & ~a17198;
assign a17210 = a17204 & i290;
assign a17212 = ~a17210 & ~a17208;
assign a17214 = ~a17162 & ~a16930;
assign a17216 = a17162 & ~a16898;
assign a17218 = ~a17216 & ~a17214;
assign a17220 = ~a17218 & ~i292;
assign a17222 = ~a17220 & ~a17212;
assign a17224 = a17218 & i292;
assign a17226 = ~a17224 & ~a17222;
assign a17228 = ~a17162 & ~a17026;
assign a17230 = a17162 & ~a17002;
assign a17232 = ~a17230 & ~a17228;
assign a17234 = ~a17232 & ~i294;
assign a17236 = ~a17234 & ~a17226;
assign a17238 = a17232 & i294;
assign a17240 = ~a17238 & ~a17236;
assign a17242 = ~a17162 & ~a17122;
assign a17244 = a17162 & ~a17098;
assign a17246 = ~a17244 & ~a17242;
assign a17248 = ~a17246 & ~i296;
assign a17250 = ~a17248 & ~a17240;
assign a17252 = a17246 & i296;
assign a17254 = ~a17252 & ~a17250;
assign a17256 = ~a17162 & ~a16288;
assign a17258 = a17162 & ~a16450;
assign a17260 = ~a17258 & ~a17256;
assign a17262 = ~l974 & l890;
assign a17264 = ~a2712 & i238;
assign a17266 = ~a17264 & ~l890;
assign a17268 = ~a17266 & ~a17262;
assign a17270 = a17268 & l976;
assign a17272 = a17270 & ~l886;
assign a17274 = l1026 & ~l978;
assign a17276 = ~l1026 & l978;
assign a17278 = ~a17276 & ~a17274;
assign a17280 = ~l1030 & l890;
assign a17282 = ~a11250 & ~i276;
assign a17284 = a11250 & i276;
assign a17286 = ~a17284 & ~a17282;
assign a17288 = ~a17286 & a4144;
assign a17290 = ~a2712 & ~i276;
assign a17292 = ~a17290 & ~a17288;
assign a17294 = ~a17292 & ~l890;
assign a17296 = ~a17294 & ~a17280;
assign a17298 = a17296 & ~a6254;
assign a17300 = ~l1034 & l890;
assign a17302 = ~a11250 & i276;
assign a17304 = ~a11330 & ~i282;
assign a17306 = a11330 & i282;
assign a17308 = ~a17306 & ~a17304;
assign a17310 = ~a17308 & ~a17302;
assign a17312 = a17308 & a17302;
assign a17314 = ~a17312 & ~a17310;
assign a17316 = ~a17314 & a4144;
assign a17318 = i282 & ~i276;
assign a17320 = ~i282 & i276;
assign a17322 = ~a17320 & ~a17318;
assign a17324 = ~a17322 & ~a2712;
assign a17326 = ~a17324 & ~a17316;
assign a17328 = ~a17326 & ~l890;
assign a17330 = ~a17328 & ~a17300;
assign a17332 = a17330 & ~a6262;
assign a17334 = ~a17332 & ~a17298;
assign a17336 = ~a17330 & a6262;
assign a17338 = ~a17336 & ~a17334;
assign a17340 = ~l1062 & l890;
assign a17342 = ~a11330 & i282;
assign a17344 = ~a17342 & ~a17302;
assign a17346 = a11330 & ~i282;
assign a17348 = ~a17346 & ~a17344;
assign a17350 = ~a11372 & ~i298;
assign a17352 = a11372 & i298;
assign a17354 = ~a17352 & ~a17350;
assign a17356 = ~a17354 & ~a17348;
assign a17358 = a17354 & a17348;
assign a17360 = ~a17358 & ~a17356;
assign a17362 = ~a17360 & a4144;
assign a17364 = i282 & i276;
assign a17366 = ~a17364 & i298;
assign a17368 = a17364 & ~i298;
assign a17370 = ~a17368 & ~a17366;
assign a17372 = ~a17370 & ~a2712;
assign a17374 = ~a17372 & ~a17362;
assign a17376 = ~a17374 & ~l890;
assign a17378 = ~a17376 & ~a17340;
assign a17380 = a17378 & ~a6270;
assign a17382 = ~a17380 & ~a17338;
assign a17384 = ~a17378 & a6270;
assign a17386 = ~a17384 & ~a17382;
assign a17388 = ~l1068 & l890;
assign a17390 = a17364 & i298;
assign a17392 = a17390 & ~a2712;
assign a17394 = a17392 & ~l890;
assign a17396 = ~a17394 & ~a17388;
assign a17398 = a17396 & ~a6278;
assign a17400 = ~a17398 & ~a17386;
assign a17402 = ~a17396 & a6278;
assign a17404 = ~a17402 & ~a17400;
assign a17406 = ~a6286 & ~l1072;
assign a17408 = ~a17406 & ~a17404;
assign a17410 = a6286 & l1072;
assign a17412 = ~a17410 & ~a17408;
assign a17414 = ~l1076 & l1054;
assign a17416 = ~a17414 & ~a17412;
assign a17418 = l1076 & ~l1054;
assign a17420 = ~a17418 & ~a17416;
assign a17422 = l1058 & ~l1028;
assign a17424 = ~a17422 & ~a17420;
assign a17426 = ~l1058 & l1028;
assign a17428 = ~a17426 & ~a17424;
assign a17430 = a17428 & a17278;
assign a17432 = ~a17428 & ~a17278;
assign a17434 = ~a17432 & ~a17430;
assign a17436 = ~a17434 & a17272;
assign a17438 = a17272 & l1026;
assign a17440 = ~a17272 & i312;
assign a17442 = ~a17440 & ~a17438;
assign a17444 = ~a17442 & a17436;
assign a17446 = l978 & l886;
assign a17448 = l1766 & ~l886;
assign a17450 = ~a17448 & ~a17446;
assign a17452 = ~a17450 & ~a17436;
assign a17454 = ~a17452 & ~a17444;
assign a17456 = ~a17454 & a17260;
assign a17458 = a17454 & ~a17260;
assign a17460 = ~a17458 & ~a17456;
assign a17462 = ~a17296 & a17272;
assign a17464 = ~a17272 & i324;
assign a17466 = ~a17464 & ~a17462;
assign a17468 = ~a17466 & a17436;
assign a17470 = ~a6254 & l886;
assign a17472 = ~a17470 & ~l1152;
assign a17474 = ~a17472 & ~a17436;
assign a17476 = ~a17474 & ~a17468;
assign a17478 = a17476 & i246;
assign a17480 = ~a17330 & a17272;
assign a17482 = ~a17272 & i422;
assign a17484 = ~a17482 & ~a17480;
assign a17486 = ~a17484 & a17436;
assign a17488 = ~a6262 & l886;
assign a17490 = ~a17488 & ~l1768;
assign a17492 = ~a17490 & ~a17436;
assign a17494 = ~a17492 & ~a17486;
assign a17496 = a17494 & i286;
assign a17498 = ~a17496 & ~a17478;
assign a17500 = ~a17494 & ~i286;
assign a17502 = ~a17500 & ~a17498;
assign a17504 = ~a17378 & a17272;
assign a17506 = ~a17272 & i322;
assign a17508 = ~a17506 & ~a17504;
assign a17510 = ~a17508 & a17436;
assign a17512 = ~a6270 & l886;
assign a17514 = ~a17512 & ~l1770;
assign a17516 = ~a17514 & ~a17436;
assign a17518 = ~a17516 & ~a17510;
assign a17520 = a17518 & i288;
assign a17522 = ~a17520 & ~a17502;
assign a17524 = ~a17518 & ~i288;
assign a17526 = ~a17524 & ~a17522;
assign a17528 = ~a17396 & a17272;
assign a17530 = ~a17272 & i320;
assign a17532 = ~a17530 & ~a17528;
assign a17534 = ~a17532 & a17436;
assign a17536 = ~a6278 & l886;
assign a17538 = ~a17536 & ~l1772;
assign a17540 = ~a17538 & ~a17436;
assign a17542 = ~a17540 & ~a17534;
assign a17544 = a17542 & i290;
assign a17546 = ~a17544 & ~a17526;
assign a17548 = ~a17542 & ~i290;
assign a17550 = ~a17548 & ~a17546;
assign a17552 = a17272 & l1072;
assign a17554 = ~a17272 & i318;
assign a17556 = ~a17554 & ~a17552;
assign a17558 = ~a17556 & a17436;
assign a17560 = ~a6286 & l886;
assign a17562 = ~a17560 & ~l1774;
assign a17564 = ~a17562 & ~a17436;
assign a17566 = ~a17564 & ~a17558;
assign a17568 = a17566 & i292;
assign a17570 = ~a17568 & ~a17550;
assign a17572 = ~a17566 & ~i292;
assign a17574 = ~a17572 & ~a17570;
assign a17576 = a17272 & l1076;
assign a17578 = ~a17272 & i316;
assign a17580 = ~a17578 & ~a17576;
assign a17582 = ~a17580 & a17436;
assign a17584 = l1054 & l886;
assign a17586 = l1776 & ~l886;
assign a17588 = ~a17586 & ~a17584;
assign a17590 = ~a17588 & ~a17436;
assign a17592 = ~a17590 & ~a17582;
assign a17594 = a17592 & i294;
assign a17596 = ~a17594 & ~a17574;
assign a17598 = ~a17592 & ~i294;
assign a17600 = ~a17598 & ~a17596;
assign a17602 = a17272 & l1028;
assign a17604 = ~a17272 & i314;
assign a17606 = ~a17604 & ~a17602;
assign a17608 = ~a17606 & a17436;
assign a17610 = l1058 & l886;
assign a17612 = ~a17610 & ~l1778;
assign a17614 = ~a17612 & ~a17436;
assign a17616 = ~a17614 & ~a17608;
assign a17618 = a17616 & i296;
assign a17620 = ~a17618 & ~a17600;
assign a17622 = ~a17616 & ~i296;
assign a17624 = ~a17622 & ~a17620;
assign a17626 = a17454 & i242;
assign a17628 = ~a17454 & ~i242;
assign a17630 = ~a17628 & ~a17626;
assign a17632 = a17630 & a17624;
assign a17634 = a17632 & a17460;
assign a17636 = a17634 & a17254;
assign a17638 = a17260 & i242;
assign a17640 = ~a17260 & ~i242;
assign a17642 = ~a17640 & ~a17638;
assign a17644 = a17642 & a17254;
assign a17646 = ~a17644 & ~a17632;
assign a17648 = ~a17646 & ~a17460;
assign a17650 = ~a17648 & ~a17636;
assign a17652 = ~a17650 & ~a5360;
assign a17654 = a17652 & a16226;
assign a17656 = a17654 & a5562;
assign a17658 = a17656 & a16228;
assign a17660 = ~l2068 & l890;
assign a17662 = ~a5346 & i544;
assign a17664 = a17662 & ~a2706;
assign a17666 = a17664 & ~a5178;
assign a17668 = ~a17666 & ~l890;
assign a17670 = ~a17668 & ~a17660;
assign a17672 = a17670 & ~a17658;
assign a17674 = a17672 & ~a14378;
assign a17676 = a17674 & a16226;
assign a17678 = a17676 & a16222;
assign a17680 = a17678 & a16190;
assign a17684 = ~a5562 & l1194;
assign a17686 = ~a9048 & ~l1196;
assign a17688 = ~a12354 & ~l1252;
assign a17690 = a12354 & l1252;
assign a17692 = ~a12300 & ~l1260;
assign a17694 = a12300 & l1260;
assign a17696 = ~a12238 & ~l1266;
assign a17698 = a12238 & l1266;
assign a17700 = ~a12178 & ~l1272;
assign a17702 = a12178 & l1272;
assign a17704 = ~a17702 & ~a17700;
assign a17706 = a17704 & ~a17698;
assign a17708 = a17706 & ~a17696;
assign a17710 = a17708 & ~a17694;
assign a17712 = a17710 & ~a17692;
assign a17714 = a17712 & ~a17690;
assign a17716 = a17714 & ~a17688;
assign a17718 = ~a17716 & a17686;
assign a17720 = ~a17718 & i488;
assign a17722 = a17718 & l1278;
assign a17724 = ~a17722 & ~a17720;
assign a17726 = ~a17724 & a5562;
assign a17728 = ~a17726 & ~a17684;
assign a17730 = a16356 & a12312;
assign a17732 = ~a12366 & l1314;
assign a17734 = a12366 & l1316;
assign a17736 = ~a17734 & ~a17732;
assign a17738 = ~a17736 & a17730;
assign a17740 = ~a12366 & l1318;
assign a17742 = a12366 & l1320;
assign a17744 = ~a17742 & ~a17740;
assign a17746 = ~a17744 & ~a12312;
assign a17748 = ~a12366 & l1322;
assign a17750 = a12366 & l1324;
assign a17752 = ~a17750 & ~a17748;
assign a17754 = ~a17752 & a12312;
assign a17756 = ~a17754 & ~a17746;
assign a17758 = ~a17756 & ~a12250;
assign a17760 = ~a12366 & l1326;
assign a17762 = a12366 & l1328;
assign a17764 = ~a17762 & ~a17760;
assign a17766 = ~a17764 & ~a12312;
assign a17768 = ~a12366 & l1330;
assign a17770 = a12366 & l1332;
assign a17772 = ~a17770 & ~a17768;
assign a17774 = ~a17772 & a12312;
assign a17776 = ~a17774 & ~a17766;
assign a17778 = ~a17776 & a12250;
assign a17780 = ~a17778 & ~a17758;
assign a17782 = ~a17780 & a12190;
assign a17784 = ~a17782 & ~a17738;
assign a17786 = a17784 & ~a17728;
assign a17788 = ~a17784 & a17728;
assign a17790 = ~a17788 & ~a17786;
assign a17792 = ~a12366 & l1334;
assign a17794 = a12366 & l1336;
assign a17796 = ~a17794 & ~a17792;
assign a17798 = ~a17796 & a17730;
assign a17800 = ~a12366 & l1338;
assign a17802 = a12366 & l1340;
assign a17804 = ~a17802 & ~a17800;
assign a17806 = ~a17804 & ~a12312;
assign a17808 = ~a12366 & l1342;
assign a17810 = a12366 & l1344;
assign a17812 = ~a17810 & ~a17808;
assign a17814 = ~a17812 & a12312;
assign a17816 = ~a17814 & ~a17806;
assign a17818 = ~a17816 & ~a12250;
assign a17820 = ~a12954 & ~a12366;
assign a17822 = ~a12962 & a12366;
assign a17824 = ~a17822 & ~a17820;
assign a17826 = ~a17824 & ~a12312;
assign a17828 = ~a12974 & ~a12366;
assign a17830 = a12366 & l1352;
assign a17832 = ~a17830 & ~a17828;
assign a17834 = ~a17832 & a12312;
assign a17836 = ~a17834 & ~a17826;
assign a17838 = ~a17836 & a12250;
assign a17840 = ~a17838 & ~a17818;
assign a17842 = ~a17840 & a12190;
assign a17844 = ~a17842 & ~a17798;
assign a17846 = ~a5562 & l1306;
assign a17848 = ~a17718 & i490;
assign a17850 = a17718 & ~a10652;
assign a17852 = ~a17850 & ~a17848;
assign a17854 = ~a17852 & a5562;
assign a17856 = ~a17854 & ~a17846;
assign a17858 = a17856 & ~a17844;
assign a17860 = ~a12366 & l1354;
assign a17862 = a12366 & l1356;
assign a17864 = ~a17862 & ~a17860;
assign a17866 = ~a17864 & a17730;
assign a17868 = ~a12366 & l1358;
assign a17870 = a12366 & l1360;
assign a17872 = ~a17870 & ~a17868;
assign a17874 = ~a17872 & ~a12312;
assign a17876 = ~a12366 & l1362;
assign a17878 = a12366 & l1364;
assign a17880 = ~a17878 & ~a17876;
assign a17882 = ~a17880 & a12312;
assign a17884 = ~a17882 & ~a17874;
assign a17886 = ~a17884 & ~a12250;
assign a17888 = ~a13138 & ~a12366;
assign a17890 = ~a13146 & a12366;
assign a17892 = ~a17890 & ~a17888;
assign a17894 = ~a17892 & ~a12312;
assign a17896 = ~a13158 & ~a12366;
assign a17898 = a12366 & l1372;
assign a17900 = ~a17898 & ~a17896;
assign a17902 = ~a17900 & a12312;
assign a17904 = ~a17902 & ~a17894;
assign a17906 = ~a17904 & a12250;
assign a17908 = ~a17906 & ~a17886;
assign a17910 = ~a17908 & a12190;
assign a17912 = ~a17910 & ~a17866;
assign a17914 = ~a5562 & l1302;
assign a17916 = ~a17718 & i492;
assign a17918 = a17718 & ~a10592;
assign a17920 = ~a17918 & ~a17916;
assign a17922 = ~a17920 & a5562;
assign a17924 = ~a17922 & ~a17914;
assign a17926 = a17924 & ~a17912;
assign a17928 = ~a17926 & ~a17858;
assign a17930 = ~a17924 & a17912;
assign a17932 = ~a17930 & ~a17928;
assign a17934 = ~a12366 & l1374;
assign a17936 = a12366 & l1376;
assign a17938 = ~a17936 & ~a17934;
assign a17940 = ~a17938 & a17730;
assign a17942 = ~a12366 & l1378;
assign a17944 = a12366 & l1380;
assign a17946 = ~a17944 & ~a17942;
assign a17948 = ~a17946 & ~a12312;
assign a17950 = ~a12366 & l1382;
assign a17952 = a12366 & l1384;
assign a17954 = ~a17952 & ~a17950;
assign a17956 = ~a17954 & a12312;
assign a17958 = ~a17956 & ~a17948;
assign a17960 = ~a17958 & ~a12250;
assign a17962 = ~a13328 & ~a12366;
assign a17964 = ~a13336 & a12366;
assign a17966 = ~a17964 & ~a17962;
assign a17968 = ~a17966 & ~a12312;
assign a17970 = ~a13348 & ~a12366;
assign a17972 = a12366 & l1392;
assign a17974 = ~a17972 & ~a17970;
assign a17976 = ~a17974 & a12312;
assign a17978 = ~a17976 & ~a17968;
assign a17980 = ~a17978 & a12250;
assign a17982 = ~a17980 & ~a17960;
assign a17984 = ~a17982 & a12190;
assign a17986 = ~a17984 & ~a17940;
assign a17988 = ~a5562 & l1298;
assign a17990 = ~a17718 & i494;
assign a17992 = a17718 & ~a10556;
assign a17994 = ~a17992 & ~a17990;
assign a17996 = ~a17994 & a5562;
assign a17998 = ~a17996 & ~a17988;
assign a18000 = a17998 & ~a17986;
assign a18002 = ~a18000 & ~a17932;
assign a18004 = ~a17998 & a17986;
assign a18006 = ~a18004 & ~a18002;
assign a18008 = ~a12366 & l1394;
assign a18010 = a12366 & l1396;
assign a18012 = ~a18010 & ~a18008;
assign a18014 = ~a18012 & a17730;
assign a18016 = ~a12366 & l1398;
assign a18018 = a12366 & l1400;
assign a18020 = ~a18018 & ~a18016;
assign a18022 = ~a18020 & ~a12312;
assign a18024 = ~a12366 & l1402;
assign a18026 = a12366 & l1404;
assign a18028 = ~a18026 & ~a18024;
assign a18030 = ~a18028 & a12312;
assign a18032 = ~a18030 & ~a18022;
assign a18034 = ~a18032 & ~a12250;
assign a18036 = ~a13518 & ~a12366;
assign a18038 = ~a13526 & a12366;
assign a18040 = ~a18038 & ~a18036;
assign a18042 = ~a18040 & ~a12312;
assign a18044 = ~a13538 & ~a12366;
assign a18046 = a12366 & l1412;
assign a18048 = ~a18046 & ~a18044;
assign a18050 = ~a18048 & a12312;
assign a18052 = ~a18050 & ~a18042;
assign a18054 = ~a18052 & a12250;
assign a18056 = ~a18054 & ~a18034;
assign a18058 = ~a18056 & a12190;
assign a18060 = ~a18058 & ~a18014;
assign a18062 = ~a5562 & l1294;
assign a18064 = ~a17718 & i496;
assign a18066 = a17718 & ~a10520;
assign a18068 = ~a18066 & ~a18064;
assign a18070 = ~a18068 & a5562;
assign a18072 = ~a18070 & ~a18062;
assign a18074 = a18072 & ~a18060;
assign a18076 = ~a18074 & ~a18006;
assign a18078 = ~a18072 & a18060;
assign a18080 = ~a18078 & ~a18076;
assign a18082 = ~a12366 & l1414;
assign a18084 = a12366 & l1416;
assign a18086 = ~a18084 & ~a18082;
assign a18088 = ~a18086 & a17730;
assign a18090 = ~a12366 & l1418;
assign a18092 = a12366 & l1420;
assign a18094 = ~a18092 & ~a18090;
assign a18096 = ~a18094 & ~a12312;
assign a18098 = ~a12366 & l1422;
assign a18100 = a12366 & l1424;
assign a18102 = ~a18100 & ~a18098;
assign a18104 = ~a18102 & a12312;
assign a18106 = ~a18104 & ~a18096;
assign a18108 = ~a18106 & ~a12250;
assign a18110 = ~a13708 & ~a12366;
assign a18112 = ~a13716 & a12366;
assign a18114 = ~a18112 & ~a18110;
assign a18116 = ~a18114 & ~a12312;
assign a18118 = ~a13728 & ~a12366;
assign a18120 = a12366 & l1432;
assign a18122 = ~a18120 & ~a18118;
assign a18124 = ~a18122 & a12312;
assign a18126 = ~a18124 & ~a18116;
assign a18128 = ~a18126 & a12250;
assign a18130 = ~a18128 & ~a18108;
assign a18132 = ~a18130 & a12190;
assign a18134 = ~a18132 & ~a18088;
assign a18136 = ~a5562 & l1290;
assign a18138 = ~a17718 & i498;
assign a18140 = a17718 & ~a10484;
assign a18142 = ~a18140 & ~a18138;
assign a18144 = ~a18142 & a5562;
assign a18146 = ~a18144 & ~a18136;
assign a18148 = a18146 & ~a18134;
assign a18150 = ~a18148 & ~a18080;
assign a18152 = ~a18146 & a18134;
assign a18154 = ~a18152 & ~a18150;
assign a18156 = ~a12366 & l1434;
assign a18158 = a12366 & l1436;
assign a18160 = ~a18158 & ~a18156;
assign a18162 = ~a18160 & a17730;
assign a18164 = ~a12366 & l1438;
assign a18166 = a12366 & l1440;
assign a18168 = ~a18166 & ~a18164;
assign a18170 = ~a18168 & ~a12312;
assign a18172 = ~a12366 & l1442;
assign a18174 = a12366 & l1444;
assign a18176 = ~a18174 & ~a18172;
assign a18178 = ~a18176 & a12312;
assign a18180 = ~a18178 & ~a18170;
assign a18182 = ~a18180 & ~a12250;
assign a18184 = ~a13886 & ~a12366;
assign a18186 = ~a13894 & a12366;
assign a18188 = ~a18186 & ~a18184;
assign a18190 = ~a18188 & ~a12312;
assign a18192 = ~a13906 & ~a12366;
assign a18194 = a12366 & l1452;
assign a18196 = ~a18194 & ~a18192;
assign a18198 = ~a18196 & a12312;
assign a18200 = ~a18198 & ~a18190;
assign a18202 = ~a18200 & a12250;
assign a18204 = ~a18202 & ~a18182;
assign a18206 = ~a18204 & a12190;
assign a18208 = ~a18206 & ~a18162;
assign a18210 = ~a5562 & l1286;
assign a18212 = ~a17718 & i500;
assign a18214 = a17718 & ~a9072;
assign a18216 = ~a18214 & ~a18212;
assign a18218 = ~a18216 & a5562;
assign a18220 = ~a18218 & ~a18210;
assign a18222 = a18220 & ~a18208;
assign a18224 = ~a18222 & ~a18154;
assign a18226 = ~a18220 & a18208;
assign a18228 = ~a18226 & ~a18224;
assign a18230 = ~a12366 & l1454;
assign a18232 = a12366 & l1456;
assign a18234 = ~a18232 & ~a18230;
assign a18236 = ~a18234 & a17730;
assign a18238 = ~a12366 & l1458;
assign a18240 = a12366 & l1460;
assign a18242 = ~a18240 & ~a18238;
assign a18244 = ~a18242 & ~a12312;
assign a18246 = ~a12366 & l1462;
assign a18248 = a12366 & l1464;
assign a18250 = ~a18248 & ~a18246;
assign a18252 = ~a18250 & a12312;
assign a18254 = ~a18252 & ~a18244;
assign a18256 = ~a18254 & ~a12250;
assign a18258 = ~a14050 & ~a12366;
assign a18260 = ~a14058 & a12366;
assign a18262 = ~a18260 & ~a18258;
assign a18264 = ~a18262 & ~a12312;
assign a18266 = ~a12366 & l1470;
assign a18268 = a12366 & l1472;
assign a18270 = ~a18268 & ~a18266;
assign a18272 = ~a18270 & a12312;
assign a18274 = ~a18272 & ~a18264;
assign a18276 = ~a18274 & a12250;
assign a18278 = ~a18276 & ~a18256;
assign a18280 = ~a18278 & a12190;
assign a18282 = ~a18280 & ~a18236;
assign a18284 = ~a5562 & l1282;
assign a18286 = ~a17718 & i502;
assign a18288 = a17718 & l1280;
assign a18290 = ~a18288 & ~a18286;
assign a18292 = ~a18290 & a5562;
assign a18294 = ~a18292 & ~a18284;
assign a18296 = a18294 & ~a18282;
assign a18298 = ~a18296 & ~a18228;
assign a18300 = ~a18294 & a18282;
assign a18302 = ~a18300 & ~a18298;
assign a18304 = ~a18302 & a17790;
assign a18306 = a18302 & ~a17790;
assign a18308 = ~a18306 & ~a18304;
assign a18310 = ~a12354 & a12328;
assign a18312 = a12354 & ~a12328;
assign a18314 = ~a12300 & a12268;
assign a18316 = a12300 & ~a12268;
assign a18318 = ~a12238 & a12206;
assign a18320 = a12238 & ~a12206;
assign a18322 = ~a12178 & a9026;
assign a18324 = a12178 & ~a9026;
assign a18326 = ~a18324 & ~a18322;
assign a18328 = a18326 & ~a18320;
assign a18330 = a18328 & ~a18318;
assign a18332 = a18330 & ~a18316;
assign a18334 = a18332 & ~a18314;
assign a18336 = a18334 & ~a18312;
assign a18338 = a18336 & ~a18310;
assign a18340 = ~a17728 & a16376;
assign a18342 = a17728 & ~a16376;
assign a18344 = ~a18342 & ~a18340;
assign a18346 = a17856 & ~a16514;
assign a18348 = a17924 & ~a16580;
assign a18350 = ~a18348 & ~a18346;
assign a18352 = ~a17924 & a16580;
assign a18354 = ~a18352 & ~a18350;
assign a18356 = a17998 & ~a16684;
assign a18358 = ~a18356 & ~a18354;
assign a18360 = ~a17998 & a16684;
assign a18362 = ~a18360 & ~a18358;
assign a18364 = a18072 & ~a16788;
assign a18366 = ~a18364 & ~a18362;
assign a18368 = ~a18072 & a16788;
assign a18370 = ~a18368 & ~a18366;
assign a18372 = a18146 & ~a16892;
assign a18374 = ~a18372 & ~a18370;
assign a18376 = ~a18146 & a16892;
assign a18378 = ~a18376 & ~a18374;
assign a18380 = a18220 & ~a16996;
assign a18382 = ~a18380 & ~a18378;
assign a18384 = ~a18220 & a16996;
assign a18386 = ~a18384 & ~a18382;
assign a18388 = a18294 & ~a17092;
assign a18390 = ~a18388 & ~a18386;
assign a18392 = ~a18294 & a17092;
assign a18394 = ~a18392 & ~a18390;
assign a18396 = a18394 & a18344;
assign a18398 = ~a18394 & ~a18344;
assign a18400 = ~a18398 & ~a18396;
assign a18402 = ~a18400 & ~a18338;
assign a18404 = ~a17728 & a12824;
assign a18406 = a17728 & ~a12824;
assign a18408 = ~a18406 & ~a18404;
assign a18410 = a17856 & ~a13012;
assign a18412 = a17924 & ~a13196;
assign a18414 = ~a18412 & ~a18410;
assign a18416 = ~a17924 & a13196;
assign a18418 = ~a18416 & ~a18414;
assign a18420 = a17998 & ~a13386;
assign a18422 = ~a18420 & ~a18418;
assign a18424 = ~a17998 & a13386;
assign a18426 = ~a18424 & ~a18422;
assign a18428 = a18072 & ~a13576;
assign a18430 = ~a18428 & ~a18426;
assign a18432 = ~a18072 & a13576;
assign a18434 = ~a18432 & ~a18430;
assign a18436 = a18146 & ~a13766;
assign a18438 = ~a18436 & ~a18434;
assign a18440 = ~a18146 & a13766;
assign a18442 = ~a18440 & ~a18438;
assign a18444 = a18220 & ~a13944;
assign a18446 = ~a18444 & ~a18442;
assign a18448 = ~a18220 & a13944;
assign a18450 = ~a18448 & ~a18446;
assign a18452 = a18294 & ~a14102;
assign a18454 = ~a18452 & ~a18450;
assign a18456 = ~a18294 & a14102;
assign a18458 = ~a18456 & ~a18454;
assign a18460 = a18458 & a18408;
assign a18462 = ~a18458 & ~a18408;
assign a18464 = ~a18462 & ~a18460;
assign a18466 = ~a18464 & a18338;
assign a18468 = ~a18466 & ~a18402;
assign a18470 = ~a18468 & ~a18308;
assign a18472 = a18470 & a5562;
assign a18474 = a18472 & i158;
assign a18476 = a12160 & a12138;
assign a18478 = ~a12160 & a12142;
assign a18480 = ~a18478 & ~a18476;
assign a18482 = ~a18480 & ~a12116;
assign a18484 = a12160 & ~a12150;
assign a18486 = a12160 & a12142;
assign a18488 = ~a18486 & ~a18484;
assign a18490 = ~a18488 & a5562;
assign a18492 = ~a18490 & a18480;
assign a18494 = a18492 & ~a18482;
assign a18496 = a18494 & i504;
assign a18498 = ~a18496 & ~a18482;
assign a18500 = a18498 & ~a17718;
assign a18502 = a18500 & ~a18474;
assign a18504 = ~l1102 & ~l908;
assign a18506 = a18504 & ~a18502;
assign a18508 = a18506 & a12110;
assign a18510 = a18508 & ~a9064;
assign a18512 = ~a18510 & l910;
assign a18516 = a16218 & l990;
assign a18518 = ~a18516 & ~a18512;
assign a18522 = a18514 & i508;
assign a18524 = ~a18522 & ~a9048;
assign a18526 = a18524 & ~l892;
assign a18528 = ~l2064 & l890;
assign a18530 = a4142 & ~l890;
assign a18532 = ~a18530 & ~a18528;
assign a18534 = ~l2066 & ~l1190;
assign a18536 = a18534 & a18532;
assign a18538 = ~a18536 & ~a12110;
assign a18540 = ~a18538 & ~l886;
assign a18544 = ~a16190 & ~a9038;
assign a18546 = a14378 & i506;
assign a18548 = a18546 & a16198;
assign a18550 = ~a18548 & ~a9038;
assign a18552 = ~a18550 & a16190;
assign a18554 = ~a18552 & ~a18544;
assign a18558 = ~a18508 & ~a5562;
assign a18560 = ~a18558 & a17686;
assign a18564 = ~l922 & l890;
assign a18566 = a2710 & ~l890;
assign a18568 = ~a18566 & ~a18564;
assign a18570 = ~l1006 & ~l1004;
assign a18572 = a18570 & ~l1002;
assign a18574 = a18572 & a18568;
assign a18576 = a18574 & l880;
assign a18578 = ~l1954 & l890;
assign a18580 = a2712 & ~l890;
assign a18582 = ~a18580 & ~a18578;
assign a18584 = a18582 & ~l1002;
assign a18586 = a18570 & ~l880;
assign a18588 = a18586 & a18584;
assign a18590 = ~a18588 & ~a18576;
assign a18592 = ~l1972 & l890;
assign a18594 = ~a2722 & ~l890;
assign a18596 = ~a18594 & ~a18592;
assign a18598 = ~l1006 & ~l1002;
assign a18600 = a18598 & a18596;
assign a18602 = a18600 & a2746;
assign a18604 = ~a18602 & a18590;
assign a18606 = ~l1006 & l1004;
assign a18608 = a18606 & ~l1002;
assign a18610 = a18608 & l1974;
assign a18612 = a18610 & l880;
assign a18614 = ~a18612 & a18604;
assign a18616 = l1976 & ~l1006;
assign a18618 = a2530 & ~l880;
assign a18620 = a18618 & a18616;
assign a18622 = ~a18620 & a18614;
assign a18624 = a2530 & l1978;
assign a18626 = a18624 & l880;
assign a18628 = ~a18626 & a18622;
assign a18630 = ~l1006 & l1002;
assign a18632 = a18630 & l1980;
assign a18634 = a18632 & a2746;
assign a18636 = ~a18634 & a18628;
assign a18638 = a18606 & l1002;
assign a18640 = a18638 & l1982;
assign a18642 = a18640 & l880;
assign a18644 = ~a18642 & a18636;
assign a18646 = l1984 & ~l884;
assign a18648 = l1006 & ~l1002;
assign a18650 = a18648 & ~l880;
assign a18652 = a18650 & a18646;
assign a18654 = ~a18652 & a18644;
assign a18656 = a18648 & l1986;
assign a18658 = a18656 & l880;
assign a18660 = ~a18658 & a18654;
assign a18662 = a18574 & ~l880;
assign a18664 = l1006 & l880;
assign a18666 = a18664 & a18584;
assign a18668 = ~a18666 & ~a18662;
assign a18670 = ~l1004 & l880;
assign a18672 = a18670 & a18600;
assign a18674 = ~a18672 & a18668;
assign a18676 = a18610 & ~l880;
assign a18678 = ~a18676 & a18674;
assign a18680 = a18616 & a2526;
assign a18682 = ~a18680 & a18678;
assign a18684 = a18624 & ~l880;
assign a18686 = ~a18684 & a18682;
assign a18688 = a18670 & a18632;
assign a18690 = ~a18688 & a18686;
assign a18692 = a18640 & ~l880;
assign a18694 = ~a18692 & a18690;
assign a18696 = a18638 & l880;
assign a18698 = a18696 & a18646;
assign a18700 = ~a18698 & a18694;
assign a18702 = a18656 & ~l880;
assign a18704 = ~a18702 & a18700;
assign a18706 = ~a18704 & ~a18660;
assign a18708 = ~l1244 & l1006;
assign a18710 = l1244 & ~l1006;
assign a18712 = ~a18710 & ~a18708;
assign a18714 = l1156 & ~l1002;
assign a18716 = ~a18714 & a18712;
assign a18718 = ~l1156 & l1002;
assign a18720 = ~a18718 & a18716;
assign a18722 = ~a2740 & ~l1004;
assign a18724 = ~a18722 & a18720;
assign a18726 = a2740 & l1004;
assign a18728 = ~a18726 & a18724;
assign a18730 = ~a2768 & ~l880;
assign a18732 = ~a18730 & a18728;
assign a18734 = a2768 & l880;
assign a18736 = ~a18734 & a18732;
assign a18738 = ~a18736 & a18706;
assign a18740 = ~a18738 & ~a18660;
assign a18742 = ~a17658 & l2062;
assign a18744 = ~a18742 & ~a5360;
assign a18746 = a18572 & l1932;
assign a18748 = a18746 & ~l880;
assign a18750 = l1936 & ~l1002;
assign a18752 = a18750 & a18664;
assign a18754 = ~a18752 & ~a18748;
assign a18756 = a18598 & l1938;
assign a18758 = a18756 & a18670;
assign a18760 = ~a18758 & a18754;
assign a18762 = a18608 & l1940;
assign a18764 = a18762 & ~l880;
assign a18766 = ~a18764 & a18760;
assign a18768 = l1942 & ~l1006;
assign a18770 = a18768 & a2526;
assign a18772 = ~a18770 & a18766;
assign a18774 = a2530 & l1944;
assign a18776 = a18774 & ~l880;
assign a18778 = ~a18776 & a18772;
assign a18780 = a18630 & l1946;
assign a18782 = a18780 & a18670;
assign a18784 = ~a18782 & a18778;
assign a18786 = a18638 & l1948;
assign a18788 = a18786 & ~l880;
assign a18790 = ~a18788 & a18784;
assign a18792 = a18696 & l1950;
assign a18794 = ~a18792 & a18790;
assign a18796 = a18650 & l1952;
assign a18798 = ~a18796 & a18794;
assign a18800 = a18746 & l880;
assign a18802 = a18750 & a18586;
assign a18804 = ~a18802 & ~a18800;
assign a18806 = a18756 & a2746;
assign a18808 = ~a18806 & a18804;
assign a18810 = a18762 & l880;
assign a18812 = ~a18810 & a18808;
assign a18814 = a18768 & a18618;
assign a18816 = ~a18814 & a18812;
assign a18818 = a18774 & l880;
assign a18820 = ~a18818 & a18816;
assign a18822 = a18780 & a2746;
assign a18824 = ~a18822 & a18820;
assign a18826 = a18786 & l880;
assign a18828 = ~a18826 & a18824;
assign a18830 = a18650 & l1950;
assign a18832 = ~a18830 & a18828;
assign a18834 = a18664 & ~l1002;
assign a18836 = a18834 & l1952;
assign a18838 = ~a18836 & a18832;
assign a18840 = ~a18838 & a18798;
assign a18842 = a18838 & ~a18798;
assign a18844 = ~a18842 & ~a18840;
assign a18846 = a17658 & i246;
assign a18848 = ~a17658 & ~a6254;
assign a18852 = ~l1780 & l890;
assign a18854 = ~a4108 & ~l890;
assign a18856 = ~a18854 & ~a18852;
assign a18858 = ~a18856 & a18572;
assign a18860 = a18858 & l880;
assign a18862 = l1784 & ~l1002;
assign a18864 = a18862 & a18586;
assign a18866 = ~a18864 & ~a18860;
assign a18868 = ~l1154 & l890;
assign a18870 = a11094 & ~l890;
assign a18872 = ~a18870 & ~a18868;
assign a18874 = ~a18872 & a18598;
assign a18876 = a18874 & a2746;
assign a18878 = ~a18876 & a18866;
assign a18880 = a18608 & l1786;
assign a18882 = a18880 & l880;
assign a18884 = ~a18882 & a18878;
assign a18886 = l1788 & ~l1006;
assign a18888 = a18886 & a18618;
assign a18890 = ~a18888 & a18884;
assign a18892 = a2530 & l1790;
assign a18894 = a18892 & l880;
assign a18896 = ~a18894 & a18890;
assign a18898 = a18630 & l1792;
assign a18900 = a18898 & a2746;
assign a18902 = ~a18900 & a18896;
assign a18904 = a18638 & l1794;
assign a18906 = a18904 & l880;
assign a18908 = ~a18906 & a18902;
assign a18910 = a18650 & l1796;
assign a18912 = ~a18910 & a18908;
assign a18914 = a18834 & l1798;
assign a18916 = ~a18914 & a18912;
assign a18918 = ~a18916 & a18850;
assign a18920 = a17658 & i286;
assign a18922 = ~a17658 & ~a6262;
assign a18926 = ~l1800 & l890;
assign a18928 = ~a4224 & ~l890;
assign a18930 = ~a18928 & ~a18926;
assign a18932 = ~a18930 & a18572;
assign a18934 = a18932 & l880;
assign a18936 = l1804 & ~l1002;
assign a18938 = a18936 & a18586;
assign a18940 = ~a18938 & ~a18934;
assign a18942 = ~l1806 & l890;
assign a18944 = a11108 & ~l890;
assign a18946 = ~a18944 & ~a18942;
assign a18948 = ~a18946 & a18598;
assign a18950 = a18948 & a2746;
assign a18952 = ~a18950 & a18940;
assign a18954 = a18608 & l1808;
assign a18956 = a18954 & l880;
assign a18958 = ~a18956 & a18952;
assign a18960 = l1810 & ~l1006;
assign a18962 = a18960 & a18618;
assign a18964 = ~a18962 & a18958;
assign a18966 = a2530 & l1812;
assign a18968 = a18966 & l880;
assign a18970 = ~a18968 & a18964;
assign a18972 = a18630 & l1814;
assign a18974 = a18972 & a2746;
assign a18976 = ~a18974 & a18970;
assign a18978 = a18638 & l1816;
assign a18980 = a18978 & l880;
assign a18982 = ~a18980 & a18976;
assign a18984 = a18650 & l1818;
assign a18986 = ~a18984 & a18982;
assign a18988 = a18834 & l1820;
assign a18990 = ~a18988 & a18986;
assign a18992 = ~a18990 & a18924;
assign a18994 = ~a18992 & ~a18918;
assign a18996 = a18990 & ~a18924;
assign a18998 = ~a18996 & ~a18994;
assign a19000 = a17658 & i288;
assign a19002 = ~a17658 & ~a6270;
assign a19006 = ~l1822 & l890;
assign a19008 = ~a4370 & ~l890;
assign a19010 = ~a19008 & ~a19006;
assign a19012 = ~a19010 & a18572;
assign a19014 = a19012 & l880;
assign a19016 = l1826 & ~l1002;
assign a19018 = a19016 & a18586;
assign a19020 = ~a19018 & ~a19014;
assign a19022 = ~l1828 & l890;
assign a19024 = a11128 & ~l890;
assign a19026 = ~a19024 & ~a19022;
assign a19028 = ~a19026 & a18598;
assign a19030 = a19028 & a2746;
assign a19032 = ~a19030 & a19020;
assign a19034 = a18608 & l1830;
assign a19036 = a19034 & l880;
assign a19038 = ~a19036 & a19032;
assign a19040 = l1832 & ~l1006;
assign a19042 = a19040 & a18618;
assign a19044 = ~a19042 & a19038;
assign a19046 = a2530 & l1834;
assign a19048 = a19046 & l880;
assign a19050 = ~a19048 & a19044;
assign a19052 = a18630 & l1836;
assign a19054 = a19052 & a2746;
assign a19056 = ~a19054 & a19050;
assign a19058 = a18638 & l1838;
assign a19060 = a19058 & l880;
assign a19062 = ~a19060 & a19056;
assign a19064 = a18650 & l1840;
assign a19066 = ~a19064 & a19062;
assign a19068 = a18648 & l1842;
assign a19070 = a19068 & l880;
assign a19072 = ~a19070 & a19066;
assign a19074 = ~a19072 & a19004;
assign a19076 = ~a19074 & ~a18998;
assign a19078 = a19072 & ~a19004;
assign a19080 = ~a19078 & ~a19076;
assign a19082 = a17658 & i290;
assign a19084 = ~a17658 & ~a6278;
assign a19088 = ~l1844 & l890;
assign a19090 = ~a4530 & ~l890;
assign a19092 = ~a19090 & ~a19088;
assign a19094 = ~a19092 & a18572;
assign a19096 = a19094 & l880;
assign a19098 = l1848 & ~l1002;
assign a19100 = a19098 & a18586;
assign a19102 = ~a19100 & ~a19096;
assign a19104 = ~l1850 & l890;
assign a19106 = a11148 & ~l890;
assign a19108 = ~a19106 & ~a19104;
assign a19110 = ~a19108 & a18598;
assign a19112 = a19110 & a2746;
assign a19114 = ~a19112 & a19102;
assign a19116 = a18608 & l1852;
assign a19118 = a19116 & l880;
assign a19120 = ~a19118 & a19114;
assign a19122 = l1854 & ~l1006;
assign a19124 = a19122 & a18618;
assign a19126 = ~a19124 & a19120;
assign a19128 = a2530 & l1856;
assign a19130 = a19128 & l880;
assign a19132 = ~a19130 & a19126;
assign a19134 = a18630 & l1858;
assign a19136 = a19134 & a2746;
assign a19138 = ~a19136 & a19132;
assign a19140 = a18638 & l1860;
assign a19142 = a19140 & l880;
assign a19144 = ~a19142 & a19138;
assign a19146 = a18650 & l1862;
assign a19148 = ~a19146 & a19144;
assign a19150 = a18648 & l1864;
assign a19152 = a19150 & l880;
assign a19154 = ~a19152 & a19148;
assign a19156 = ~a19154 & a19086;
assign a19158 = ~a19156 & ~a19080;
assign a19160 = a19154 & ~a19086;
assign a19162 = ~a19160 & ~a19158;
assign a19164 = a17658 & i292;
assign a19166 = ~a17658 & ~a6286;
assign a19170 = ~l1866 & l890;
assign a19172 = ~a4690 & ~l890;
assign a19174 = ~a19172 & ~a19170;
assign a19176 = ~a19174 & a18572;
assign a19178 = a19176 & l880;
assign a19180 = l1870 & ~l1002;
assign a19182 = a19180 & a18586;
assign a19184 = ~a19182 & ~a19178;
assign a19186 = ~l1872 & l890;
assign a19188 = a11168 & ~l890;
assign a19190 = ~a19188 & ~a19186;
assign a19192 = ~a19190 & a18598;
assign a19194 = a19192 & a2746;
assign a19196 = ~a19194 & a19184;
assign a19198 = a18608 & l1874;
assign a19200 = a19198 & l880;
assign a19202 = ~a19200 & a19196;
assign a19204 = l1876 & ~l1006;
assign a19206 = a19204 & a18618;
assign a19208 = ~a19206 & a19202;
assign a19210 = a2530 & l1878;
assign a19212 = a19210 & l880;
assign a19214 = ~a19212 & a19208;
assign a19216 = a18630 & l1880;
assign a19218 = a19216 & a2746;
assign a19220 = ~a19218 & a19214;
assign a19222 = a18638 & l1882;
assign a19224 = a19222 & l880;
assign a19226 = ~a19224 & a19220;
assign a19228 = a18650 & l1884;
assign a19230 = ~a19228 & a19226;
assign a19232 = a18648 & l1886;
assign a19234 = a19232 & l880;
assign a19236 = ~a19234 & a19230;
assign a19238 = ~a19236 & a19168;
assign a19240 = ~a19238 & ~a19162;
assign a19242 = a19236 & ~a19168;
assign a19244 = ~a19242 & ~a19240;
assign a19246 = a17658 & i294;
assign a19248 = ~a17658 & l1054;
assign a19250 = ~a19248 & ~a19246;
assign a19252 = ~l1888 & l890;
assign a19254 = ~a4832 & ~l890;
assign a19256 = ~a19254 & ~a19252;
assign a19258 = ~a19256 & a18572;
assign a19260 = a19258 & l880;
assign a19262 = l1892 & ~l1002;
assign a19264 = a19262 & a18586;
assign a19266 = ~a19264 & ~a19260;
assign a19268 = ~l1894 & l890;
assign a19270 = a11188 & ~l890;
assign a19272 = ~a19270 & ~a19268;
assign a19274 = ~a19272 & a18598;
assign a19276 = a19274 & a2746;
assign a19278 = ~a19276 & a19266;
assign a19280 = a18608 & l1896;
assign a19282 = a19280 & l880;
assign a19284 = ~a19282 & a19278;
assign a19286 = l1898 & ~l1006;
assign a19288 = a19286 & a18618;
assign a19290 = ~a19288 & a19284;
assign a19292 = a2530 & l1900;
assign a19294 = a19292 & l880;
assign a19296 = ~a19294 & a19290;
assign a19298 = a18630 & l1902;
assign a19300 = a19298 & a2746;
assign a19302 = ~a19300 & a19296;
assign a19304 = a18638 & l1904;
assign a19306 = a19304 & l880;
assign a19308 = ~a19306 & a19302;
assign a19310 = a18650 & l1906;
assign a19312 = ~a19310 & a19308;
assign a19314 = a18648 & l1908;
assign a19316 = a19314 & l880;
assign a19318 = ~a19316 & a19312;
assign a19320 = ~a19318 & a19250;
assign a19322 = ~a19320 & ~a19244;
assign a19324 = a19318 & ~a19250;
assign a19326 = ~a19324 & ~a19322;
assign a19328 = a17658 & i296;
assign a19330 = ~a17658 & l1058;
assign a19332 = ~a19330 & ~a19328;
assign a19334 = a18572 & l1910;
assign a19336 = a19334 & l880;
assign a19338 = l1914 & ~l1002;
assign a19340 = a19338 & a18586;
assign a19342 = ~a19340 & ~a19336;
assign a19344 = ~l1916 & l890;
assign a19346 = a11208 & ~l890;
assign a19348 = ~a19346 & ~a19344;
assign a19350 = ~a19348 & a18598;
assign a19352 = a19350 & a2746;
assign a19354 = ~a19352 & a19342;
assign a19356 = a18608 & l1918;
assign a19358 = a19356 & l880;
assign a19360 = ~a19358 & a19354;
assign a19362 = l1920 & ~l1006;
assign a19364 = a19362 & a18618;
assign a19366 = ~a19364 & a19360;
assign a19368 = a2530 & l1922;
assign a19370 = a19368 & l880;
assign a19372 = ~a19370 & a19366;
assign a19374 = a18630 & l1924;
assign a19376 = a19374 & a2746;
assign a19378 = ~a19376 & a19372;
assign a19380 = a18638 & l1926;
assign a19382 = a19380 & l880;
assign a19384 = ~a19382 & a19378;
assign a19386 = a18650 & l1928;
assign a19388 = ~a19386 & a19384;
assign a19390 = a18648 & l1930;
assign a19392 = a19390 & l880;
assign a19394 = ~a19392 & a19388;
assign a19396 = ~a19394 & a19332;
assign a19398 = ~a19396 & ~a19326;
assign a19400 = a19394 & ~a19332;
assign a19402 = ~a19400 & ~a19398;
assign a19404 = a17658 & i242;
assign a19406 = ~a17658 & l978;
assign a19408 = ~a19406 & ~a19404;
assign a19410 = ~a19408 & a18838;
assign a19412 = a19408 & ~a18838;
assign a19414 = ~a19412 & ~a19410;
assign a19416 = a19414 & ~a19402;
assign a19418 = a18650 & l1798;
assign a19420 = a18858 & ~l880;
assign a19422 = a18862 & a18664;
assign a19424 = ~a19422 & ~a19420;
assign a19426 = a18874 & a18670;
assign a19428 = ~a19426 & a19424;
assign a19430 = a18880 & ~l880;
assign a19432 = ~a19430 & a19428;
assign a19434 = a18886 & a2526;
assign a19436 = ~a19434 & a19432;
assign a19438 = a18892 & ~l880;
assign a19440 = ~a19438 & a19436;
assign a19442 = a18898 & a18670;
assign a19444 = ~a19442 & a19440;
assign a19446 = a18904 & ~l880;
assign a19448 = ~a19446 & a19444;
assign a19450 = a18696 & l1796;
assign a19452 = ~a19450 & a19448;
assign a19454 = a19452 & ~a19418;
assign a19456 = ~a19454 & a18850;
assign a19458 = a18650 & l1820;
assign a19460 = a18932 & ~l880;
assign a19462 = a18936 & a18664;
assign a19464 = ~a19462 & ~a19460;
assign a19466 = a18948 & a18670;
assign a19468 = ~a19466 & a19464;
assign a19470 = a18954 & ~l880;
assign a19472 = ~a19470 & a19468;
assign a19474 = a18960 & a2526;
assign a19476 = ~a19474 & a19472;
assign a19478 = a18966 & ~l880;
assign a19480 = ~a19478 & a19476;
assign a19482 = a18972 & a18670;
assign a19484 = ~a19482 & a19480;
assign a19486 = a18978 & ~l880;
assign a19488 = ~a19486 & a19484;
assign a19490 = a18696 & l1818;
assign a19492 = ~a19490 & a19488;
assign a19494 = a19492 & ~a19458;
assign a19496 = ~a19494 & a18924;
assign a19498 = ~a19496 & ~a19456;
assign a19500 = a19494 & ~a18924;
assign a19502 = ~a19500 & ~a19498;
assign a19504 = a19068 & ~l880;
assign a19506 = a18696 & l1840;
assign a19508 = a19058 & ~l880;
assign a19510 = a19052 & a18670;
assign a19512 = a19046 & ~l880;
assign a19514 = a19040 & a2526;
assign a19516 = a19034 & ~l880;
assign a19518 = a19028 & a18670;
assign a19520 = a19012 & ~l880;
assign a19522 = a19016 & a18664;
assign a19524 = ~a19522 & ~a19520;
assign a19526 = a19524 & ~a19518;
assign a19528 = a19526 & ~a19516;
assign a19530 = a19528 & ~a19514;
assign a19532 = a19530 & ~a19512;
assign a19534 = a19532 & ~a19510;
assign a19536 = a19534 & ~a19508;
assign a19538 = a19536 & ~a19506;
assign a19540 = a19538 & ~a19504;
assign a19542 = ~a19540 & a19004;
assign a19544 = ~a19542 & ~a19502;
assign a19546 = a19540 & ~a19004;
assign a19548 = ~a19546 & ~a19544;
assign a19550 = a19150 & ~l880;
assign a19552 = a18696 & l1862;
assign a19554 = a19140 & ~l880;
assign a19556 = a19134 & a18670;
assign a19558 = a19128 & ~l880;
assign a19560 = a19122 & a2526;
assign a19562 = a19116 & ~l880;
assign a19564 = a19110 & a18670;
assign a19566 = a19094 & ~l880;
assign a19568 = a19098 & a18664;
assign a19570 = ~a19568 & ~a19566;
assign a19572 = a19570 & ~a19564;
assign a19574 = a19572 & ~a19562;
assign a19576 = a19574 & ~a19560;
assign a19578 = a19576 & ~a19558;
assign a19580 = a19578 & ~a19556;
assign a19582 = a19580 & ~a19554;
assign a19584 = a19582 & ~a19552;
assign a19586 = a19584 & ~a19550;
assign a19588 = ~a19586 & a19086;
assign a19590 = ~a19588 & ~a19548;
assign a19592 = a19586 & ~a19086;
assign a19594 = ~a19592 & ~a19590;
assign a19596 = a19232 & ~l880;
assign a19598 = a18696 & l1884;
assign a19600 = a19222 & ~l880;
assign a19602 = a19216 & a18670;
assign a19604 = a19210 & ~l880;
assign a19606 = a19204 & a2526;
assign a19608 = a19198 & ~l880;
assign a19610 = a19192 & a18670;
assign a19612 = a19176 & ~l880;
assign a19614 = a19180 & a18664;
assign a19616 = ~a19614 & ~a19612;
assign a19618 = a19616 & ~a19610;
assign a19620 = a19618 & ~a19608;
assign a19622 = a19620 & ~a19606;
assign a19624 = a19622 & ~a19604;
assign a19626 = a19624 & ~a19602;
assign a19628 = a19626 & ~a19600;
assign a19630 = a19628 & ~a19598;
assign a19632 = a19630 & ~a19596;
assign a19634 = ~a19632 & a19168;
assign a19636 = ~a19634 & ~a19594;
assign a19638 = a19632 & ~a19168;
assign a19640 = ~a19638 & ~a19636;
assign a19642 = a19314 & ~l880;
assign a19644 = a18696 & l1906;
assign a19646 = a19304 & ~l880;
assign a19648 = a19298 & a18670;
assign a19650 = a19292 & ~l880;
assign a19652 = a19286 & a2526;
assign a19654 = a19280 & ~l880;
assign a19656 = a19274 & a18670;
assign a19658 = a19258 & ~l880;
assign a19660 = a19262 & a18664;
assign a19662 = ~a19660 & ~a19658;
assign a19664 = a19662 & ~a19656;
assign a19666 = a19664 & ~a19654;
assign a19668 = a19666 & ~a19652;
assign a19670 = a19668 & ~a19650;
assign a19672 = a19670 & ~a19648;
assign a19674 = a19672 & ~a19646;
assign a19676 = a19674 & ~a19644;
assign a19678 = a19676 & ~a19642;
assign a19680 = ~a19678 & a19250;
assign a19682 = ~a19680 & ~a19640;
assign a19684 = a19678 & ~a19250;
assign a19686 = ~a19684 & ~a19682;
assign a19688 = a19390 & ~l880;
assign a19690 = a18696 & l1928;
assign a19692 = a19380 & ~l880;
assign a19694 = a19374 & a18670;
assign a19696 = a19368 & ~l880;
assign a19698 = a19362 & a2526;
assign a19700 = a19356 & ~l880;
assign a19702 = a19350 & a18670;
assign a19704 = a19334 & ~l880;
assign a19706 = a19338 & a18664;
assign a19708 = ~a19706 & ~a19704;
assign a19710 = a19708 & ~a19702;
assign a19712 = a19710 & ~a19700;
assign a19714 = a19712 & ~a19698;
assign a19716 = a19714 & ~a19696;
assign a19718 = a19716 & ~a19694;
assign a19720 = a19718 & ~a19692;
assign a19722 = a19720 & ~a19690;
assign a19724 = a19722 & ~a19688;
assign a19726 = ~a19724 & a19332;
assign a19728 = ~a19726 & ~a19686;
assign a19730 = a19724 & ~a19332;
assign a19732 = ~a19730 & ~a19728;
assign a19734 = ~a19408 & a18798;
assign a19736 = a19408 & ~a18798;
assign a19738 = ~a19736 & ~a19734;
assign a19740 = a19738 & a19732;
assign a19742 = ~a19740 & ~a19416;
assign a19744 = ~a19742 & ~a18844;
assign a19746 = a19416 & a18844;
assign a19748 = a19746 & a19732;
assign a19750 = ~a19748 & ~a19744;
assign a19752 = a19750 & a18744;
assign a19754 = ~a19752 & a18738;
assign a19758 = a2768 & l1960;
assign a19760 = l1964 & l1244;
assign a19762 = a19760 & a19758;
assign a19764 = ~l1968 & ~l1960;
assign a19766 = ~l1964 & ~l1956;
assign a19768 = a19766 & l1244;
assign a19770 = a19768 & a19764;
assign a19772 = ~a19770 & ~a19762;
assign a19774 = a19758 & ~l1968;
assign a19776 = a19774 & ~l1156;
assign a19778 = ~a2740 & l1956;
assign a19780 = a19778 & a19776;
assign a19782 = l1968 & l1156;
assign a19784 = a19782 & a19758;
assign a19786 = a19784 & a2740;
assign a19788 = a19786 & ~l1956;
assign a19790 = l1968 & l1956;
assign a19792 = a2740 & l1156;
assign a19794 = a19792 & a19790;
assign a19796 = a19784 & a19778;
assign a19798 = ~a19796 & ~a19794;
assign a19800 = a19798 & ~a19788;
assign a19802 = a19800 & ~a19780;
assign a19804 = l1968 & ~l1156;
assign a19806 = a19804 & ~a2740;
assign a19808 = ~a19806 & a19802;
assign a19810 = a19808 & a19772;
assign a19812 = l1964 & l1156;
assign a19814 = ~a2740 & l1964;
assign a19816 = l1964 & ~l1244;
assign a19818 = a19816 & ~a2768;
assign a19820 = ~l1960 & ~l1956;
assign a19822 = a19820 & ~l1156;
assign a19824 = a19822 & ~a2740;
assign a19826 = a19764 & l1156;
assign a19828 = a19826 & ~l1956;
assign a19830 = a19804 & ~l1244;
assign a19832 = a19830 & ~a2768;
assign a19834 = a2740 & l1956;
assign a19836 = a19834 & ~l1156;
assign a19838 = a19836 & ~l1244;
assign a19840 = a19838 & ~a2768;
assign a19842 = ~a2768 & ~l1244;
assign a19844 = a19842 & a19822;
assign a19846 = ~a19844 & ~a19840;
assign a19848 = a19846 & ~a19832;
assign a19850 = a19848 & ~a19828;
assign a19852 = a19850 & ~a19824;
assign a19854 = a19852 & ~a19818;
assign a19856 = a19854 & ~a19814;
assign a19858 = a19856 & ~a19812;
assign a19860 = a19858 & a19810;
assign a19862 = ~a19860 & l924;
assign a19864 = ~l1164 & ~l1162;
assign a19866 = l1150 & l1148;
assign a19868 = a19866 & ~l1166;
assign a19870 = a19868 & a19864;
assign a19872 = ~l1526 & l890;
assign a19874 = ~l890 & ~i92;
assign a19876 = ~a19874 & ~a19872;
assign a19878 = a19876 & ~a2768;
assign a19880 = a19878 & ~l1244;
assign a19882 = a19880 & ~l1156;
assign a19884 = a19882 & a2740;
assign a19886 = ~a19884 & ~a18568;
assign a19888 = ~a19886 & ~l886;
assign a19890 = a19888 & ~a19870;
assign a19896 = ~l936 & l890;
assign a19898 = ~a5366 & ~l890;
assign a19902 = ~a5408 & l1058;
assign a19904 = l1144 & l1100;
assign a19906 = ~a17686 & ~a17112;
assign a19908 = ~a14378 & l1142;
assign a19910 = ~a19908 & ~a14514;
assign a19912 = ~a19910 & a17686;
assign a19914 = ~a19912 & ~a19906;
assign a19916 = ~a19914 & ~l1100;
assign a19918 = ~a19916 & ~a19904;
assign a19920 = ~a19918 & a5408;
assign a19922 = ~a19920 & ~a19902;
assign a19924 = a19922 & ~a14090;
assign a19926 = ~a19922 & a14090;
assign a19928 = ~a19926 & ~a19924;
assign a19930 = ~a5408 & l1054;
assign a19932 = l1136 & l1100;
assign a19934 = ~a17686 & ~a17016;
assign a19936 = ~a14378 & l1134;
assign a19938 = ~a19936 & ~a14494;
assign a19940 = ~a19938 & a17686;
assign a19942 = ~a19940 & ~a19934;
assign a19944 = ~a19942 & ~l1100;
assign a19946 = ~a19944 & ~a19932;
assign a19948 = ~a19946 & a5408;
assign a19950 = ~a19948 & ~a19930;
assign a19952 = a19950 & ~a13932;
assign a19954 = ~a19950 & a13932;
assign a19956 = ~a6286 & ~a5408;
assign a19958 = ~a16906 & l1100;
assign a19960 = ~a17686 & ~a16920;
assign a19962 = ~a14378 & ~a14298;
assign a19964 = ~a19962 & ~a14474;
assign a19966 = ~a19964 & a17686;
assign a19968 = ~a19966 & ~a19960;
assign a19970 = ~a19968 & ~l1100;
assign a19972 = ~a19970 & ~a19958;
assign a19974 = ~a19972 & a5408;
assign a19978 = a19976 & ~a13754;
assign a19980 = ~a19976 & a13754;
assign a19982 = ~a6278 & ~a5408;
assign a19984 = ~a16802 & l1100;
assign a19986 = ~a17686 & ~a16816;
assign a19988 = ~a14378 & ~a14312;
assign a19990 = ~a19988 & ~a14454;
assign a19992 = ~a19990 & a17686;
assign a19994 = ~a19992 & ~a19986;
assign a19996 = ~a19994 & ~l1100;
assign a19998 = ~a19996 & ~a19984;
assign a20000 = ~a19998 & a5408;
assign a20004 = a20002 & ~a13564;
assign a20006 = ~a20002 & a13564;
assign a20008 = ~a6270 & ~a5408;
assign a20010 = ~a16698 & l1100;
assign a20012 = ~a17686 & ~a16712;
assign a20014 = ~a14378 & ~a14326;
assign a20016 = ~a20014 & ~a14434;
assign a20018 = ~a20016 & a17686;
assign a20020 = ~a20018 & ~a20012;
assign a20022 = ~a20020 & ~l1100;
assign a20024 = ~a20022 & ~a20010;
assign a20026 = ~a20024 & a5408;
assign a20030 = a20028 & ~a13374;
assign a20032 = ~a20028 & a13374;
assign a20034 = ~a6262 & ~a5408;
assign a20036 = ~a16594 & l1100;
assign a20038 = ~a17686 & ~a16608;
assign a20040 = ~a14378 & ~a14340;
assign a20042 = ~a20040 & ~a14414;
assign a20044 = ~a20042 & a17686;
assign a20046 = ~a20044 & ~a20038;
assign a20048 = ~a20046 & ~l1100;
assign a20050 = ~a20048 & ~a20036;
assign a20052 = ~a20050 & a5408;
assign a20056 = a20054 & ~a13184;
assign a20058 = ~a6254 & ~a5408;
assign a20060 = ~a16236 & l1100;
assign a20062 = ~a17686 & ~a16250;
assign a20064 = ~a14378 & ~a14354;
assign a20066 = ~a20064 & ~a14400;
assign a20068 = ~a20066 & a17686;
assign a20070 = ~a20068 & ~a20062;
assign a20072 = ~a20070 & ~l1100;
assign a20074 = ~a20072 & ~a20060;
assign a20076 = ~a20074 & a5408;
assign a20080 = ~a20078 & a13000;
assign a20082 = ~a20054 & a13184;
assign a20084 = ~a20082 & ~a20080;
assign a20086 = ~a20084 & ~a20056;
assign a20088 = ~a20086 & ~a20032;
assign a20090 = ~a20088 & ~a20030;
assign a20092 = ~a20090 & ~a20006;
assign a20094 = ~a20092 & ~a20004;
assign a20096 = ~a20094 & ~a19980;
assign a20098 = ~a20096 & ~a19978;
assign a20100 = ~a20098 & ~a19954;
assign a20102 = ~a20100 & ~a19952;
assign a20104 = ~a20102 & ~a19928;
assign a20106 = a20102 & a19928;
assign a20108 = ~a20106 & ~a20104;
assign a20110 = ~a19954 & ~a19952;
assign a20112 = ~a20110 & ~a20098;
assign a20114 = a20110 & a20098;
assign a20116 = ~a20114 & ~a20112;
assign a20118 = ~a19980 & ~a19978;
assign a20120 = ~a20118 & ~a20094;
assign a20122 = a20118 & a20094;
assign a20124 = ~a20122 & ~a20120;
assign a20126 = ~a20006 & ~a20004;
assign a20128 = ~a20126 & ~a20090;
assign a20130 = a20126 & a20090;
assign a20132 = ~a20130 & ~a20128;
assign a20134 = ~a20032 & ~a20030;
assign a20136 = ~a20134 & ~a20086;
assign a20138 = a20134 & a20086;
assign a20140 = ~a20138 & ~a20136;
assign a20142 = ~a20082 & ~a20056;
assign a20144 = ~a20142 & ~a20080;
assign a20146 = a20142 & a20080;
assign a20148 = ~a20146 & ~a20144;
assign a20150 = a20078 & ~a13000;
assign a20152 = ~a20150 & ~a20080;
assign a20154 = ~a5408 & l978;
assign a20156 = l1100 & l996;
assign a20158 = ~a17686 & ~a16278;
assign a20160 = ~a14378 & l994;
assign a20162 = ~a20160 & ~a14382;
assign a20164 = ~a20162 & a17686;
assign a20166 = ~a20164 & ~a20158;
assign a20168 = ~a20166 & ~l1100;
assign a20170 = ~a20168 & ~a20156;
assign a20172 = ~a20170 & a5408;
assign a20174 = ~a20172 & ~a20154;
assign a20176 = a20174 & ~a12726;
assign a20178 = ~a20174 & a12726;
assign a20180 = ~a20178 & ~a20176;
assign a20182 = ~a20180 & a20152;
assign a20184 = a20182 & a20142;
assign a20186 = a20184 & a20134;
assign a20188 = a20186 & a20126;
assign a20190 = a20188 & a20118;
assign a20192 = a20190 & a20110;
assign a20194 = a20192 & a19928;
assign a20196 = ~a20194 & a20152;
assign a20198 = a20196 & a20148;
assign a20200 = a20198 & a20140;
assign a20202 = a20200 & a20132;
assign a20204 = a20202 & a20124;
assign a20206 = a20204 & a20116;
assign a20208 = a20206 & a20108;
assign a20210 = ~i522 & ~i520;
assign a20212 = ~a20210 & i524;
assign a20214 = a20212 & i518;
assign a20216 = a20214 & i516;
assign a20218 = a20216 & i514;
assign a20220 = a20218 & i512;
assign a20222 = i526 & i510;
assign a20224 = a20222 & i528;
assign a20226 = a20224 & i530;
assign a20228 = a20226 & i522;
assign a20230 = a20228 & i520;
assign a20232 = ~a20230 & i524;
assign a20234 = a20230 & ~i524;
assign a20236 = ~a20234 & ~a20232;
assign a20238 = a20236 & ~a20220;
assign a20240 = ~a20152 & a20108;
assign a20242 = a20240 & a20116;
assign a20244 = a20238 & ~a20152;
assign a20246 = a20230 & i524;
assign a20248 = ~a20246 & i518;
assign a20250 = a20246 & ~i518;
assign a20252 = ~a20250 & ~a20248;
assign a20254 = a20252 & ~a20220;
assign a20256 = a20242 & a20124;
assign a20258 = a20254 & ~a20152;
assign a20260 = a20246 & i518;
assign a20262 = ~a20260 & i516;
assign a20264 = a20260 & ~i516;
assign a20266 = ~a20264 & ~a20262;
assign a20268 = a20266 & ~a20220;
assign a20270 = a20256 & a20132;
assign a20272 = a20268 & ~a20152;
assign a20274 = a20260 & i516;
assign a20276 = ~a20274 & i514;
assign a20278 = a20274 & ~i514;
assign a20280 = ~a20278 & ~a20276;
assign a20282 = a20280 & ~a20220;
assign a20284 = a20270 & a20140;
assign a20286 = a20282 & ~a20152;
assign a20288 = a20274 & i514;
assign a20290 = ~a20288 & i512;
assign a20292 = a20288 & ~i512;
assign a20294 = ~a20292 & ~a20290;
assign a20296 = a20294 & ~a20220;
assign a20298 = a20296 & ~a20152;
assign a20300 = ~a20298 & a20284;
assign a20302 = a20300 & a20148;
assign a20304 = ~a20302 & ~a20296;
assign a20306 = ~a20304 & ~a20148;
assign a20308 = ~a20306 & ~a20286;
assign a20310 = a20304 & a20148;
assign a20312 = ~a20310 & ~a20308;
assign a20314 = ~a20312 & a20284;
assign a20316 = ~a20314 & ~a20282;
assign a20318 = ~a20316 & ~a20148;
assign a20320 = ~a20318 & ~a20272;
assign a20322 = a20316 & a20148;
assign a20324 = ~a20322 & ~a20320;
assign a20326 = ~a20148 & a20108;
assign a20328 = a20326 & a20116;
assign a20330 = a20328 & a20124;
assign a20332 = a20330 & a20132;
assign a20334 = a20332 & ~a20312;
assign a20336 = a20334 & a20140;
assign a20338 = ~a20336 & a20304;
assign a20340 = ~a20338 & ~a20140;
assign a20342 = ~a20340 & ~a20324;
assign a20344 = a20338 & a20140;
assign a20346 = ~a20344 & ~a20342;
assign a20348 = ~a20346 & a20270;
assign a20350 = ~a20348 & ~a20268;
assign a20352 = a20348 & a20268;
assign a20354 = ~a20352 & ~a20350;
assign a20356 = a20354 & ~a20148;
assign a20358 = ~a20356 & ~a20258;
assign a20360 = ~a20354 & a20148;
assign a20362 = ~a20360 & ~a20358;
assign a20364 = ~a20346 & a20332;
assign a20366 = ~a20364 & a20316;
assign a20368 = a20364 & ~a20316;
assign a20370 = ~a20368 & ~a20366;
assign a20372 = ~a20370 & ~a20352;
assign a20374 = ~a20372 & ~a20140;
assign a20376 = ~a20374 & ~a20362;
assign a20378 = a20372 & a20140;
assign a20380 = ~a20378 & ~a20376;
assign a20382 = ~a20140 & a20108;
assign a20384 = a20382 & a20116;
assign a20386 = a20384 & a20124;
assign a20388 = a20386 & ~a20346;
assign a20390 = a20388 & a20132;
assign a20392 = ~a20390 & ~a20368;
assign a20394 = a20392 & a20338;
assign a20396 = ~a20394 & ~a20132;
assign a20398 = ~a20396 & ~a20380;
assign a20400 = a20394 & a20132;
assign a20402 = ~a20400 & ~a20398;
assign a20404 = ~a20402 & a20256;
assign a20406 = ~a20404 & ~a20254;
assign a20408 = a20404 & a20254;
assign a20410 = ~a20408 & ~a20406;
assign a20412 = a20410 & ~a20148;
assign a20414 = ~a20412 & ~a20244;
assign a20416 = ~a20410 & a20148;
assign a20418 = ~a20416 & ~a20414;
assign a20420 = ~a20402 & a20330;
assign a20422 = ~a20420 & ~a20354;
assign a20424 = a20420 & a20354;
assign a20426 = ~a20424 & ~a20422;
assign a20428 = ~a20426 & ~a20408;
assign a20430 = a20426 & a20408;
assign a20432 = ~a20430 & ~a20428;
assign a20434 = a20432 & ~a20140;
assign a20436 = ~a20434 & ~a20418;
assign a20438 = ~a20432 & a20140;
assign a20440 = ~a20438 & ~a20436;
assign a20442 = ~a20402 & a20386;
assign a20444 = ~a20442 & a20372;
assign a20446 = a20442 & ~a20372;
assign a20448 = ~a20446 & ~a20444;
assign a20450 = ~a20424 & ~a20408;
assign a20452 = ~a20450 & ~a20422;
assign a20454 = ~a20452 & ~a20448;
assign a20456 = a20452 & a20448;
assign a20458 = ~a20456 & ~a20454;
assign a20460 = a20458 & ~a20132;
assign a20462 = ~a20460 & ~a20440;
assign a20464 = ~a20458 & a20132;
assign a20466 = ~a20464 & ~a20462;
assign a20468 = ~a20132 & a20108;
assign a20470 = a20468 & a20116;
assign a20472 = a20470 & ~a20402;
assign a20474 = a20472 & a20124;
assign a20476 = ~a20452 & ~a20446;
assign a20478 = ~a20476 & ~a20444;
assign a20480 = ~a20478 & ~a20474;
assign a20482 = a20480 & a20394;
assign a20484 = ~a20482 & ~a20124;
assign a20486 = ~a20484 & ~a20466;
assign a20488 = a20482 & a20124;
assign a20490 = ~a20488 & ~a20486;
assign a20492 = ~a20490 & a20242;
assign a20494 = a20492 & a20238;
assign a20496 = ~a20490 & a20328;
assign a20498 = ~a20496 & ~a20410;
assign a20500 = a20496 & a20410;
assign a20502 = ~a20500 & ~a20498;
assign a20504 = ~a20502 & ~a20494;
assign a20506 = a20502 & a20494;
assign a20508 = ~a20506 & ~a20504;
assign a20510 = ~a20228 & i520;
assign a20512 = a20228 & ~i520;
assign a20514 = ~a20512 & ~a20510;
assign a20516 = ~a20514 & ~a20220;
assign a20518 = ~a20516 & ~a20152;
assign a20520 = ~a20492 & ~a20238;
assign a20522 = ~a20520 & ~a20494;
assign a20524 = a20522 & ~a20148;
assign a20526 = ~a20524 & ~a20518;
assign a20528 = ~a20522 & a20148;
assign a20530 = ~a20528 & ~a20526;
assign a20532 = a20508 & ~a20140;
assign a20534 = ~a20532 & ~a20530;
assign a20536 = ~a20508 & a20140;
assign a20538 = ~a20536 & ~a20534;
assign a20540 = ~a20490 & a20384;
assign a20542 = ~a20540 & ~a20432;
assign a20544 = a20540 & a20432;
assign a20546 = ~a20544 & ~a20542;
assign a20548 = ~a20500 & ~a20494;
assign a20550 = ~a20548 & ~a20498;
assign a20552 = ~a20550 & ~a20546;
assign a20554 = a20550 & a20546;
assign a20556 = ~a20554 & ~a20552;
assign a20558 = a20556 & ~a20132;
assign a20560 = ~a20558 & ~a20538;
assign a20562 = ~a20556 & a20132;
assign a20564 = ~a20562 & ~a20560;
assign a20566 = ~a20490 & a20470;
assign a20568 = ~a20566 & ~a20458;
assign a20570 = a20566 & a20458;
assign a20572 = ~a20570 & ~a20568;
assign a20574 = ~a20550 & ~a20544;
assign a20576 = ~a20574 & ~a20542;
assign a20578 = ~a20576 & ~a20572;
assign a20580 = a20576 & a20572;
assign a20582 = ~a20580 & ~a20578;
assign a20584 = a20582 & ~a20124;
assign a20586 = ~a20584 & ~a20564;
assign a20588 = ~a20582 & a20124;
assign a20590 = ~a20588 & ~a20586;
assign a20592 = ~a20124 & a20108;
assign a20594 = a20592 & ~a20490;
assign a20596 = a20594 & a20116;
assign a20598 = ~a20576 & ~a20570;
assign a20600 = ~a20598 & ~a20568;
assign a20602 = ~a20600 & ~a20596;
assign a20604 = a20602 & a20482;
assign a20606 = ~a20604 & ~a20116;
assign a20608 = ~a20606 & ~a20590;
assign a20610 = a20604 & a20116;
assign a20612 = ~a20610 & ~a20608;
assign a20614 = ~a20612 & a20382;
assign a20616 = ~a20614 & ~a20508;
assign a20618 = a20614 & a20508;
assign a20620 = ~a20618 & ~a20616;
assign a20622 = ~a20612 & a20326;
assign a20624 = ~a20622 & ~a20522;
assign a20626 = ~a20612 & a20240;
assign a20628 = a20626 & ~a20516;
assign a20630 = a20622 & a20522;
assign a20632 = ~a20630 & ~a20628;
assign a20634 = ~a20632 & ~a20624;
assign a20636 = ~a20634 & ~a20620;
assign a20638 = a20634 & a20620;
assign a20640 = ~a20638 & ~a20636;
assign a20642 = ~a20226 & i522;
assign a20644 = a20226 & ~i522;
assign a20646 = ~a20644 & ~a20642;
assign a20648 = a20646 & ~a20220;
assign a20650 = a20648 & ~a20152;
assign a20652 = ~a20626 & a20516;
assign a20654 = ~a20652 & ~a20628;
assign a20656 = a20654 & ~a20148;
assign a20658 = ~a20656 & ~a20650;
assign a20660 = ~a20654 & a20148;
assign a20662 = ~a20660 & ~a20658;
assign a20664 = ~a20630 & ~a20624;
assign a20666 = ~a20664 & ~a20628;
assign a20668 = a20664 & a20628;
assign a20670 = ~a20668 & ~a20666;
assign a20672 = a20670 & ~a20140;
assign a20674 = ~a20672 & ~a20662;
assign a20676 = ~a20670 & a20140;
assign a20678 = ~a20676 & ~a20674;
assign a20680 = a20640 & ~a20132;
assign a20682 = ~a20680 & ~a20678;
assign a20684 = ~a20640 & a20132;
assign a20686 = ~a20684 & ~a20682;
assign a20688 = ~a20612 & a20468;
assign a20690 = ~a20688 & ~a20556;
assign a20692 = a20688 & a20556;
assign a20694 = ~a20692 & ~a20690;
assign a20696 = ~a20634 & ~a20618;
assign a20698 = ~a20696 & ~a20616;
assign a20700 = ~a20698 & ~a20694;
assign a20702 = a20698 & a20694;
assign a20704 = ~a20702 & ~a20700;
assign a20706 = a20704 & ~a20124;
assign a20708 = ~a20706 & ~a20686;
assign a20710 = ~a20704 & a20124;
assign a20712 = ~a20710 & ~a20708;
assign a20714 = ~a20612 & a20592;
assign a20716 = ~a20714 & ~a20582;
assign a20718 = a20714 & a20582;
assign a20720 = ~a20718 & ~a20716;
assign a20722 = ~a20698 & ~a20692;
assign a20724 = ~a20722 & ~a20690;
assign a20726 = ~a20724 & ~a20720;
assign a20728 = a20724 & a20720;
assign a20730 = ~a20728 & ~a20726;
assign a20732 = a20730 & ~a20116;
assign a20734 = ~a20732 & ~a20712;
assign a20736 = ~a20730 & a20116;
assign a20738 = ~a20736 & ~a20734;
assign a20740 = ~a20612 & ~a20116;
assign a20742 = a20740 & a20108;
assign a20744 = ~a20724 & ~a20718;
assign a20746 = ~a20744 & ~a20716;
assign a20748 = ~a20746 & ~a20742;
assign a20750 = a20748 & a20604;
assign a20752 = ~a20750 & ~a20108;
assign a20754 = ~a20752 & ~a20738;
assign a20756 = a20750 & a20108;
assign a20758 = ~a20756 & ~a20754;
assign a20760 = ~a20758 & ~a20132;
assign a20762 = ~a20760 & ~a20640;
assign a20764 = a20760 & a20640;
assign a20766 = ~a20764 & ~a20762;
assign a20768 = ~a20758 & ~a20140;
assign a20770 = ~a20768 & ~a20670;
assign a20772 = a20768 & a20670;
assign a20774 = ~a20758 & ~a20148;
assign a20776 = ~a20774 & ~a20654;
assign a20778 = ~a20758 & ~a20152;
assign a20780 = a20778 & a20648;
assign a20782 = a20774 & a20654;
assign a20784 = ~a20782 & ~a20780;
assign a20786 = ~a20784 & ~a20776;
assign a20788 = ~a20786 & ~a20772;
assign a20790 = ~a20788 & ~a20770;
assign a20792 = ~a20790 & ~a20766;
assign a20794 = a20790 & a20766;
assign a20796 = ~a20794 & ~a20792;
assign a20798 = ~a20224 & i530;
assign a20800 = a20224 & ~i530;
assign a20802 = ~a20800 & ~a20798;
assign a20804 = ~a20802 & ~a20220;
assign a20806 = ~a20804 & ~a20152;
assign a20808 = ~a20778 & ~a20648;
assign a20810 = ~a20808 & ~a20780;
assign a20812 = a20810 & ~a20148;
assign a20814 = ~a20812 & ~a20806;
assign a20816 = ~a20810 & a20148;
assign a20818 = ~a20816 & ~a20814;
assign a20820 = ~a20782 & ~a20776;
assign a20822 = ~a20820 & ~a20780;
assign a20824 = a20820 & a20780;
assign a20826 = ~a20824 & ~a20822;
assign a20828 = a20826 & ~a20140;
assign a20830 = ~a20828 & ~a20818;
assign a20832 = ~a20826 & a20140;
assign a20834 = ~a20832 & ~a20830;
assign a20836 = ~a20772 & ~a20770;
assign a20838 = ~a20836 & ~a20786;
assign a20840 = a20836 & a20786;
assign a20842 = ~a20840 & ~a20838;
assign a20844 = a20842 & ~a20132;
assign a20846 = ~a20844 & ~a20834;
assign a20848 = ~a20842 & a20132;
assign a20850 = ~a20848 & ~a20846;
assign a20852 = a20796 & ~a20124;
assign a20854 = ~a20852 & ~a20850;
assign a20856 = ~a20796 & a20124;
assign a20858 = ~a20856 & ~a20854;
assign a20860 = ~a20758 & ~a20124;
assign a20862 = ~a20860 & ~a20704;
assign a20864 = a20860 & a20704;
assign a20866 = ~a20864 & ~a20862;
assign a20868 = ~a20790 & ~a20764;
assign a20870 = ~a20868 & ~a20762;
assign a20872 = ~a20870 & ~a20866;
assign a20874 = a20870 & a20866;
assign a20876 = ~a20874 & ~a20872;
assign a20878 = a20876 & ~a20116;
assign a20880 = ~a20878 & ~a20858;
assign a20882 = ~a20876 & a20116;
assign a20884 = ~a20882 & ~a20880;
assign a20886 = ~a20758 & ~a20116;
assign a20888 = ~a20886 & ~a20730;
assign a20890 = a20886 & a20730;
assign a20892 = ~a20890 & ~a20888;
assign a20894 = ~a20870 & ~a20864;
assign a20896 = ~a20894 & ~a20862;
assign a20898 = ~a20896 & ~a20892;
assign a20900 = a20896 & a20892;
assign a20902 = ~a20900 & ~a20898;
assign a20904 = a20902 & ~a20108;
assign a20906 = ~a20904 & ~a20884;
assign a20908 = ~a20902 & a20108;
assign a20910 = ~a20908 & ~a20906;
assign a20912 = ~a20758 & ~a20108;
assign a20914 = ~a20896 & ~a20890;
assign a20916 = ~a20914 & ~a20888;
assign a20918 = ~a20916 & ~a20912;
assign a20920 = a20918 & a20750;
assign a20922 = ~a20920 & a20194;
assign a20924 = ~a20922 & ~a20910;
assign a20926 = a20920 & ~a20194;
assign a20928 = ~a20926 & ~a20924;
assign a20930 = ~a20928 & ~a20124;
assign a20932 = ~a20930 & ~a20796;
assign a20934 = a20930 & a20796;
assign a20936 = ~a20934 & ~a20932;
assign a20938 = ~a20928 & ~a20132;
assign a20940 = ~a20938 & ~a20842;
assign a20942 = a20938 & a20842;
assign a20944 = ~a20928 & ~a20140;
assign a20946 = ~a20944 & ~a20826;
assign a20948 = a20944 & a20826;
assign a20950 = ~a20928 & ~a20148;
assign a20952 = ~a20950 & ~a20810;
assign a20954 = ~a20928 & ~a20152;
assign a20956 = a20954 & ~a20804;
assign a20958 = a20950 & a20810;
assign a20960 = ~a20958 & ~a20956;
assign a20962 = ~a20960 & ~a20952;
assign a20964 = ~a20962 & ~a20948;
assign a20966 = ~a20964 & ~a20946;
assign a20968 = ~a20966 & ~a20942;
assign a20970 = ~a20968 & ~a20940;
assign a20972 = ~a20970 & ~a20936;
assign a20974 = a20970 & a20936;
assign a20976 = ~a20974 & ~a20972;
assign a20978 = ~a20222 & i528;
assign a20980 = a20222 & ~i528;
assign a20982 = ~a20980 & ~a20978;
assign a20984 = ~a20982 & ~a20220;
assign a20986 = ~a20984 & ~a20152;
assign a20988 = ~a20954 & a20804;
assign a20990 = ~a20988 & ~a20956;
assign a20992 = a20990 & ~a20148;
assign a20994 = ~a20992 & ~a20986;
assign a20996 = ~a20990 & a20148;
assign a20998 = ~a20996 & ~a20994;
assign a21000 = ~a20958 & ~a20952;
assign a21002 = ~a21000 & ~a20956;
assign a21004 = a21000 & a20956;
assign a21006 = ~a21004 & ~a21002;
assign a21008 = a21006 & ~a20140;
assign a21010 = ~a21008 & ~a20998;
assign a21012 = ~a21006 & a20140;
assign a21014 = ~a21012 & ~a21010;
assign a21016 = ~a20948 & ~a20946;
assign a21018 = ~a21016 & ~a20962;
assign a21020 = a21016 & a20962;
assign a21022 = ~a21020 & ~a21018;
assign a21024 = a21022 & ~a20132;
assign a21026 = ~a21024 & ~a21014;
assign a21028 = ~a21022 & a20132;
assign a21030 = ~a21028 & ~a21026;
assign a21032 = ~a20942 & ~a20940;
assign a21034 = ~a21032 & ~a20966;
assign a21036 = a21032 & a20966;
assign a21038 = ~a21036 & ~a21034;
assign a21040 = a21038 & ~a20124;
assign a21042 = ~a21040 & ~a21030;
assign a21044 = ~a21038 & a20124;
assign a21046 = ~a21044 & ~a21042;
assign a21048 = a20976 & ~a20116;
assign a21050 = ~a21048 & ~a21046;
assign a21052 = ~a20976 & a20116;
assign a21054 = ~a21052 & ~a21050;
assign a21056 = ~a20928 & ~a20116;
assign a21058 = ~a21056 & ~a20876;
assign a21060 = a21056 & a20876;
assign a21062 = ~a21060 & ~a21058;
assign a21064 = ~a20970 & ~a20934;
assign a21066 = ~a21064 & ~a20932;
assign a21068 = ~a21066 & ~a21062;
assign a21070 = a21066 & a21062;
assign a21072 = ~a21070 & ~a21068;
assign a21074 = a21072 & ~a20108;
assign a21076 = ~a21074 & ~a21054;
assign a21078 = ~a21072 & a20108;
assign a21080 = ~a21078 & ~a21076;
assign a21082 = ~a20928 & ~a20108;
assign a21084 = ~a21082 & ~a20902;
assign a21086 = a21082 & a20902;
assign a21088 = ~a21086 & ~a21084;
assign a21090 = ~a21066 & ~a21060;
assign a21092 = ~a21090 & ~a21058;
assign a21094 = ~a21092 & ~a21088;
assign a21096 = a21092 & a21088;
assign a21098 = ~a21096 & ~a21094;
assign a21100 = a21098 & a20194;
assign a21102 = ~a21100 & ~a21080;
assign a21104 = ~a21098 & ~a20194;
assign a21106 = ~a21104 & ~a21102;
assign a21108 = ~a21106 & ~a20116;
assign a21110 = ~a21108 & ~a20976;
assign a21112 = a21108 & a20976;
assign a21114 = ~a21112 & ~a21110;
assign a21116 = ~a21106 & ~a20124;
assign a21118 = ~a21116 & ~a21038;
assign a21120 = a21116 & a21038;
assign a21122 = ~a21106 & ~a20132;
assign a21124 = ~a21122 & ~a21022;
assign a21126 = a21122 & a21022;
assign a21128 = ~a21106 & ~a20140;
assign a21130 = ~a21128 & ~a21006;
assign a21132 = a21128 & a21006;
assign a21134 = ~a21106 & ~a20148;
assign a21136 = ~a21134 & ~a20990;
assign a21138 = ~a21106 & ~a20152;
assign a21140 = a21138 & ~a20984;
assign a21142 = a21134 & a20990;
assign a21144 = ~a21142 & ~a21140;
assign a21146 = ~a21144 & ~a21136;
assign a21148 = ~a21146 & ~a21132;
assign a21150 = ~a21148 & ~a21130;
assign a21152 = ~a21150 & ~a21126;
assign a21154 = ~a21152 & ~a21124;
assign a21156 = ~a21154 & ~a21120;
assign a21158 = ~a21156 & ~a21118;
assign a21160 = ~a21158 & ~a21114;
assign a21162 = a21158 & a21114;
assign a21164 = ~a21162 & ~a21160;
assign a21166 = i526 & ~i510;
assign a21168 = ~i526 & i510;
assign a21170 = ~a21168 & ~a21166;
assign a21172 = ~a21170 & ~a20220;
assign a21174 = ~a21172 & ~a20152;
assign a21176 = ~a21138 & a20984;
assign a21178 = ~a21176 & ~a21140;
assign a21180 = a21178 & ~a20148;
assign a21182 = ~a21180 & ~a21174;
assign a21184 = ~a21178 & a20148;
assign a21186 = ~a21184 & ~a21182;
assign a21188 = ~a21142 & ~a21136;
assign a21190 = ~a21188 & ~a21140;
assign a21192 = a21188 & a21140;
assign a21194 = ~a21192 & ~a21190;
assign a21196 = a21194 & ~a20140;
assign a21198 = ~a21196 & ~a21186;
assign a21200 = ~a21194 & a20140;
assign a21202 = ~a21200 & ~a21198;
assign a21204 = ~a21132 & ~a21130;
assign a21206 = ~a21204 & ~a21146;
assign a21208 = a21204 & a21146;
assign a21210 = ~a21208 & ~a21206;
assign a21212 = a21210 & ~a20132;
assign a21214 = ~a21212 & ~a21202;
assign a21216 = ~a21210 & a20132;
assign a21218 = ~a21216 & ~a21214;
assign a21220 = ~a21126 & ~a21124;
assign a21222 = ~a21220 & ~a21150;
assign a21224 = a21220 & a21150;
assign a21226 = ~a21224 & ~a21222;
assign a21228 = a21226 & ~a20124;
assign a21230 = ~a21228 & ~a21218;
assign a21232 = ~a21226 & a20124;
assign a21234 = ~a21232 & ~a21230;
assign a21236 = ~a21120 & ~a21118;
assign a21238 = ~a21236 & ~a21154;
assign a21240 = a21236 & a21154;
assign a21242 = ~a21240 & ~a21238;
assign a21244 = a21242 & ~a20116;
assign a21246 = ~a21244 & ~a21234;
assign a21248 = ~a21242 & a20116;
assign a21250 = ~a21248 & ~a21246;
assign a21252 = a21164 & ~a20108;
assign a21254 = ~a21252 & ~a21250;
assign a21256 = ~a21164 & a20108;
assign a21258 = ~a21256 & ~a21254;
assign a21260 = ~a21106 & ~a20108;
assign a21262 = ~a21260 & ~a21072;
assign a21264 = a21260 & a21072;
assign a21266 = ~a21264 & ~a21262;
assign a21268 = ~a21158 & ~a21112;
assign a21270 = ~a21268 & ~a21110;
assign a21272 = ~a21270 & ~a21266;
assign a21274 = a21270 & a21266;
assign a21276 = ~a21274 & ~a21272;
assign a21278 = a21276 & a20194;
assign a21280 = ~a21278 & ~a21258;
assign a21282 = ~a21276 & ~a20194;
assign a21284 = ~a21282 & ~a21280;
assign a21286 = ~a21284 & ~a20108;
assign a21288 = ~a21286 & ~a21164;
assign a21290 = a21286 & a21164;
assign a21292 = ~a21290 & ~a21288;
assign a21294 = ~a21284 & ~a20116;
assign a21296 = ~a21294 & ~a21242;
assign a21298 = a21294 & a21242;
assign a21300 = ~a21284 & ~a20124;
assign a21302 = ~a21300 & ~a21226;
assign a21304 = a21300 & a21226;
assign a21306 = ~a21284 & ~a20132;
assign a21308 = ~a21306 & ~a21210;
assign a21310 = a21306 & a21210;
assign a21312 = ~a21284 & ~a20140;
assign a21314 = ~a21312 & ~a21194;
assign a21316 = a21312 & a21194;
assign a21318 = ~a21284 & ~a20148;
assign a21320 = ~a21318 & ~a21178;
assign a21322 = ~a21284 & ~a20152;
assign a21324 = a21322 & ~a21172;
assign a21326 = a21318 & a21178;
assign a21328 = ~a21326 & ~a21324;
assign a21330 = ~a21328 & ~a21320;
assign a21332 = ~a21330 & ~a21316;
assign a21334 = ~a21332 & ~a21314;
assign a21336 = ~a21334 & ~a21310;
assign a21338 = ~a21336 & ~a21308;
assign a21340 = ~a21338 & ~a21304;
assign a21342 = ~a21340 & ~a21302;
assign a21344 = ~a21342 & ~a21298;
assign a21346 = ~a21344 & ~a21296;
assign a21348 = ~a21346 & ~a21292;
assign a21350 = a21346 & a21292;
assign a21352 = ~a21350 & ~a21348;
assign a21354 = ~a21352 & ~a20194;
assign a21356 = ~a21298 & ~a21296;
assign a21358 = ~a21356 & ~a21342;
assign a21360 = a21356 & a21342;
assign a21362 = ~a21360 & ~a21358;
assign a21364 = ~a20220 & ~i510;
assign a21366 = ~a21364 & ~a20152;
assign a21368 = ~a21322 & a21172;
assign a21370 = ~a21368 & ~a21324;
assign a21372 = a21370 & ~a20148;
assign a21374 = ~a21372 & ~a21366;
assign a21376 = ~a21370 & a20148;
assign a21378 = ~a21376 & ~a21374;
assign a21380 = ~a21326 & ~a21320;
assign a21382 = ~a21380 & ~a21324;
assign a21384 = a21380 & a21324;
assign a21386 = ~a21384 & ~a21382;
assign a21388 = a21386 & ~a20140;
assign a21390 = ~a21388 & ~a21378;
assign a21392 = ~a21386 & a20140;
assign a21394 = ~a21392 & ~a21390;
assign a21396 = ~a21316 & ~a21314;
assign a21398 = ~a21396 & ~a21330;
assign a21400 = a21396 & a21330;
assign a21402 = ~a21400 & ~a21398;
assign a21404 = a21402 & ~a20132;
assign a21406 = ~a21404 & ~a21394;
assign a21408 = ~a21402 & a20132;
assign a21410 = ~a21408 & ~a21406;
assign a21412 = ~a21310 & ~a21308;
assign a21414 = ~a21412 & ~a21334;
assign a21416 = a21412 & a21334;
assign a21418 = ~a21416 & ~a21414;
assign a21420 = a21418 & ~a20124;
assign a21422 = ~a21420 & ~a21410;
assign a21424 = ~a21418 & a20124;
assign a21426 = ~a21424 & ~a21422;
assign a21428 = ~a21304 & ~a21302;
assign a21430 = ~a21428 & ~a21338;
assign a21432 = a21428 & a21338;
assign a21434 = ~a21432 & ~a21430;
assign a21436 = a21434 & ~a20116;
assign a21438 = ~a21436 & ~a21426;
assign a21440 = ~a21434 & a20116;
assign a21442 = ~a21440 & ~a21438;
assign a21444 = a21362 & ~a20108;
assign a21446 = ~a21444 & ~a21442;
assign a21448 = ~a21362 & a20108;
assign a21450 = ~a21448 & ~a21446;
assign a21452 = a21352 & a20194;
assign a21454 = ~a21452 & ~a21450;
assign a21456 = ~a21454 & ~a21354;
assign a21458 = ~a21456 & ~a20108;
assign a21460 = ~a21458 & ~a21362;
assign a21462 = a21458 & a21362;
assign a21464 = ~a21456 & ~a20116;
assign a21466 = ~a21464 & ~a21434;
assign a21468 = a21464 & a21434;
assign a21470 = ~a21456 & ~a20124;
assign a21472 = ~a21470 & ~a21418;
assign a21474 = a21470 & a21418;
assign a21476 = ~a21456 & ~a20132;
assign a21478 = ~a21476 & ~a21402;
assign a21480 = a21476 & a21402;
assign a21482 = ~a21456 & ~a20140;
assign a21484 = ~a21482 & ~a21386;
assign a21486 = a21482 & a21386;
assign a21488 = ~a21456 & ~a20148;
assign a21490 = ~a21488 & ~a21370;
assign a21492 = ~a21456 & ~a20152;
assign a21494 = a21492 & ~a21364;
assign a21496 = a21488 & a21370;
assign a21498 = ~a21496 & ~a21494;
assign a21500 = ~a21498 & ~a21490;
assign a21502 = ~a21500 & ~a21486;
assign a21504 = ~a21502 & ~a21484;
assign a21506 = ~a21504 & ~a21480;
assign a21508 = ~a21506 & ~a21478;
assign a21510 = ~a21508 & ~a21474;
assign a21512 = ~a21510 & ~a21472;
assign a21514 = ~a21512 & ~a21468;
assign a21516 = ~a21514 & ~a21466;
assign a21518 = ~a21516 & ~a21462;
assign a21520 = ~a21518 & ~a21460;
assign a21522 = ~a21520 & a21354;
assign a21524 = ~a21462 & ~a21460;
assign a21526 = ~a21524 & ~a21516;
assign a21528 = a21524 & a21516;
assign a21530 = ~a21528 & ~a21526;
assign a21532 = ~a21468 & ~a21466;
assign a21534 = ~a21532 & ~a21512;
assign a21536 = a21532 & a21512;
assign a21538 = ~a21536 & ~a21534;
assign a21540 = ~a21474 & ~a21472;
assign a21542 = ~a21540 & ~a21508;
assign a21544 = a21540 & a21508;
assign a21546 = ~a21544 & ~a21542;
assign a21548 = ~a21480 & ~a21478;
assign a21550 = ~a21548 & ~a21504;
assign a21552 = a21548 & a21504;
assign a21554 = ~a21552 & ~a21550;
assign a21556 = ~a21486 & ~a21484;
assign a21558 = ~a21556 & ~a21500;
assign a21560 = a21556 & a21500;
assign a21562 = ~a21560 & ~a21558;
assign a21564 = ~a21492 & a21364;
assign a21566 = ~a21564 & ~a21494;
assign a21568 = ~a21496 & ~a21490;
assign a21570 = ~a21568 & ~a21494;
assign a21572 = a21568 & a21494;
assign a21574 = ~a21572 & ~a21570;
assign a21576 = ~a21574 & ~a21566;
assign a21578 = a21576 & ~a21562;
assign a21580 = a21578 & ~a21554;
assign a21582 = a21580 & ~a21546;
assign a21584 = a21582 & ~a21538;
assign a21586 = a21584 & ~a21530;
assign a21588 = ~a21586 & a21522;
assign a21590 = a21586 & ~a21522;
assign a21592 = ~a21590 & ~a21588;
assign a21594 = ~a21592 & ~a20208;
assign a21596 = ~a21584 & ~a21530;
assign a21598 = a21584 & a21530;
assign a21600 = ~a21598 & ~a21596;
assign a21602 = ~a21600 & ~a20208;
assign a21604 = ~a21582 & ~a21538;
assign a21606 = a21582 & a21538;
assign a21608 = ~a21606 & ~a21604;
assign a21610 = ~a21608 & ~a20208;
assign a21612 = ~a21580 & ~a21546;
assign a21614 = a21580 & a21546;
assign a21616 = ~a21614 & ~a21612;
assign a21618 = ~a21616 & ~a20208;
assign a21620 = ~a21578 & ~a21554;
assign a21622 = a21578 & a21554;
assign a21624 = ~a21622 & ~a21620;
assign a21626 = ~a21624 & ~a20208;
assign a21628 = ~a21576 & ~a21562;
assign a21630 = a21576 & a21562;
assign a21632 = ~a21630 & ~a21628;
assign a21634 = ~a21632 & ~a20208;
assign a21636 = ~a21574 & a21566;
assign a21638 = a21574 & ~a21566;
assign a21640 = ~a21638 & ~a21636;
assign a21642 = ~a21640 & ~a20208;
assign a21644 = a21566 & ~a20208;
assign a21646 = ~a21644 & ~a14368;
assign a21648 = a21646 & ~a21642;
assign a21650 = a21648 & ~a21634;
assign a21652 = a21650 & ~a21626;
assign a21654 = a21652 & ~a21618;
assign a21656 = a21654 & ~a21610;
assign a21658 = a21656 & ~a21602;
assign a21660 = a21658 & ~a21594;
assign a21662 = a18504 & i542;
assign a21666 = ~a5760 & a5748;
assign a21668 = ~a5748 & i280;
assign a21672 = ~a7316 & a5748;
assign a21674 = ~a5748 & i338;
assign a21676 = ~a21674 & ~a21672;
assign a21678 = ~a7328 & a5748;
assign a21680 = ~a5748 & i340;
assign a21682 = ~a21680 & ~a21678;
assign a21684 = ~a7322 & a5748;
assign a21686 = ~a5748 & i342;
assign a21688 = ~a21686 & ~a21684;
assign a21690 = a21688 & a21682;
assign a21692 = a5748 & ~l886;
assign a21694 = a5748 & l1246;
assign a21696 = ~a5748 & i330;
assign a21698 = ~a21696 & ~a21694;
assign a21700 = ~a21698 & a21692;
assign a21702 = a21700 & a21690;
assign a21704 = a21702 & ~a21676;
assign a21706 = a21704 & ~a21670;
assign a21708 = ~a21704 & l1334;
assign a21710 = ~a21708 & ~a21706;
assign a21712 = ~a21710 & ~a11996;
assign a21714 = a21702 & a21676;
assign a21716 = a21714 & ~a21670;
assign a21718 = ~a21714 & l1336;
assign a21720 = ~a21718 & ~a21716;
assign a21722 = ~a21720 & a11996;
assign a21724 = ~a21722 & ~a21712;
assign a21726 = ~a21724 & l1000;
assign a21728 = a21692 & ~a21682;
assign a21730 = a21728 & a21698;
assign a21732 = a21730 & ~a21676;
assign a21734 = a21732 & ~a21688;
assign a21736 = a21734 & ~a21670;
assign a21738 = ~a21734 & l1338;
assign a21740 = ~a21738 & ~a21736;
assign a21742 = ~a21740 & ~a11996;
assign a21744 = a21730 & a21676;
assign a21746 = a21744 & ~a21688;
assign a21748 = a21746 & ~a21670;
assign a21750 = ~a21746 & l1340;
assign a21752 = ~a21750 & ~a21748;
assign a21754 = ~a21752 & a11996;
assign a21756 = ~a21754 & ~a21742;
assign a21758 = ~a21756 & ~a11974;
assign a21760 = a21732 & a21688;
assign a21762 = a21760 & ~a21670;
assign a21764 = ~a21760 & l1342;
assign a21766 = ~a21764 & ~a21762;
assign a21768 = ~a21766 & ~a11996;
assign a21770 = a21744 & a21688;
assign a21772 = a21770 & ~a21670;
assign a21774 = ~a21770 & l1344;
assign a21776 = ~a21774 & ~a21772;
assign a21778 = ~a21776 & a11996;
assign a21780 = ~a21778 & ~a21768;
assign a21782 = ~a21780 & a11974;
assign a21784 = ~a21782 & ~a21758;
assign a21786 = ~a21784 & l1308;
assign a21788 = a21692 & ~a21688;
assign a21790 = a21698 & a21682;
assign a21792 = a21790 & a21788;
assign a21794 = a21792 & ~a21676;
assign a21796 = a21794 & ~a21670;
assign a21798 = ~a21794 & ~a12954;
assign a21802 = ~a21800 & ~a11996;
assign a21804 = a21792 & a21676;
assign a21806 = a21804 & ~a21670;
assign a21808 = ~a21804 & ~a12962;
assign a21812 = ~a21810 & a11996;
assign a21814 = ~a21812 & ~a21802;
assign a21816 = ~a21814 & ~a11974;
assign a21818 = a21692 & ~a21676;
assign a21820 = a21698 & a21690;
assign a21822 = a21820 & a21818;
assign a21824 = a21822 & ~a21670;
assign a21826 = ~a21822 & ~a12974;
assign a21830 = ~a21828 & ~a11996;
assign a21832 = a21820 & a21692;
assign a21834 = a21832 & a21676;
assign a21836 = a21834 & ~a21670;
assign a21838 = ~a21834 & l1352;
assign a21840 = ~a21838 & ~a21836;
assign a21842 = ~a21840 & a11996;
assign a21844 = ~a21842 & ~a21830;
assign a21846 = ~a21844 & a11974;
assign a21848 = ~a21846 & ~a21816;
assign a21850 = ~a21848 & ~l1308;
assign a21852 = ~a21850 & ~a21786;
assign a21854 = ~a21852 & ~l1000;
assign a21856 = ~a21854 & ~a21726;
assign a21858 = ~a21856 & ~a5624;
assign a21860 = ~a5760 & a5624;
assign a21862 = ~a21860 & ~a21858;
assign a21864 = i356 & ~i354;
assign a21866 = a21864 & i352;
assign a21868 = a21866 & i350;
assign a21870 = a21868 & i348;
assign a21872 = ~a21870 & i346;
assign a21874 = ~a21872 & ~a21862;
assign a21876 = ~a5778 & a5748;
assign a21878 = ~a5748 & i302;
assign a21882 = ~a21880 & a21704;
assign a21884 = ~a21704 & l1354;
assign a21886 = ~a21884 & ~a21882;
assign a21888 = ~a21886 & ~a11996;
assign a21890 = ~a21880 & a21714;
assign a21892 = ~a21714 & l1356;
assign a21894 = ~a21892 & ~a21890;
assign a21896 = ~a21894 & a11996;
assign a21898 = ~a21896 & ~a21888;
assign a21900 = ~a21898 & l1000;
assign a21902 = ~a21880 & a21734;
assign a21904 = ~a21734 & l1358;
assign a21906 = ~a21904 & ~a21902;
assign a21908 = ~a21906 & ~a11996;
assign a21910 = ~a21880 & a21746;
assign a21912 = ~a21746 & l1360;
assign a21914 = ~a21912 & ~a21910;
assign a21916 = ~a21914 & a11996;
assign a21918 = ~a21916 & ~a21908;
assign a21920 = ~a21918 & ~a11974;
assign a21922 = ~a21880 & a21760;
assign a21924 = ~a21760 & l1362;
assign a21926 = ~a21924 & ~a21922;
assign a21928 = ~a21926 & ~a11996;
assign a21930 = ~a21880 & a21770;
assign a21932 = ~a21770 & l1364;
assign a21934 = ~a21932 & ~a21930;
assign a21936 = ~a21934 & a11996;
assign a21938 = ~a21936 & ~a21928;
assign a21940 = ~a21938 & a11974;
assign a21942 = ~a21940 & ~a21920;
assign a21944 = ~a21942 & l1308;
assign a21946 = ~a21880 & a21794;
assign a21948 = ~a21794 & ~a13138;
assign a21952 = ~a21950 & ~a11996;
assign a21954 = ~a21880 & a21804;
assign a21956 = ~a21804 & ~a13146;
assign a21960 = ~a21958 & a11996;
assign a21962 = ~a21960 & ~a21952;
assign a21964 = ~a21962 & ~a11974;
assign a21966 = ~a21880 & a21822;
assign a21968 = ~a21822 & ~a13158;
assign a21972 = ~a21970 & ~a11996;
assign a21974 = ~a21880 & a21834;
assign a21976 = ~a21834 & l1372;
assign a21978 = ~a21976 & ~a21974;
assign a21980 = ~a21978 & a11996;
assign a21982 = ~a21980 & ~a21972;
assign a21984 = ~a21982 & a11974;
assign a21986 = ~a21984 & ~a21964;
assign a21988 = ~a21986 & ~l1308;
assign a21990 = ~a21988 & ~a21944;
assign a21992 = ~a21990 & ~l1000;
assign a21994 = ~a21992 & ~a21900;
assign a21996 = ~a21994 & ~a5624;
assign a21998 = ~a5778 & a5624;
assign a22000 = ~a21998 & ~a21996;
assign a22002 = ~a22000 & ~i348;
assign a22004 = ~a22002 & ~a21874;
assign a22006 = a22000 & i348;
assign a22008 = ~a22006 & ~a22004;
assign a22010 = ~a5796 & a5748;
assign a22012 = ~a5748 & i304;
assign a22016 = ~a22014 & a21704;
assign a22018 = ~a21704 & l1374;
assign a22020 = ~a22018 & ~a22016;
assign a22022 = ~a22020 & ~a11996;
assign a22024 = ~a22014 & a21714;
assign a22026 = ~a21714 & l1376;
assign a22028 = ~a22026 & ~a22024;
assign a22030 = ~a22028 & a11996;
assign a22032 = ~a22030 & ~a22022;
assign a22034 = ~a22032 & l1000;
assign a22036 = ~a22014 & a21734;
assign a22038 = ~a21734 & l1378;
assign a22040 = ~a22038 & ~a22036;
assign a22042 = ~a22040 & ~a11996;
assign a22044 = ~a22014 & a21746;
assign a22046 = ~a21746 & l1380;
assign a22048 = ~a22046 & ~a22044;
assign a22050 = ~a22048 & a11996;
assign a22052 = ~a22050 & ~a22042;
assign a22054 = ~a22052 & ~a11974;
assign a22056 = ~a22014 & a21760;
assign a22058 = ~a21760 & l1382;
assign a22060 = ~a22058 & ~a22056;
assign a22062 = ~a22060 & ~a11996;
assign a22064 = ~a22014 & a21770;
assign a22066 = ~a21770 & l1384;
assign a22068 = ~a22066 & ~a22064;
assign a22070 = ~a22068 & a11996;
assign a22072 = ~a22070 & ~a22062;
assign a22074 = ~a22072 & a11974;
assign a22076 = ~a22074 & ~a22054;
assign a22078 = ~a22076 & l1308;
assign a22080 = ~a22014 & a21794;
assign a22082 = ~a21794 & ~a13328;
assign a22086 = ~a22084 & ~a11996;
assign a22088 = ~a22014 & a21804;
assign a22090 = ~a21804 & ~a13336;
assign a22094 = ~a22092 & a11996;
assign a22096 = ~a22094 & ~a22086;
assign a22098 = ~a22096 & ~a11974;
assign a22100 = ~a22014 & a21822;
assign a22102 = ~a21822 & ~a13348;
assign a22106 = ~a22104 & ~a11996;
assign a22108 = ~a22014 & a21834;
assign a22110 = ~a21834 & l1392;
assign a22112 = ~a22110 & ~a22108;
assign a22114 = ~a22112 & a11996;
assign a22116 = ~a22114 & ~a22106;
assign a22118 = ~a22116 & a11974;
assign a22120 = ~a22118 & ~a22098;
assign a22122 = ~a22120 & ~l1308;
assign a22124 = ~a22122 & ~a22078;
assign a22126 = ~a22124 & ~l1000;
assign a22128 = ~a22126 & ~a22034;
assign a22130 = ~a22128 & ~a5624;
assign a22132 = ~a5796 & a5624;
assign a22134 = ~a22132 & ~a22130;
assign a22136 = ~a22134 & ~i350;
assign a22138 = ~a22136 & ~a22008;
assign a22140 = a22134 & i350;
assign a22142 = ~a22140 & ~a22138;
assign a22144 = ~a5814 & a5748;
assign a22146 = ~a5748 & i306;
assign a22150 = ~a22148 & a21704;
assign a22152 = ~a21704 & l1394;
assign a22154 = ~a22152 & ~a22150;
assign a22156 = ~a22154 & ~a11996;
assign a22158 = ~a22148 & a21714;
assign a22160 = ~a21714 & l1396;
assign a22162 = ~a22160 & ~a22158;
assign a22164 = ~a22162 & a11996;
assign a22166 = ~a22164 & ~a22156;
assign a22168 = ~a22166 & l1000;
assign a22170 = ~a22148 & a21734;
assign a22172 = ~a21734 & l1398;
assign a22174 = ~a22172 & ~a22170;
assign a22176 = ~a22174 & ~a11996;
assign a22178 = ~a22148 & a21746;
assign a22180 = ~a21746 & l1400;
assign a22182 = ~a22180 & ~a22178;
assign a22184 = ~a22182 & a11996;
assign a22186 = ~a22184 & ~a22176;
assign a22188 = ~a22186 & ~a11974;
assign a22190 = ~a22148 & a21760;
assign a22192 = ~a21760 & l1402;
assign a22194 = ~a22192 & ~a22190;
assign a22196 = ~a22194 & ~a11996;
assign a22198 = ~a22148 & a21770;
assign a22200 = ~a21770 & l1404;
assign a22202 = ~a22200 & ~a22198;
assign a22204 = ~a22202 & a11996;
assign a22206 = ~a22204 & ~a22196;
assign a22208 = ~a22206 & a11974;
assign a22210 = ~a22208 & ~a22188;
assign a22212 = ~a22210 & l1308;
assign a22214 = ~a22148 & a21794;
assign a22216 = ~a21794 & ~a13518;
assign a22220 = ~a22218 & ~a11996;
assign a22222 = ~a22148 & a21804;
assign a22224 = ~a21804 & ~a13526;
assign a22228 = ~a22226 & a11996;
assign a22230 = ~a22228 & ~a22220;
assign a22232 = ~a22230 & ~a11974;
assign a22234 = ~a22148 & a21822;
assign a22236 = ~a21822 & ~a13538;
assign a22240 = ~a22238 & ~a11996;
assign a22242 = ~a22148 & a21834;
assign a22244 = ~a21834 & l1412;
assign a22246 = ~a22244 & ~a22242;
assign a22248 = ~a22246 & a11996;
assign a22250 = ~a22248 & ~a22240;
assign a22252 = ~a22250 & a11974;
assign a22254 = ~a22252 & ~a22232;
assign a22256 = ~a22254 & ~l1308;
assign a22258 = ~a22256 & ~a22212;
assign a22260 = ~a22258 & ~l1000;
assign a22262 = ~a22260 & ~a22168;
assign a22264 = ~a22262 & ~a5624;
assign a22266 = ~a5814 & a5624;
assign a22268 = ~a22266 & ~a22264;
assign a22270 = ~a22268 & ~i352;
assign a22272 = ~a22270 & ~a22142;
assign a22274 = a22268 & i352;
assign a22276 = ~a22274 & ~a22272;
assign a22278 = ~a5832 & a5748;
assign a22280 = ~a5748 & i308;
assign a22284 = ~a22282 & a21704;
assign a22286 = ~a21704 & l1414;
assign a22288 = ~a22286 & ~a22284;
assign a22290 = ~a22288 & ~a11996;
assign a22292 = ~a22282 & a21714;
assign a22294 = ~a21714 & l1416;
assign a22296 = ~a22294 & ~a22292;
assign a22298 = ~a22296 & a11996;
assign a22300 = ~a22298 & ~a22290;
assign a22302 = ~a22300 & l1000;
assign a22304 = ~a22282 & a21734;
assign a22306 = ~a21734 & l1418;
assign a22308 = ~a22306 & ~a22304;
assign a22310 = ~a22308 & ~a11996;
assign a22312 = ~a22282 & a21746;
assign a22314 = ~a21746 & l1420;
assign a22316 = ~a22314 & ~a22312;
assign a22318 = ~a22316 & a11996;
assign a22320 = ~a22318 & ~a22310;
assign a22322 = ~a22320 & ~a11974;
assign a22324 = ~a22282 & a21760;
assign a22326 = ~a21760 & l1422;
assign a22328 = ~a22326 & ~a22324;
assign a22330 = ~a22328 & ~a11996;
assign a22332 = ~a22282 & a21770;
assign a22334 = ~a21770 & l1424;
assign a22336 = ~a22334 & ~a22332;
assign a22338 = ~a22336 & a11996;
assign a22340 = ~a22338 & ~a22330;
assign a22342 = ~a22340 & a11974;
assign a22344 = ~a22342 & ~a22322;
assign a22346 = ~a22344 & l1308;
assign a22348 = ~a22282 & a21794;
assign a22350 = ~a21794 & ~a13708;
assign a22354 = ~a22352 & ~a11996;
assign a22356 = ~a22282 & a21804;
assign a22358 = ~a21804 & ~a13716;
assign a22362 = ~a22360 & a11996;
assign a22364 = ~a22362 & ~a22354;
assign a22366 = ~a22364 & ~a11974;
assign a22368 = ~a22282 & a21822;
assign a22370 = ~a21822 & ~a13728;
assign a22374 = ~a22372 & ~a11996;
assign a22376 = ~a22282 & a21834;
assign a22378 = ~a21834 & l1432;
assign a22380 = ~a22378 & ~a22376;
assign a22382 = ~a22380 & a11996;
assign a22384 = ~a22382 & ~a22374;
assign a22386 = ~a22384 & a11974;
assign a22388 = ~a22386 & ~a22366;
assign a22390 = ~a22388 & ~l1308;
assign a22392 = ~a22390 & ~a22346;
assign a22394 = ~a22392 & ~l1000;
assign a22396 = ~a22394 & ~a22302;
assign a22398 = ~a22396 & ~a5624;
assign a22400 = ~a5832 & a5624;
assign a22402 = ~a22400 & ~a22398;
assign a22404 = ~a22402 & ~i356;
assign a22406 = ~a22404 & ~a22276;
assign a22408 = a22402 & i356;
assign a22410 = ~a22408 & ~a22406;
assign a22412 = ~a5850 & a5748;
assign a22414 = ~a5748 & i310;
assign a22418 = ~a22416 & a21704;
assign a22420 = ~a21704 & l1434;
assign a22422 = ~a22420 & ~a22418;
assign a22424 = ~a22422 & ~a11996;
assign a22426 = ~a22416 & a21714;
assign a22428 = ~a21714 & l1436;
assign a22430 = ~a22428 & ~a22426;
assign a22432 = ~a22430 & a11996;
assign a22434 = ~a22432 & ~a22424;
assign a22436 = ~a22434 & l1000;
assign a22438 = ~a22416 & a21734;
assign a22440 = ~a21734 & l1438;
assign a22442 = ~a22440 & ~a22438;
assign a22444 = ~a22442 & ~a11996;
assign a22446 = ~a22416 & a21746;
assign a22448 = ~a21746 & l1440;
assign a22450 = ~a22448 & ~a22446;
assign a22452 = ~a22450 & a11996;
assign a22454 = ~a22452 & ~a22444;
assign a22456 = ~a22454 & ~a11974;
assign a22458 = ~a22416 & a21760;
assign a22460 = ~a21760 & l1442;
assign a22462 = ~a22460 & ~a22458;
assign a22464 = ~a22462 & ~a11996;
assign a22466 = ~a22416 & a21770;
assign a22468 = ~a21770 & l1444;
assign a22470 = ~a22468 & ~a22466;
assign a22472 = ~a22470 & a11996;
assign a22474 = ~a22472 & ~a22464;
assign a22476 = ~a22474 & a11974;
assign a22478 = ~a22476 & ~a22456;
assign a22480 = ~a22478 & l1308;
assign a22482 = ~a22416 & a21794;
assign a22484 = ~a21794 & ~a13886;
assign a22488 = ~a22486 & ~a11996;
assign a22490 = ~a22416 & a21804;
assign a22492 = ~a21804 & ~a13894;
assign a22496 = ~a22494 & a11996;
assign a22498 = ~a22496 & ~a22488;
assign a22500 = ~a22498 & ~a11974;
assign a22502 = ~a22416 & a21822;
assign a22504 = ~a21822 & ~a13906;
assign a22508 = ~a22506 & ~a11996;
assign a22510 = ~a22416 & a21834;
assign a22512 = ~a21834 & l1452;
assign a22514 = ~a22512 & ~a22510;
assign a22516 = ~a22514 & a11996;
assign a22518 = ~a22516 & ~a22508;
assign a22520 = ~a22518 & a11974;
assign a22522 = ~a22520 & ~a22500;
assign a22524 = ~a22522 & ~l1308;
assign a22526 = ~a22524 & ~a22480;
assign a22528 = ~a22526 & ~l1000;
assign a22530 = ~a22528 & ~a22436;
assign a22532 = ~a22530 & ~a5624;
assign a22534 = ~a5850 & a5624;
assign a22536 = ~a22534 & ~a22532;
assign a22538 = ~a22536 & i354;
assign a22540 = ~a22538 & ~a22410;
assign a22542 = a22536 & ~i354;
assign a22544 = ~a22542 & ~a22540;
assign a22546 = ~a5868 & a5748;
assign a22548 = ~a5748 & i358;
assign a22552 = ~a22550 & a21704;
assign a22554 = ~a21704 & l1454;
assign a22556 = ~a22554 & ~a22552;
assign a22558 = ~a22556 & ~a11996;
assign a22560 = ~a22550 & a21714;
assign a22562 = ~a21714 & l1456;
assign a22564 = ~a22562 & ~a22560;
assign a22566 = ~a22564 & a11996;
assign a22568 = ~a22566 & ~a22558;
assign a22570 = ~a22568 & l1000;
assign a22572 = ~a22550 & a21734;
assign a22574 = ~a21734 & l1458;
assign a22576 = ~a22574 & ~a22572;
assign a22578 = ~a22576 & ~a11996;
assign a22580 = ~a22550 & a21746;
assign a22582 = ~a21746 & l1460;
assign a22584 = ~a22582 & ~a22580;
assign a22586 = ~a22584 & a11996;
assign a22588 = ~a22586 & ~a22578;
assign a22590 = ~a22588 & ~a11974;
assign a22592 = ~a22550 & a21760;
assign a22594 = ~a21760 & l1462;
assign a22596 = ~a22594 & ~a22592;
assign a22598 = ~a22596 & ~a11996;
assign a22600 = ~a22550 & a21770;
assign a22602 = ~a21770 & l1464;
assign a22604 = ~a22602 & ~a22600;
assign a22606 = ~a22604 & a11996;
assign a22608 = ~a22606 & ~a22598;
assign a22610 = ~a22608 & a11974;
assign a22612 = ~a22610 & ~a22590;
assign a22614 = ~a22612 & l1308;
assign a22616 = ~a22550 & a21794;
assign a22618 = ~a21794 & ~a14050;
assign a22622 = ~a22620 & ~a11996;
assign a22624 = ~a22550 & a21804;
assign a22626 = ~a21804 & ~a14058;
assign a22630 = ~a22628 & a11996;
assign a22632 = ~a22630 & ~a22622;
assign a22634 = ~a22632 & ~a11974;
assign a22636 = ~a22550 & a21822;
assign a22638 = ~a21822 & l1470;
assign a22640 = ~a22638 & ~a22636;
assign a22642 = ~a22640 & ~a11996;
assign a22644 = ~a22550 & a21834;
assign a22646 = ~a21834 & l1472;
assign a22648 = ~a22646 & ~a22644;
assign a22650 = ~a22648 & a11996;
assign a22652 = ~a22650 & ~a22642;
assign a22654 = ~a22652 & a11974;
assign a22656 = ~a22654 & ~a22634;
assign a22658 = ~a22656 & ~l1308;
assign a22660 = ~a22658 & ~a22614;
assign a22662 = ~a22660 & ~l1000;
assign a22664 = ~a22662 & ~a22570;
assign a22666 = ~a22664 & ~a5624;
assign a22668 = ~a5868 & a5624;
assign a22670 = ~a22668 & ~a22666;
assign a22672 = ~a22670 & ~a22544;
assign a22674 = a22670 & a22544;
assign a22676 = ~a22674 & ~a22672;
assign a22678 = ~a22676 & ~a12380;
assign a22680 = l1060 & ~l998;
assign a22682 = ~l1060 & l998;
assign a22684 = ~a22682 & ~a22680;
assign a22686 = a12836 & ~l972;
assign a22688 = a13020 & ~l1024;
assign a22690 = ~a22688 & ~a22686;
assign a22692 = ~a13020 & l1024;
assign a22694 = ~a22692 & ~a22690;
assign a22696 = a13210 & ~l1092;
assign a22698 = ~a22696 & ~a22694;
assign a22700 = ~a13210 & l1092;
assign a22702 = ~a22700 & ~a22698;
assign a22704 = a13400 & ~l1090;
assign a22706 = ~a22704 & ~a22702;
assign a22708 = ~a13400 & l1090;
assign a22710 = ~a22708 & ~a22706;
assign a22712 = a13590 & ~l1088;
assign a22714 = ~a22712 & ~a22710;
assign a22716 = ~a13590 & l1088;
assign a22718 = ~a22716 & ~a22714;
assign a22720 = a13780 & ~l1086;
assign a22722 = ~a22720 & ~a22718;
assign a22724 = ~a13780 & l1086;
assign a22726 = ~a22724 & ~a22722;
assign a22728 = ~a13958 & ~l1084;
assign a22730 = ~a22728 & ~a22726;
assign a22732 = a13958 & l1084;
assign a22734 = ~a22732 & ~a22730;
assign a22736 = a22734 & ~a22684;
assign a22738 = ~a22734 & a22684;
assign a22740 = ~l1486 & l890;
assign a22742 = a11316 & ~i360;
assign a22744 = ~a22742 & a11318;
assign a22746 = a22744 & ~a11220;
assign a22748 = ~a22746 & ~a22742;
assign a22750 = ~a22748 & ~l890;
assign a22752 = ~a22750 & ~a22740;
assign a22754 = ~a21862 & ~a12836;
assign a22756 = ~a22000 & ~a13020;
assign a22758 = ~a22756 & ~a22754;
assign a22760 = a22000 & a13020;
assign a22762 = ~a22760 & ~a22758;
assign a22764 = ~a22134 & ~a13210;
assign a22766 = ~a22764 & ~a22762;
assign a22768 = a22134 & a13210;
assign a22770 = ~a22768 & ~a22766;
assign a22772 = ~a22268 & ~a13400;
assign a22774 = ~a22772 & ~a22770;
assign a22776 = a22268 & a13400;
assign a22778 = ~a22776 & ~a22774;
assign a22780 = ~a22402 & ~a13590;
assign a22782 = ~a22780 & ~a22778;
assign a22784 = a22402 & a13590;
assign a22786 = ~a22784 & ~a22782;
assign a22788 = ~a22536 & ~a13780;
assign a22790 = ~a22788 & ~a22786;
assign a22792 = a22536 & a13780;
assign a22794 = ~a22792 & ~a22790;
assign a22796 = ~a22670 & a13958;
assign a22798 = ~a22796 & ~a22794;
assign a22800 = a22670 & ~a13958;
assign a22802 = ~a22800 & ~a22798;
assign a22804 = ~a5874 & a5748;
assign a22806 = ~a5748 & i344;
assign a22810 = ~a22808 & a21704;
assign a22812 = ~a21704 & l1314;
assign a22814 = ~a22812 & ~a22810;
assign a22816 = ~a22814 & ~a11996;
assign a22818 = ~a22808 & a21714;
assign a22820 = ~a21714 & l1316;
assign a22822 = ~a22820 & ~a22818;
assign a22824 = ~a22822 & a11996;
assign a22826 = ~a22824 & ~a22816;
assign a22828 = ~a22826 & l1000;
assign a22830 = ~a22808 & a21734;
assign a22832 = ~a21734 & l1318;
assign a22834 = ~a22832 & ~a22830;
assign a22836 = ~a22834 & ~a11996;
assign a22838 = ~a22808 & a21746;
assign a22840 = ~a21746 & l1320;
assign a22842 = ~a22840 & ~a22838;
assign a22844 = ~a22842 & a11996;
assign a22846 = ~a22844 & ~a22836;
assign a22848 = ~a22846 & ~a11974;
assign a22850 = ~a22808 & a21760;
assign a22852 = ~a21760 & l1322;
assign a22854 = ~a22852 & ~a22850;
assign a22856 = ~a22854 & ~a11996;
assign a22858 = ~a22808 & a21770;
assign a22860 = ~a21770 & l1324;
assign a22862 = ~a22860 & ~a22858;
assign a22864 = ~a22862 & a11996;
assign a22866 = ~a22864 & ~a22856;
assign a22868 = ~a22866 & a11974;
assign a22870 = ~a22868 & ~a22848;
assign a22872 = ~a22870 & l1308;
assign a22874 = ~a22808 & a21794;
assign a22876 = ~a21794 & l1326;
assign a22878 = ~a22876 & ~a22874;
assign a22880 = ~a22878 & ~a11996;
assign a22882 = ~a22808 & a21804;
assign a22884 = ~a21804 & l1328;
assign a22886 = ~a22884 & ~a22882;
assign a22888 = ~a22886 & a11996;
assign a22890 = ~a22888 & ~a22880;
assign a22892 = ~a22890 & ~a11974;
assign a22894 = ~a22808 & a21822;
assign a22896 = ~a21822 & l1330;
assign a22898 = ~a22896 & ~a22894;
assign a22900 = ~a22898 & ~a11996;
assign a22902 = ~a22808 & a21834;
assign a22904 = ~a21834 & l1332;
assign a22906 = ~a22904 & ~a22902;
assign a22908 = ~a22906 & a11996;
assign a22910 = ~a22908 & ~a22900;
assign a22912 = ~a22910 & a11974;
assign a22914 = ~a22912 & ~a22892;
assign a22916 = ~a22914 & ~l1308;
assign a22918 = ~a22916 & ~a22872;
assign a22920 = ~a22918 & ~l1000;
assign a22922 = ~a22920 & ~a22828;
assign a22924 = ~a22922 & ~a5624;
assign a22926 = ~a5874 & a5624;
assign a22928 = ~a22926 & ~a22924;
assign a22930 = ~a22928 & ~l998;
assign a22932 = a22928 & l998;
assign a22934 = ~a22932 & ~a22930;
assign a22936 = a22934 & ~a22802;
assign a22938 = a12328 & ~a11996;
assign a22940 = ~a12328 & a11996;
assign a22942 = a12268 & ~a11974;
assign a22944 = ~a12268 & a11974;
assign a22946 = a12206 & l1308;
assign a22948 = ~a12206 & ~l1308;
assign a22950 = a9026 & l1000;
assign a22952 = ~a9026 & ~l1000;
assign a22954 = ~a22952 & ~a22950;
assign a22956 = a22954 & ~a22948;
assign a22958 = a22956 & ~a22946;
assign a22960 = a22958 & ~a22944;
assign a22962 = a22960 & ~a22942;
assign a22964 = a22962 & ~a22940;
assign a22966 = a22964 & ~a22938;
assign a22968 = ~a11996 & l968;
assign a22970 = a11996 & l970;
assign a22972 = ~a22970 & ~a22968;
assign a22974 = ~a22972 & l1000;
assign a22976 = ~a11996 & l966;
assign a22978 = a11996 & l964;
assign a22980 = ~a22978 & ~a22976;
assign a22982 = ~a22980 & ~a11974;
assign a22984 = ~a11996 & l962;
assign a22986 = a11996 & l960;
assign a22988 = ~a22986 & ~a22984;
assign a22990 = ~a22988 & a11974;
assign a22992 = ~a22990 & ~a22982;
assign a22994 = ~a22992 & l1308;
assign a22996 = ~a11996 & a5606;
assign a22998 = a11996 & a5600;
assign a23000 = ~a22998 & ~a22996;
assign a23002 = ~a23000 & ~a11974;
assign a23004 = ~a11996 & a5594;
assign a23006 = a11996 & a5568;
assign a23008 = ~a23006 & ~a23004;
assign a23010 = ~a23008 & a11974;
assign a23012 = ~a23010 & ~a23002;
assign a23014 = ~a23012 & ~l1308;
assign a23016 = ~a23014 & ~a22994;
assign a23018 = ~a23016 & ~l1000;
assign a23020 = ~a23018 & ~a22974;
assign a23022 = ~a23020 & ~a22966;
assign a23024 = ~a23022 & ~a5760;
assign a23026 = ~a11996 & a11974;
assign a23028 = a23026 & l1000;
assign a23030 = a23028 & ~l1308;
assign a23032 = ~a11996 & ~a11974;
assign a23034 = a23032 & l1308;
assign a23036 = ~a23034 & l1000;
assign a23038 = a23034 & ~l1000;
assign a23040 = ~a23038 & ~a23036;
assign a23042 = ~a21710 & a11996;
assign a23044 = ~a21720 & ~a11996;
assign a23046 = ~a23044 & ~a23042;
assign a23048 = ~a23046 & ~a23040;
assign a23050 = ~a23032 & l1308;
assign a23052 = a23032 & ~l1308;
assign a23054 = ~a23052 & ~a23050;
assign a23056 = a11996 & ~a11974;
assign a23058 = ~a23056 & ~a23026;
assign a23060 = ~a21740 & a11996;
assign a23062 = ~a21752 & ~a11996;
assign a23064 = ~a23062 & ~a23060;
assign a23066 = ~a23064 & ~a23058;
assign a23068 = ~a21766 & a11996;
assign a23070 = ~a21776 & ~a11996;
assign a23072 = ~a23070 & ~a23068;
assign a23074 = ~a23072 & a23058;
assign a23076 = ~a23074 & ~a23066;
assign a23078 = ~a23076 & ~a23054;
assign a23080 = ~a21800 & a11996;
assign a23082 = ~a21810 & ~a11996;
assign a23084 = ~a23082 & ~a23080;
assign a23086 = ~a23084 & ~a23058;
assign a23088 = ~a21828 & a11996;
assign a23090 = ~a21840 & ~a11996;
assign a23092 = ~a23090 & ~a23088;
assign a23094 = ~a23092 & a23058;
assign a23096 = ~a23094 & ~a23086;
assign a23098 = ~a23096 & a23054;
assign a23100 = ~a23098 & ~a23078;
assign a23102 = ~a23100 & a23040;
assign a23104 = ~a23102 & ~a23048;
assign a23106 = ~a23104 & ~a23030;
assign a23108 = a23030 & ~a21840;
assign a23110 = ~a23108 & ~a23106;
assign a23112 = ~a23110 & a23022;
assign a23114 = ~a23112 & ~a23024;
assign a23116 = ~a23114 & ~a12836;
assign a23118 = ~a23022 & ~a5778;
assign a23120 = ~a21886 & a11996;
assign a23122 = ~a21894 & ~a11996;
assign a23124 = ~a23122 & ~a23120;
assign a23126 = ~a23124 & ~a23040;
assign a23128 = ~a21906 & a11996;
assign a23130 = ~a21914 & ~a11996;
assign a23132 = ~a23130 & ~a23128;
assign a23134 = ~a23132 & ~a23058;
assign a23136 = ~a21926 & a11996;
assign a23138 = ~a21934 & ~a11996;
assign a23140 = ~a23138 & ~a23136;
assign a23142 = ~a23140 & a23058;
assign a23144 = ~a23142 & ~a23134;
assign a23146 = ~a23144 & ~a23054;
assign a23148 = ~a21950 & a11996;
assign a23150 = ~a21958 & ~a11996;
assign a23152 = ~a23150 & ~a23148;
assign a23154 = ~a23152 & ~a23058;
assign a23156 = ~a21970 & a11996;
assign a23158 = ~a21978 & ~a11996;
assign a23160 = ~a23158 & ~a23156;
assign a23162 = ~a23160 & a23058;
assign a23164 = ~a23162 & ~a23154;
assign a23166 = ~a23164 & a23054;
assign a23168 = ~a23166 & ~a23146;
assign a23170 = ~a23168 & a23040;
assign a23172 = ~a23170 & ~a23126;
assign a23174 = ~a23172 & ~a23030;
assign a23176 = a23030 & ~a21978;
assign a23178 = ~a23176 & ~a23174;
assign a23180 = ~a23178 & a23022;
assign a23182 = ~a23180 & ~a23118;
assign a23184 = ~a23182 & ~a13020;
assign a23186 = ~a23184 & ~a23116;
assign a23188 = a23182 & a13020;
assign a23190 = ~a23188 & ~a23186;
assign a23192 = ~a23022 & ~a5796;
assign a23194 = ~a22020 & a11996;
assign a23196 = ~a22028 & ~a11996;
assign a23198 = ~a23196 & ~a23194;
assign a23200 = ~a23198 & ~a23040;
assign a23202 = ~a22040 & a11996;
assign a23204 = ~a22048 & ~a11996;
assign a23206 = ~a23204 & ~a23202;
assign a23208 = ~a23206 & ~a23058;
assign a23210 = ~a22060 & a11996;
assign a23212 = ~a22068 & ~a11996;
assign a23214 = ~a23212 & ~a23210;
assign a23216 = ~a23214 & a23058;
assign a23218 = ~a23216 & ~a23208;
assign a23220 = ~a23218 & ~a23054;
assign a23222 = ~a22084 & a11996;
assign a23224 = ~a22092 & ~a11996;
assign a23226 = ~a23224 & ~a23222;
assign a23228 = ~a23226 & ~a23058;
assign a23230 = ~a22104 & a11996;
assign a23232 = ~a22112 & ~a11996;
assign a23234 = ~a23232 & ~a23230;
assign a23236 = ~a23234 & a23058;
assign a23238 = ~a23236 & ~a23228;
assign a23240 = ~a23238 & a23054;
assign a23242 = ~a23240 & ~a23220;
assign a23244 = ~a23242 & a23040;
assign a23246 = ~a23244 & ~a23200;
assign a23248 = ~a23246 & ~a23030;
assign a23250 = a23030 & ~a22112;
assign a23252 = ~a23250 & ~a23248;
assign a23254 = ~a23252 & a23022;
assign a23256 = ~a23254 & ~a23192;
assign a23258 = ~a23256 & ~a13210;
assign a23260 = ~a23258 & ~a23190;
assign a23262 = a23256 & a13210;
assign a23264 = ~a23262 & ~a23260;
assign a23266 = ~a23022 & ~a5814;
assign a23268 = ~a22154 & a11996;
assign a23270 = ~a22162 & ~a11996;
assign a23272 = ~a23270 & ~a23268;
assign a23274 = ~a23272 & ~a23040;
assign a23276 = ~a22174 & a11996;
assign a23278 = ~a22182 & ~a11996;
assign a23280 = ~a23278 & ~a23276;
assign a23282 = ~a23280 & ~a23058;
assign a23284 = ~a22194 & a11996;
assign a23286 = ~a22202 & ~a11996;
assign a23288 = ~a23286 & ~a23284;
assign a23290 = ~a23288 & a23058;
assign a23292 = ~a23290 & ~a23282;
assign a23294 = ~a23292 & ~a23054;
assign a23296 = ~a22218 & a11996;
assign a23298 = ~a22226 & ~a11996;
assign a23300 = ~a23298 & ~a23296;
assign a23302 = ~a23300 & ~a23058;
assign a23304 = ~a22238 & a11996;
assign a23306 = ~a22246 & ~a11996;
assign a23308 = ~a23306 & ~a23304;
assign a23310 = ~a23308 & a23058;
assign a23312 = ~a23310 & ~a23302;
assign a23314 = ~a23312 & a23054;
assign a23316 = ~a23314 & ~a23294;
assign a23318 = ~a23316 & a23040;
assign a23320 = ~a23318 & ~a23274;
assign a23322 = ~a23320 & ~a23030;
assign a23324 = a23030 & ~a22246;
assign a23326 = ~a23324 & ~a23322;
assign a23328 = ~a23326 & a23022;
assign a23330 = ~a23328 & ~a23266;
assign a23332 = ~a23330 & ~a13400;
assign a23334 = ~a23332 & ~a23264;
assign a23336 = a23330 & a13400;
assign a23338 = ~a23336 & ~a23334;
assign a23340 = ~a23022 & ~a5832;
assign a23342 = ~a22288 & a11996;
assign a23344 = ~a22296 & ~a11996;
assign a23346 = ~a23344 & ~a23342;
assign a23348 = ~a23346 & ~a23040;
assign a23350 = ~a22308 & a11996;
assign a23352 = ~a22316 & ~a11996;
assign a23354 = ~a23352 & ~a23350;
assign a23356 = ~a23354 & ~a23058;
assign a23358 = ~a22328 & a11996;
assign a23360 = ~a22336 & ~a11996;
assign a23362 = ~a23360 & ~a23358;
assign a23364 = ~a23362 & a23058;
assign a23366 = ~a23364 & ~a23356;
assign a23368 = ~a23366 & ~a23054;
assign a23370 = ~a22352 & a11996;
assign a23372 = ~a22360 & ~a11996;
assign a23374 = ~a23372 & ~a23370;
assign a23376 = ~a23374 & ~a23058;
assign a23378 = ~a22372 & a11996;
assign a23380 = ~a22380 & ~a11996;
assign a23382 = ~a23380 & ~a23378;
assign a23384 = ~a23382 & a23058;
assign a23386 = ~a23384 & ~a23376;
assign a23388 = ~a23386 & a23054;
assign a23390 = ~a23388 & ~a23368;
assign a23392 = ~a23390 & a23040;
assign a23394 = ~a23392 & ~a23348;
assign a23396 = ~a23394 & ~a23030;
assign a23398 = a23030 & ~a22380;
assign a23400 = ~a23398 & ~a23396;
assign a23402 = ~a23400 & a23022;
assign a23404 = ~a23402 & ~a23340;
assign a23406 = ~a23404 & ~a13590;
assign a23408 = ~a23406 & ~a23338;
assign a23410 = a23404 & a13590;
assign a23412 = ~a23410 & ~a23408;
assign a23414 = ~a23022 & ~a5850;
assign a23416 = ~a22422 & a11996;
assign a23418 = ~a22430 & ~a11996;
assign a23420 = ~a23418 & ~a23416;
assign a23422 = ~a23420 & ~a23040;
assign a23424 = ~a22442 & a11996;
assign a23426 = ~a22450 & ~a11996;
assign a23428 = ~a23426 & ~a23424;
assign a23430 = ~a23428 & ~a23058;
assign a23432 = ~a22462 & a11996;
assign a23434 = ~a22470 & ~a11996;
assign a23436 = ~a23434 & ~a23432;
assign a23438 = ~a23436 & a23058;
assign a23440 = ~a23438 & ~a23430;
assign a23442 = ~a23440 & ~a23054;
assign a23444 = ~a22486 & a11996;
assign a23446 = ~a22494 & ~a11996;
assign a23448 = ~a23446 & ~a23444;
assign a23450 = ~a23448 & ~a23058;
assign a23452 = ~a22506 & a11996;
assign a23454 = ~a22514 & ~a11996;
assign a23456 = ~a23454 & ~a23452;
assign a23458 = ~a23456 & a23058;
assign a23460 = ~a23458 & ~a23450;
assign a23462 = ~a23460 & a23054;
assign a23464 = ~a23462 & ~a23442;
assign a23466 = ~a23464 & a23040;
assign a23468 = ~a23466 & ~a23422;
assign a23470 = ~a23468 & ~a23030;
assign a23472 = a23030 & ~a22514;
assign a23474 = ~a23472 & ~a23470;
assign a23476 = ~a23474 & a23022;
assign a23478 = ~a23476 & ~a23414;
assign a23480 = ~a23478 & ~a13780;
assign a23482 = ~a23480 & ~a23412;
assign a23484 = a23478 & a13780;
assign a23486 = ~a23484 & ~a23482;
assign a23488 = ~a23022 & ~a5868;
assign a23490 = ~a22556 & a11996;
assign a23492 = ~a22564 & ~a11996;
assign a23494 = ~a23492 & ~a23490;
assign a23496 = ~a23494 & ~a23040;
assign a23498 = ~a22576 & a11996;
assign a23500 = ~a22584 & ~a11996;
assign a23502 = ~a23500 & ~a23498;
assign a23504 = ~a23502 & ~a23058;
assign a23506 = ~a22596 & a11996;
assign a23508 = ~a22604 & ~a11996;
assign a23510 = ~a23508 & ~a23506;
assign a23512 = ~a23510 & a23058;
assign a23514 = ~a23512 & ~a23504;
assign a23516 = ~a23514 & ~a23054;
assign a23518 = ~a22620 & a11996;
assign a23520 = ~a22628 & ~a11996;
assign a23522 = ~a23520 & ~a23518;
assign a23524 = ~a23522 & ~a23058;
assign a23526 = ~a22640 & a11996;
assign a23528 = ~a22648 & ~a11996;
assign a23530 = ~a23528 & ~a23526;
assign a23532 = ~a23530 & a23058;
assign a23534 = ~a23532 & ~a23524;
assign a23536 = ~a23534 & a23054;
assign a23538 = ~a23536 & ~a23516;
assign a23540 = ~a23538 & a23040;
assign a23542 = ~a23540 & ~a23496;
assign a23544 = ~a23542 & ~a23030;
assign a23546 = a23030 & ~a22648;
assign a23548 = ~a23546 & ~a23544;
assign a23550 = ~a23548 & a23022;
assign a23552 = ~a23550 & ~a23488;
assign a23554 = ~a23552 & a13958;
assign a23556 = ~a23554 & ~a23486;
assign a23558 = a23552 & ~a13958;
assign a23560 = ~a23558 & ~a23556;
assign a23562 = ~a23022 & ~a5874;
assign a23564 = ~a22814 & a11996;
assign a23566 = ~a22822 & ~a11996;
assign a23568 = ~a23566 & ~a23564;
assign a23570 = ~a23568 & ~a23040;
assign a23572 = ~a22834 & a11996;
assign a23574 = ~a22842 & ~a11996;
assign a23576 = ~a23574 & ~a23572;
assign a23578 = ~a23576 & ~a23058;
assign a23580 = ~a22854 & a11996;
assign a23582 = ~a22862 & ~a11996;
assign a23584 = ~a23582 & ~a23580;
assign a23586 = ~a23584 & a23058;
assign a23588 = ~a23586 & ~a23578;
assign a23590 = ~a23588 & ~a23054;
assign a23592 = ~a22878 & a11996;
assign a23594 = ~a22886 & ~a11996;
assign a23596 = ~a23594 & ~a23592;
assign a23598 = ~a23596 & ~a23058;
assign a23600 = ~a22898 & a11996;
assign a23602 = ~a22906 & ~a11996;
assign a23604 = ~a23602 & ~a23600;
assign a23606 = ~a23604 & a23058;
assign a23608 = ~a23606 & ~a23598;
assign a23610 = ~a23608 & a23054;
assign a23612 = ~a23610 & ~a23590;
assign a23614 = ~a23612 & a23040;
assign a23616 = ~a23614 & ~a23570;
assign a23618 = ~a23616 & ~a23030;
assign a23620 = a23030 & ~a22906;
assign a23622 = ~a23620 & ~a23618;
assign a23624 = ~a23622 & a23022;
assign a23626 = ~a23624 & ~a23562;
assign a23628 = a23626 & ~a22928;
assign a23630 = ~a23626 & a22928;
assign a23632 = ~a23630 & ~a23628;
assign a23634 = a23632 & a23560;
assign a23636 = a23634 & a22936;
assign a23638 = ~a23626 & ~l998;
assign a23640 = a23626 & l998;
assign a23642 = ~a23640 & ~a23638;
assign a23644 = a23642 & a23560;
assign a23646 = ~a23644 & ~a22936;
assign a23648 = ~a23646 & ~a23632;
assign a23650 = ~a23648 & ~a23636;
assign a23652 = ~a23650 & ~a22752;
assign a23654 = a23652 & ~a22738;
assign a23656 = a23654 & ~a22736;
assign a23658 = ~l1488 & l890;
assign a23660 = a11960 & i362;
assign a23662 = a23660 & ~i364;
assign a23664 = ~a23662 & ~l890;
assign a23666 = ~a23664 & ~a23658;
assign a23668 = a12380 & ~l886;
assign a23670 = a23668 & a23666;
assign a23672 = a23670 & a22752;
assign a23674 = a22934 & a22802;
assign a23676 = ~a23674 & ~a23672;
assign a23678 = a23676 & ~a23656;
assign a23680 = ~a21872 & a12836;
assign a23682 = a13020 & ~i348;
assign a23684 = ~a23682 & ~a23680;
assign a23686 = ~a13020 & i348;
assign a23688 = ~a23686 & ~a23684;
assign a23690 = a13210 & ~i350;
assign a23692 = ~a23690 & ~a23688;
assign a23694 = ~a13210 & i350;
assign a23696 = ~a23694 & ~a23692;
assign a23698 = a13400 & ~i352;
assign a23700 = ~a23698 & ~a23696;
assign a23702 = ~a13400 & i352;
assign a23704 = ~a23702 & ~a23700;
assign a23706 = a13590 & ~i356;
assign a23708 = ~a23706 & ~a23704;
assign a23710 = ~a13590 & i356;
assign a23712 = ~a23710 & ~a23708;
assign a23714 = a13780 & i354;
assign a23716 = ~a23714 & ~a23712;
assign a23718 = ~a13780 & ~i354;
assign a23720 = ~a23718 & ~a23716;
assign a23722 = ~a23720 & ~a13958;
assign a23724 = a23720 & a13958;
assign a23726 = ~a23724 & ~a23722;
assign a23728 = ~a23726 & ~a23678;
assign a23730 = a23678 & ~a13958;
assign a23732 = ~a23730 & ~a23728;
assign a23734 = ~a23732 & a12380;
assign a23738 = ~a21692 & ~a12380;
assign a23740 = ~a23738 & ~l886;
assign a23744 = a8986 & a8954;
assign a23746 = a23744 & a8924;
assign a23748 = a23746 & a8870;
assign a23750 = a8814 & l1516;
assign a23752 = a8818 & l1518;
assign a23754 = ~a23752 & ~a23750;
assign a23756 = l1544 & l1172;
assign a23758 = ~a23756 & a23754;
assign a23760 = a8974 & ~a8860;
assign a23762 = a23760 & a8826;
assign a23764 = ~a23762 & ~a23758;
assign a23766 = a23762 & a23758;
assign a23768 = ~a23766 & ~a23764;
assign a23770 = ~a23768 & ~a8812;
assign a23772 = a8812 & l1546;
assign a23774 = ~a23772 & ~a23770;
assign a23776 = ~a23774 & ~l1582;
assign a23778 = a23774 & l1582;
assign a23780 = ~a23778 & ~a23776;
assign a23782 = a23780 & a23748;
assign a23784 = ~a8954 & l968;
assign a23786 = a8954 & l970;
assign a23788 = ~a23786 & ~a23784;
assign a23790 = ~a23788 & ~a8870;
assign a23792 = ~a8954 & l966;
assign a23794 = a8954 & l964;
assign a23796 = ~a23794 & ~a23792;
assign a23798 = ~a23796 & ~a8986;
assign a23800 = ~a8954 & l962;
assign a23802 = a8954 & l960;
assign a23804 = ~a23802 & ~a23800;
assign a23806 = ~a23804 & a8986;
assign a23808 = ~a23806 & ~a23798;
assign a23810 = ~a23808 & ~a8924;
assign a23812 = ~a8954 & a5606;
assign a23814 = a8954 & a5600;
assign a23816 = ~a23814 & ~a23812;
assign a23818 = ~a23816 & ~a8986;
assign a23820 = ~a8954 & a5594;
assign a23822 = a8954 & a5568;
assign a23824 = ~a23822 & ~a23820;
assign a23826 = ~a23824 & a8986;
assign a23828 = ~a23826 & ~a23818;
assign a23830 = ~a23828 & a8924;
assign a23832 = ~a23830 & ~a23810;
assign a23834 = ~a23832 & a8870;
assign a23836 = ~a23834 & ~a23790;
assign a23838 = ~a8954 & ~l1550;
assign a23840 = a8954 & l1550;
assign a23842 = ~a8986 & ~l1552;
assign a23844 = a8986 & l1552;
assign a23846 = ~a8924 & ~l1556;
assign a23848 = a8924 & l1556;
assign a23850 = ~a8870 & ~l1554;
assign a23852 = a8870 & l1554;
assign a23854 = ~a23852 & ~a23850;
assign a23856 = a23854 & ~a23848;
assign a23858 = a23856 & ~a23846;
assign a23860 = a23858 & ~a23844;
assign a23862 = a23860 & ~a23842;
assign a23864 = a23862 & ~a23840;
assign a23866 = a23864 & ~a23838;
assign a23868 = ~a14546 & l1560;
assign a23870 = a14546 & l1564;
assign a23872 = ~a23870 & ~a23868;
assign a23874 = ~a23872 & l1558;
assign a23876 = ~a14546 & l1548;
assign a23878 = a14546 & l1570;
assign a23880 = ~a23878 & ~a23876;
assign a23882 = ~a23880 & ~a14552;
assign a23884 = ~a14546 & l1572;
assign a23886 = a14546 & l1574;
assign a23888 = ~a23886 & ~a23884;
assign a23890 = ~a23888 & a14552;
assign a23892 = ~a23890 & ~a23882;
assign a23894 = ~a23892 & l1566;
assign a23896 = ~a14546 & l1576;
assign a23898 = a14546 & l1578;
assign a23900 = ~a23898 & ~a23896;
assign a23902 = ~a23900 & ~a14552;
assign a23904 = ~a14546 & l1580;
assign a23906 = a14546 & l1582;
assign a23908 = ~a23906 & ~a23904;
assign a23910 = ~a23908 & a14552;
assign a23912 = ~a23910 & ~a23902;
assign a23914 = ~a23912 & ~l1566;
assign a23916 = ~a23914 & ~a23894;
assign a23918 = ~a23916 & ~l1558;
assign a23920 = ~a23918 & ~a23874;
assign a23922 = a23920 & ~a23774;
assign a23924 = ~a23920 & a23774;
assign a23926 = ~a23924 & ~a23922;
assign a23928 = ~a23926 & ~a23866;
assign a23930 = a23928 & ~a23836;
assign a23932 = a23930 & ~a23780;
assign a23934 = ~a23932 & ~a23782;
assign a23936 = ~a23934 & l948;
assign a23938 = ~a17442 & ~l1330;
assign a23940 = a17442 & l1330;
assign a23942 = ~a23940 & ~a23938;
assign a23944 = a17466 & ~a12974;
assign a23946 = a17484 & ~a13158;
assign a23948 = ~a23946 & ~a23944;
assign a23950 = ~a17484 & a13158;
assign a23952 = ~a23950 & ~a23948;
assign a23954 = a17508 & ~a13348;
assign a23956 = ~a23954 & ~a23952;
assign a23958 = ~a17508 & a13348;
assign a23960 = ~a23958 & ~a23956;
assign a23962 = a17532 & ~a13538;
assign a23964 = ~a23962 & ~a23960;
assign a23966 = ~a17532 & a13538;
assign a23968 = ~a23966 & ~a23964;
assign a23970 = a17556 & ~a13728;
assign a23972 = ~a23970 & ~a23968;
assign a23974 = ~a17556 & a13728;
assign a23976 = ~a23974 & ~a23972;
assign a23978 = a17580 & ~a13906;
assign a23980 = ~a23978 & ~a23976;
assign a23982 = ~a17580 & a13906;
assign a23984 = ~a23982 & ~a23980;
assign a23986 = a17606 & l1470;
assign a23988 = ~a23986 & ~a23984;
assign a23990 = ~a17606 & ~l1470;
assign a23992 = ~a23990 & ~a23988;
assign a23994 = ~a23992 & a23942;
assign a23996 = ~a17466 & a12974;
assign a23998 = ~a23996 & ~a23950;
assign a24000 = ~a23998 & ~a23946;
assign a24002 = ~a24000 & ~a23958;
assign a24004 = ~a24002 & ~a23954;
assign a24006 = ~a24004 & ~a23966;
assign a24008 = ~a24006 & ~a23962;
assign a24010 = ~a24008 & ~a23974;
assign a24012 = ~a24010 & ~a23970;
assign a24014 = ~a24012 & ~a23982;
assign a24016 = ~a24014 & ~a23978;
assign a24018 = ~a24016 & ~a23990;
assign a24020 = ~a24018 & ~a23986;
assign a24022 = ~a24020 & ~a23942;
assign a24024 = ~a24022 & ~a23994;
assign a24026 = a5748 & l1530;
assign a24028 = ~a5748 & i420;
assign a24030 = ~a24028 & ~a24026;
assign a24032 = ~a24030 & a21822;
assign a24034 = ~a21822 & l1580;
assign a24036 = ~a24034 & ~a24032;
assign a24038 = ~a24036 & ~l1582;
assign a24040 = a24036 & l1582;
assign a24042 = ~a24040 & ~a24038;
assign a24044 = a24042 & ~a24024;
assign a24046 = a24044 & a17436;
assign a24048 = a24046 & a5594;
assign a24050 = ~a24048 & a5568;
assign a24052 = ~a24050 & ~a21834;
assign a24054 = ~a24052 & ~l886;
assign a24058 = ~a23774 & ~l1580;
assign a24060 = a23774 & l1580;
assign a24062 = ~a24060 & ~a24058;
assign a24064 = a8986 & a8924;
assign a24066 = a24064 & a8870;
assign a24068 = a24066 & a24062;
assign a24070 = ~a24062 & a23930;
assign a24072 = ~a24070 & ~a24068;
assign a24074 = ~a24072 & l948;
assign a24076 = ~a17442 & ~l1328;
assign a24078 = a17442 & l1328;
assign a24080 = ~a24078 & ~a24076;
assign a24082 = a17466 & ~a12962;
assign a24084 = a17484 & ~a13146;
assign a24086 = ~a24084 & ~a24082;
assign a24088 = ~a17484 & a13146;
assign a24090 = ~a24088 & ~a24086;
assign a24092 = a17508 & ~a13336;
assign a24094 = ~a24092 & ~a24090;
assign a24096 = ~a17508 & a13336;
assign a24098 = ~a24096 & ~a24094;
assign a24100 = a17532 & ~a13526;
assign a24102 = ~a24100 & ~a24098;
assign a24104 = ~a17532 & a13526;
assign a24106 = ~a24104 & ~a24102;
assign a24108 = a17556 & ~a13716;
assign a24110 = ~a24108 & ~a24106;
assign a24112 = ~a17556 & a13716;
assign a24114 = ~a24112 & ~a24110;
assign a24116 = a17580 & ~a13894;
assign a24118 = ~a24116 & ~a24114;
assign a24120 = ~a17580 & a13894;
assign a24122 = ~a24120 & ~a24118;
assign a24124 = a17606 & ~a14058;
assign a24126 = ~a24124 & ~a24122;
assign a24128 = ~a17606 & a14058;
assign a24130 = ~a24128 & ~a24126;
assign a24132 = ~a24130 & a24080;
assign a24134 = ~a17466 & a12962;
assign a24136 = ~a24134 & ~a24088;
assign a24138 = ~a24136 & ~a24084;
assign a24140 = ~a24138 & ~a24096;
assign a24142 = ~a24140 & ~a24092;
assign a24144 = ~a24142 & ~a24104;
assign a24146 = ~a24144 & ~a24100;
assign a24148 = ~a24146 & ~a24112;
assign a24150 = ~a24148 & ~a24108;
assign a24152 = ~a24150 & ~a24120;
assign a24154 = ~a24152 & ~a24116;
assign a24156 = ~a24154 & ~a24128;
assign a24158 = ~a24156 & ~a24124;
assign a24160 = ~a24158 & ~a24080;
assign a24162 = ~a24160 & ~a24132;
assign a24164 = ~a24030 & a21804;
assign a24166 = ~a21804 & l1578;
assign a24168 = ~a24166 & ~a24164;
assign a24170 = ~a24168 & ~l1580;
assign a24172 = a24168 & l1580;
assign a24174 = ~a24172 & ~a24170;
assign a24176 = a24174 & ~a24162;
assign a24178 = a24176 & a17436;
assign a24180 = a24178 & a5600;
assign a24182 = ~a24180 & a5594;
assign a24184 = ~a24182 & ~a21822;
assign a24186 = ~a24184 & ~l886;
assign a24190 = ~a23774 & ~l1578;
assign a24192 = a23774 & l1578;
assign a24194 = ~a24192 & ~a24190;
assign a24196 = ~a8986 & ~a8954;
assign a24198 = a8924 & a8870;
assign a24200 = a24198 & ~a24196;
assign a24202 = a24200 & a24194;
assign a24204 = ~a24194 & a23930;
assign a24206 = ~a24204 & ~a24202;
assign a24208 = ~a24206 & l948;
assign a24210 = ~a17442 & ~l1326;
assign a24212 = a17442 & l1326;
assign a24214 = ~a24212 & ~a24210;
assign a24216 = a17466 & ~a12954;
assign a24218 = a17484 & ~a13138;
assign a24220 = ~a24218 & ~a24216;
assign a24222 = ~a17484 & a13138;
assign a24224 = ~a24222 & ~a24220;
assign a24226 = a17508 & ~a13328;
assign a24228 = ~a24226 & ~a24224;
assign a24230 = ~a17508 & a13328;
assign a24232 = ~a24230 & ~a24228;
assign a24234 = a17532 & ~a13518;
assign a24236 = ~a24234 & ~a24232;
assign a24238 = ~a17532 & a13518;
assign a24240 = ~a24238 & ~a24236;
assign a24242 = a17556 & ~a13708;
assign a24244 = ~a24242 & ~a24240;
assign a24246 = ~a17556 & a13708;
assign a24248 = ~a24246 & ~a24244;
assign a24250 = a17580 & ~a13886;
assign a24252 = ~a24250 & ~a24248;
assign a24254 = ~a17580 & a13886;
assign a24256 = ~a24254 & ~a24252;
assign a24258 = a17606 & ~a14050;
assign a24260 = ~a24258 & ~a24256;
assign a24262 = ~a17606 & a14050;
assign a24264 = ~a24262 & ~a24260;
assign a24266 = ~a24264 & a24214;
assign a24268 = ~a17466 & a12954;
assign a24270 = ~a24268 & ~a24222;
assign a24272 = ~a24270 & ~a24218;
assign a24274 = ~a24272 & ~a24230;
assign a24276 = ~a24274 & ~a24226;
assign a24278 = ~a24276 & ~a24238;
assign a24280 = ~a24278 & ~a24234;
assign a24282 = ~a24280 & ~a24246;
assign a24284 = ~a24282 & ~a24242;
assign a24286 = ~a24284 & ~a24254;
assign a24288 = ~a24286 & ~a24250;
assign a24290 = ~a24288 & ~a24262;
assign a24292 = ~a24290 & ~a24258;
assign a24294 = ~a24292 & ~a24214;
assign a24296 = ~a24294 & ~a24266;
assign a24298 = ~a24030 & a21794;
assign a24300 = ~a21794 & l1576;
assign a24302 = ~a24300 & ~a24298;
assign a24304 = ~a24302 & ~l1578;
assign a24306 = a24302 & l1578;
assign a24308 = ~a24306 & ~a24304;
assign a24310 = a24308 & ~a24296;
assign a24312 = a24310 & a17436;
assign a24314 = a24312 & a5606;
assign a24316 = ~a24314 & a5600;
assign a24318 = ~a24316 & ~a21804;
assign a24320 = ~a24318 & ~l886;
assign a24324 = ~a23774 & ~l1576;
assign a24326 = a23774 & l1576;
assign a24328 = ~a24326 & ~a24324;
assign a24330 = a24328 & a24198;
assign a24332 = ~a24328 & a23930;
assign a24334 = ~a24332 & ~a24330;
assign a24336 = ~a24334 & l948;
assign a24338 = ~a17442 & ~l1324;
assign a24340 = a17442 & l1324;
assign a24342 = ~a24340 & ~a24338;
assign a24344 = a17466 & l1344;
assign a24346 = a17484 & l1364;
assign a24348 = ~a24346 & ~a24344;
assign a24350 = ~a17484 & ~l1364;
assign a24352 = ~a24350 & ~a24348;
assign a24354 = a17508 & l1384;
assign a24356 = ~a24354 & ~a24352;
assign a24358 = ~a17508 & ~l1384;
assign a24360 = ~a24358 & ~a24356;
assign a24362 = a17532 & l1404;
assign a24364 = ~a24362 & ~a24360;
assign a24366 = ~a17532 & ~l1404;
assign a24368 = ~a24366 & ~a24364;
assign a24370 = a17556 & l1424;
assign a24372 = ~a24370 & ~a24368;
assign a24374 = ~a17556 & ~l1424;
assign a24376 = ~a24374 & ~a24372;
assign a24378 = a17580 & l1444;
assign a24380 = ~a24378 & ~a24376;
assign a24382 = ~a17580 & ~l1444;
assign a24384 = ~a24382 & ~a24380;
assign a24386 = a17606 & l1464;
assign a24388 = ~a24386 & ~a24384;
assign a24390 = ~a17606 & ~l1464;
assign a24392 = ~a24390 & ~a24388;
assign a24394 = ~a24392 & a24342;
assign a24396 = ~a17466 & ~l1344;
assign a24398 = ~a24396 & ~a24350;
assign a24400 = ~a24398 & ~a24346;
assign a24402 = ~a24400 & ~a24358;
assign a24404 = ~a24402 & ~a24354;
assign a24406 = ~a24404 & ~a24366;
assign a24408 = ~a24406 & ~a24362;
assign a24410 = ~a24408 & ~a24374;
assign a24412 = ~a24410 & ~a24370;
assign a24414 = ~a24412 & ~a24382;
assign a24416 = ~a24414 & ~a24378;
assign a24418 = ~a24416 & ~a24390;
assign a24420 = ~a24418 & ~a24386;
assign a24422 = ~a24420 & ~a24342;
assign a24424 = ~a24422 & ~a24394;
assign a24426 = ~a24030 & a21770;
assign a24428 = ~a21770 & l1574;
assign a24430 = ~a24428 & ~a24426;
assign a24432 = ~a24430 & ~l1576;
assign a24434 = a24430 & l1576;
assign a24436 = ~a24434 & ~a24432;
assign a24438 = a24436 & ~a24424;
assign a24440 = a24438 & a17436;
assign a24442 = a24440 & l960;
assign a24444 = ~a24442 & a5606;
assign a24446 = ~a24444 & ~a21794;
assign a24448 = ~a24446 & ~l886;
assign a24452 = ~a23774 & ~l1574;
assign a24454 = a23774 & l1574;
assign a24456 = ~a24454 & ~a24452;
assign a24458 = ~a23744 & ~a8924;
assign a24460 = ~a24458 & a8870;
assign a24462 = a24460 & a24456;
assign a24464 = ~a24456 & a23930;
assign a24466 = ~a24464 & ~a24462;
assign a24468 = ~a24466 & l948;
assign a24470 = ~a17442 & ~l1322;
assign a24472 = a17442 & l1322;
assign a24474 = ~a24472 & ~a24470;
assign a24476 = a17466 & l1342;
assign a24478 = a17484 & l1362;
assign a24480 = ~a24478 & ~a24476;
assign a24482 = ~a17484 & ~l1362;
assign a24484 = ~a24482 & ~a24480;
assign a24486 = a17508 & l1382;
assign a24488 = ~a24486 & ~a24484;
assign a24490 = ~a17508 & ~l1382;
assign a24492 = ~a24490 & ~a24488;
assign a24494 = a17532 & l1402;
assign a24496 = ~a24494 & ~a24492;
assign a24498 = ~a17532 & ~l1402;
assign a24500 = ~a24498 & ~a24496;
assign a24502 = a17556 & l1422;
assign a24504 = ~a24502 & ~a24500;
assign a24506 = ~a17556 & ~l1422;
assign a24508 = ~a24506 & ~a24504;
assign a24510 = a17580 & l1442;
assign a24512 = ~a24510 & ~a24508;
assign a24514 = ~a17580 & ~l1442;
assign a24516 = ~a24514 & ~a24512;
assign a24518 = a17606 & l1462;
assign a24520 = ~a24518 & ~a24516;
assign a24522 = ~a17606 & ~l1462;
assign a24524 = ~a24522 & ~a24520;
assign a24526 = ~a24524 & a24474;
assign a24528 = ~a17466 & ~l1342;
assign a24530 = ~a24528 & ~a24482;
assign a24532 = ~a24530 & ~a24478;
assign a24534 = ~a24532 & ~a24490;
assign a24536 = ~a24534 & ~a24486;
assign a24538 = ~a24536 & ~a24498;
assign a24540 = ~a24538 & ~a24494;
assign a24542 = ~a24540 & ~a24506;
assign a24544 = ~a24542 & ~a24502;
assign a24546 = ~a24544 & ~a24514;
assign a24548 = ~a24546 & ~a24510;
assign a24550 = ~a24548 & ~a24522;
assign a24552 = ~a24550 & ~a24518;
assign a24554 = ~a24552 & ~a24474;
assign a24556 = ~a24554 & ~a24526;
assign a24558 = ~a24030 & a21760;
assign a24560 = ~a21760 & l1572;
assign a24562 = ~a24560 & ~a24558;
assign a24564 = ~a24562 & ~l1574;
assign a24566 = a24562 & l1574;
assign a24568 = ~a24566 & ~a24564;
assign a24570 = a24568 & ~a24556;
assign a24572 = a24570 & a17436;
assign a24574 = a24572 & l962;
assign a24576 = ~a24574 & l960;
assign a24578 = ~a24576 & ~a21770;
assign a24580 = ~a24578 & ~l886;
assign a24584 = ~a23774 & ~l1572;
assign a24586 = a23774 & l1572;
assign a24588 = ~a24586 & ~a24584;
assign a24590 = ~a8986 & ~a8924;
assign a24592 = ~a24590 & a8870;
assign a24594 = a24592 & a24588;
assign a24596 = ~a24588 & a23930;
assign a24598 = ~a24596 & ~a24594;
assign a24600 = ~a24598 & l948;
assign a24602 = ~a17442 & ~l1320;
assign a24604 = a17442 & l1320;
assign a24606 = ~a24604 & ~a24602;
assign a24608 = a17466 & l1340;
assign a24610 = a17484 & l1360;
assign a24612 = ~a24610 & ~a24608;
assign a24614 = ~a17484 & ~l1360;
assign a24616 = ~a24614 & ~a24612;
assign a24618 = a17508 & l1380;
assign a24620 = ~a24618 & ~a24616;
assign a24622 = ~a17508 & ~l1380;
assign a24624 = ~a24622 & ~a24620;
assign a24626 = a17532 & l1400;
assign a24628 = ~a24626 & ~a24624;
assign a24630 = ~a17532 & ~l1400;
assign a24632 = ~a24630 & ~a24628;
assign a24634 = a17556 & l1420;
assign a24636 = ~a24634 & ~a24632;
assign a24638 = ~a17556 & ~l1420;
assign a24640 = ~a24638 & ~a24636;
assign a24642 = a17580 & l1440;
assign a24644 = ~a24642 & ~a24640;
assign a24646 = ~a17580 & ~l1440;
assign a24648 = ~a24646 & ~a24644;
assign a24650 = a17606 & l1460;
assign a24652 = ~a24650 & ~a24648;
assign a24654 = ~a17606 & ~l1460;
assign a24656 = ~a24654 & ~a24652;
assign a24658 = ~a24656 & a24606;
assign a24660 = ~a17466 & ~l1340;
assign a24662 = ~a24660 & ~a24614;
assign a24664 = ~a24662 & ~a24610;
assign a24666 = ~a24664 & ~a24622;
assign a24668 = ~a24666 & ~a24618;
assign a24670 = ~a24668 & ~a24630;
assign a24672 = ~a24670 & ~a24626;
assign a24674 = ~a24672 & ~a24638;
assign a24676 = ~a24674 & ~a24634;
assign a24678 = ~a24676 & ~a24646;
assign a24680 = ~a24678 & ~a24642;
assign a24682 = ~a24680 & ~a24654;
assign a24684 = ~a24682 & ~a24650;
assign a24686 = ~a24684 & ~a24606;
assign a24688 = ~a24686 & ~a24658;
assign a24690 = ~a24030 & a21746;
assign a24692 = ~a21746 & l1570;
assign a24694 = ~a24692 & ~a24690;
assign a24696 = ~a24694 & ~l1572;
assign a24698 = a24694 & l1572;
assign a24700 = ~a24698 & ~a24696;
assign a24702 = a24700 & ~a24688;
assign a24704 = a24702 & a17436;
assign a24706 = a24704 & l964;
assign a24708 = ~a24706 & l962;
assign a24710 = ~a24708 & ~a21760;
assign a24712 = ~a24710 & ~l886;
assign a24716 = ~a23774 & ~l1570;
assign a24718 = a23774 & l1570;
assign a24720 = ~a24718 & ~a24716;
assign a24722 = a24196 & ~a8924;
assign a24724 = ~a24722 & a8870;
assign a24726 = a24724 & a24720;
assign a24728 = ~a24720 & a23930;
assign a24730 = ~a24728 & ~a24726;
assign a24732 = ~a24730 & l948;
assign a24734 = ~a17442 & ~l1318;
assign a24736 = a17442 & l1318;
assign a24738 = ~a24736 & ~a24734;
assign a24740 = a17466 & l1338;
assign a24742 = a17484 & l1358;
assign a24744 = ~a24742 & ~a24740;
assign a24746 = ~a17484 & ~l1358;
assign a24748 = ~a24746 & ~a24744;
assign a24750 = a17508 & l1378;
assign a24752 = ~a24750 & ~a24748;
assign a24754 = ~a17508 & ~l1378;
assign a24756 = ~a24754 & ~a24752;
assign a24758 = a17532 & l1398;
assign a24760 = ~a24758 & ~a24756;
assign a24762 = ~a17532 & ~l1398;
assign a24764 = ~a24762 & ~a24760;
assign a24766 = a17556 & l1418;
assign a24768 = ~a24766 & ~a24764;
assign a24770 = ~a17556 & ~l1418;
assign a24772 = ~a24770 & ~a24768;
assign a24774 = a17580 & l1438;
assign a24776 = ~a24774 & ~a24772;
assign a24778 = ~a17580 & ~l1438;
assign a24780 = ~a24778 & ~a24776;
assign a24782 = a17606 & l1458;
assign a24784 = ~a24782 & ~a24780;
assign a24786 = ~a17606 & ~l1458;
assign a24788 = ~a24786 & ~a24784;
assign a24790 = ~a24788 & a24738;
assign a24792 = ~a17466 & ~l1338;
assign a24794 = ~a24792 & ~a24746;
assign a24796 = ~a24794 & ~a24742;
assign a24798 = ~a24796 & ~a24754;
assign a24800 = ~a24798 & ~a24750;
assign a24802 = ~a24800 & ~a24762;
assign a24804 = ~a24802 & ~a24758;
assign a24806 = ~a24804 & ~a24770;
assign a24808 = ~a24806 & ~a24766;
assign a24810 = ~a24808 & ~a24778;
assign a24812 = ~a24810 & ~a24774;
assign a24814 = ~a24812 & ~a24786;
assign a24816 = ~a24814 & ~a24782;
assign a24818 = ~a24816 & ~a24738;
assign a24820 = ~a24818 & ~a24790;
assign a24822 = ~a24030 & a21734;
assign a24824 = ~a21734 & l1548;
assign a24826 = ~a24824 & ~a24822;
assign a24828 = ~a24826 & ~l1570;
assign a24830 = a24826 & l1570;
assign a24832 = ~a24830 & ~a24828;
assign a24834 = a24832 & ~a24820;
assign a24836 = a24834 & a17436;
assign a24838 = a24836 & l966;
assign a24840 = ~a24838 & l964;
assign a24842 = ~a24840 & ~a21746;
assign a24844 = ~a24842 & ~l886;
assign a24848 = ~a23774 & ~l1548;
assign a24850 = a23774 & l1548;
assign a24852 = ~a24850 & ~a24848;
assign a24854 = a24852 & a8870;
assign a24856 = ~a24852 & a23930;
assign a24858 = ~a24856 & ~a24854;
assign a24860 = ~a24858 & l948;
assign a24862 = ~a17442 & ~l1316;
assign a24864 = a17442 & l1316;
assign a24866 = ~a24864 & ~a24862;
assign a24868 = a17466 & l1336;
assign a24870 = a17484 & l1356;
assign a24872 = ~a24870 & ~a24868;
assign a24874 = ~a17484 & ~l1356;
assign a24876 = ~a24874 & ~a24872;
assign a24878 = a17508 & l1376;
assign a24880 = ~a24878 & ~a24876;
assign a24882 = ~a17508 & ~l1376;
assign a24884 = ~a24882 & ~a24880;
assign a24886 = a17532 & l1396;
assign a24888 = ~a24886 & ~a24884;
assign a24890 = ~a17532 & ~l1396;
assign a24892 = ~a24890 & ~a24888;
assign a24894 = a17556 & l1416;
assign a24896 = ~a24894 & ~a24892;
assign a24898 = ~a17556 & ~l1416;
assign a24900 = ~a24898 & ~a24896;
assign a24902 = a17580 & l1436;
assign a24904 = ~a24902 & ~a24900;
assign a24906 = ~a17580 & ~l1436;
assign a24908 = ~a24906 & ~a24904;
assign a24910 = a17606 & l1456;
assign a24912 = ~a24910 & ~a24908;
assign a24914 = ~a17606 & ~l1456;
assign a24916 = ~a24914 & ~a24912;
assign a24918 = ~a24916 & a24866;
assign a24920 = ~a17466 & ~l1336;
assign a24922 = ~a24920 & ~a24874;
assign a24924 = ~a24922 & ~a24870;
assign a24926 = ~a24924 & ~a24882;
assign a24928 = ~a24926 & ~a24878;
assign a24930 = ~a24928 & ~a24890;
assign a24932 = ~a24930 & ~a24886;
assign a24934 = ~a24932 & ~a24898;
assign a24936 = ~a24934 & ~a24894;
assign a24938 = ~a24936 & ~a24906;
assign a24940 = ~a24938 & ~a24902;
assign a24942 = ~a24940 & ~a24914;
assign a24944 = ~a24942 & ~a24910;
assign a24946 = ~a24944 & ~a24866;
assign a24948 = ~a24946 & ~a24918;
assign a24950 = ~a24030 & a21714;
assign a24952 = ~a21714 & l1564;
assign a24954 = ~a24952 & ~a24950;
assign a24956 = ~a24954 & ~l1548;
assign a24958 = a24954 & l1548;
assign a24960 = ~a24958 & ~a24956;
assign a24962 = a24960 & ~a24948;
assign a24964 = a24962 & a17436;
assign a24966 = a24964 & l970;
assign a24968 = ~a24966 & l966;
assign a24970 = ~a24968 & ~a21734;
assign a24972 = ~a24970 & ~l886;
assign a24976 = ~a23774 & ~l1560;
assign a24978 = a23774 & l1560;
assign a24980 = ~a24978 & ~a24976;
assign a24982 = ~a24064 & ~a8870;
assign a24984 = ~a24982 & a24980;
assign a24986 = ~a24980 & a23930;
assign a24988 = ~a24986 & ~a24984;
assign a24990 = ~a24988 & l948;
assign a24992 = ~a21704 & ~l968;
assign a24994 = ~a17442 & ~l1332;
assign a24996 = a17442 & l1332;
assign a24998 = ~a24996 & ~a24994;
assign a25000 = a17466 & l1352;
assign a25002 = a17484 & l1372;
assign a25004 = ~a25002 & ~a25000;
assign a25006 = ~a17484 & ~l1372;
assign a25008 = ~a25006 & ~a25004;
assign a25010 = a17508 & l1392;
assign a25012 = ~a25010 & ~a25008;
assign a25014 = ~a17508 & ~l1392;
assign a25016 = ~a25014 & ~a25012;
assign a25018 = a17532 & l1412;
assign a25020 = ~a25018 & ~a25016;
assign a25022 = ~a17532 & ~l1412;
assign a25024 = ~a25022 & ~a25020;
assign a25026 = a17556 & l1432;
assign a25028 = ~a25026 & ~a25024;
assign a25030 = ~a17556 & ~l1432;
assign a25032 = ~a25030 & ~a25028;
assign a25034 = a17580 & l1452;
assign a25036 = ~a25034 & ~a25032;
assign a25038 = ~a17580 & ~l1452;
assign a25040 = ~a25038 & ~a25036;
assign a25042 = a17606 & l1472;
assign a25044 = ~a25042 & ~a25040;
assign a25046 = ~a17606 & ~l1472;
assign a25048 = ~a25046 & ~a25044;
assign a25050 = ~a25048 & a24998;
assign a25052 = ~a17466 & ~l1352;
assign a25054 = ~a25052 & ~a25006;
assign a25056 = ~a25054 & ~a25002;
assign a25058 = ~a25056 & ~a25014;
assign a25060 = ~a25058 & ~a25010;
assign a25062 = ~a25060 & ~a25022;
assign a25064 = ~a25062 & ~a25018;
assign a25066 = ~a25064 & ~a25030;
assign a25068 = ~a25066 & ~a25026;
assign a25070 = ~a25068 & ~a25038;
assign a25072 = ~a25070 & ~a25034;
assign a25074 = ~a25072 & ~a25046;
assign a25076 = ~a25074 & ~a25042;
assign a25078 = ~a25076 & ~a24998;
assign a25080 = ~a25078 & ~a25050;
assign a25082 = ~a24030 & a21834;
assign a25084 = ~a21834 & l1582;
assign a25086 = ~a25084 & ~a25082;
assign a25088 = ~a25086 & ~l1560;
assign a25090 = a25086 & l1560;
assign a25092 = ~a25090 & ~a25088;
assign a25094 = ~a25092 & ~a25080;
assign a25096 = a25094 & a17436;
assign a25098 = a25096 & a5568;
assign a25100 = ~a25098 & ~a24992;
assign a25102 = ~a25100 & ~a21704;
assign a25104 = ~a25102 & ~l886;
assign a25108 = ~a23746 & ~a8870;
assign a25110 = ~a23774 & ~l1564;
assign a25112 = a23774 & l1564;
assign a25114 = ~a25112 & ~a25110;
assign a25116 = a25114 & ~a25108;
assign a25118 = ~a25114 & a23930;
assign a25120 = ~a25118 & ~a25116;
assign a25122 = ~a25120 & l948;
assign a25124 = ~a17442 & ~l1314;
assign a25126 = a17442 & l1314;
assign a25128 = ~a25126 & ~a25124;
assign a25130 = a17466 & l1334;
assign a25132 = a17484 & l1354;
assign a25134 = ~a25132 & ~a25130;
assign a25136 = ~a17484 & ~l1354;
assign a25138 = ~a25136 & ~a25134;
assign a25140 = a17508 & l1374;
assign a25142 = ~a25140 & ~a25138;
assign a25144 = ~a17508 & ~l1374;
assign a25146 = ~a25144 & ~a25142;
assign a25148 = a17532 & l1394;
assign a25150 = ~a25148 & ~a25146;
assign a25152 = ~a17532 & ~l1394;
assign a25154 = ~a25152 & ~a25150;
assign a25156 = a17556 & l1414;
assign a25158 = ~a25156 & ~a25154;
assign a25160 = ~a17556 & ~l1414;
assign a25162 = ~a25160 & ~a25158;
assign a25164 = a17580 & l1434;
assign a25166 = ~a25164 & ~a25162;
assign a25168 = ~a17580 & ~l1434;
assign a25170 = ~a25168 & ~a25166;
assign a25172 = a17606 & l1454;
assign a25174 = ~a25172 & ~a25170;
assign a25176 = ~a17606 & ~l1454;
assign a25178 = ~a25176 & ~a25174;
assign a25180 = ~a25178 & a25128;
assign a25182 = ~a17466 & ~l1334;
assign a25184 = ~a25182 & ~a25136;
assign a25186 = ~a25184 & ~a25132;
assign a25188 = ~a25186 & ~a25144;
assign a25190 = ~a25188 & ~a25140;
assign a25192 = ~a25190 & ~a25152;
assign a25194 = ~a25192 & ~a25148;
assign a25196 = ~a25194 & ~a25160;
assign a25198 = ~a25196 & ~a25156;
assign a25200 = ~a25198 & ~a25168;
assign a25202 = ~a25200 & ~a25164;
assign a25204 = ~a25202 & ~a25176;
assign a25206 = ~a25204 & ~a25172;
assign a25208 = ~a25206 & ~a25128;
assign a25210 = ~a25208 & ~a25180;
assign a25212 = ~a24030 & a21704;
assign a25214 = ~a21704 & l1560;
assign a25216 = ~a25214 & ~a25212;
assign a25218 = ~a25216 & ~l1564;
assign a25220 = a25216 & l1564;
assign a25222 = ~a25220 & ~a25218;
assign a25224 = a25222 & ~a25210;
assign a25226 = a25224 & l968;
assign a25228 = a25226 & a17436;
assign a25230 = ~a25228 & l970;
assign a25232 = ~a25230 & ~a21714;
assign a25234 = ~a25232 & ~l886;
assign a25238 = ~a17436 & l972;
assign a25240 = ~a25238 & ~a17468;
assign a25244 = ~a17296 & i278;
assign a25246 = ~a17330 & i284;
assign a25248 = ~a25246 & ~a25244;
assign a25250 = a17330 & ~i284;
assign a25252 = ~a25250 & ~a25248;
assign a25254 = ~a17378 & i300;
assign a25256 = ~a25254 & ~a25252;
assign a25258 = a17378 & ~i300;
assign a25260 = ~a25258 & ~a25256;
assign a25262 = a25260 & ~a17396;
assign a25264 = a25262 & l1072;
assign a25266 = a25264 & l1076;
assign a25268 = a25266 & l1028;
assign a25270 = ~a25268 & l1026;
assign a25272 = a25268 & ~l1026;
assign a25274 = ~a25272 & ~a25270;
assign a25276 = ~a17296 & ~i278;
assign a25278 = a17296 & i278;
assign a25280 = ~a25278 & ~a25276;
assign a25282 = ~a17330 & ~i284;
assign a25284 = a17330 & i284;
assign a25286 = ~a25284 & ~a25282;
assign a25288 = ~a25286 & ~a25244;
assign a25290 = a25286 & a25244;
assign a25292 = ~a25290 & ~a25288;
assign a25294 = ~a25292 & ~a25280;
assign a25296 = ~a17378 & ~i300;
assign a25298 = a17378 & i300;
assign a25300 = ~a25298 & ~a25296;
assign a25302 = ~a25300 & ~a25252;
assign a25304 = a25300 & a25252;
assign a25306 = ~a25304 & ~a25302;
assign a25308 = ~a25306 & a25294;
assign a25310 = ~a25260 & ~a17396;
assign a25312 = a25260 & a17396;
assign a25314 = ~a25312 & ~a25310;
assign a25316 = ~a25314 & a25308;
assign a25318 = ~a25262 & l1072;
assign a25320 = a25262 & ~l1072;
assign a25322 = ~a25320 & ~a25318;
assign a25324 = ~a25322 & a25316;
assign a25326 = ~a25264 & l1076;
assign a25328 = a25264 & ~l1076;
assign a25330 = ~a25328 & ~a25326;
assign a25332 = ~a25330 & a25324;
assign a25334 = ~a25266 & l1028;
assign a25336 = a25266 & ~l1028;
assign a25338 = ~a25336 & ~a25334;
assign a25340 = ~a25338 & a25332;
assign a25342 = ~a25340 & ~a25274;
assign a25344 = a25340 & a25274;
assign a25346 = ~a25344 & ~a25342;
assign a25348 = ~a25346 & a17272;
assign a25350 = a21692 & a5624;
assign a25352 = ~a21670 & i278;
assign a25354 = ~a21880 & i284;
assign a25356 = ~a25354 & ~a25352;
assign a25358 = a21880 & ~i284;
assign a25360 = ~a25358 & ~a25356;
assign a25362 = ~a22014 & i300;
assign a25364 = ~a25362 & ~a25360;
assign a25366 = a22014 & ~i300;
assign a25368 = ~a25366 & ~a25364;
assign a25370 = a25368 & ~a22148;
assign a25372 = a25370 & ~a22282;
assign a25374 = a25372 & ~a22416;
assign a25376 = a25374 & ~a22550;
assign a25378 = ~a25376 & ~a22808;
assign a25380 = a25376 & a22808;
assign a25382 = ~a25380 & ~a25378;
assign a25384 = ~a25382 & a25350;
assign a25386 = ~a5624 & ~l976;
assign a25388 = l1032 & i278;
assign a25390 = l1064 & i284;
assign a25392 = ~a25390 & ~a25388;
assign a25394 = ~l1064 & ~i284;
assign a25396 = ~a25394 & ~a25392;
assign a25398 = l1066 & i300;
assign a25400 = ~a25398 & ~a25396;
assign a25402 = ~l1066 & ~i300;
assign a25404 = ~a25402 & ~a25400;
assign a25406 = a25404 & l1070;
assign a25408 = a25406 & l1074;
assign a25410 = a25408 & l1078;
assign a25412 = a25410 & l2058;
assign a25414 = ~a25412 & l2060;
assign a25416 = a25412 & ~l2060;
assign a25418 = ~a25416 & ~a25414;
assign a25420 = l1032 & ~i278;
assign a25422 = ~l1032 & i278;
assign a25424 = ~a25422 & ~a25420;
assign a25426 = l1064 & ~i284;
assign a25428 = ~l1064 & i284;
assign a25430 = ~a25428 & ~a25426;
assign a25432 = ~a25430 & ~a25388;
assign a25434 = a25430 & a25388;
assign a25436 = ~a25434 & ~a25432;
assign a25438 = ~a25436 & ~a25424;
assign a25440 = l1066 & ~i300;
assign a25442 = ~l1066 & i300;
assign a25444 = ~a25442 & ~a25440;
assign a25446 = ~a25444 & ~a25396;
assign a25448 = a25444 & a25396;
assign a25450 = ~a25448 & ~a25446;
assign a25452 = ~a25450 & a25438;
assign a25454 = ~a25404 & l1070;
assign a25456 = a25404 & ~l1070;
assign a25458 = ~a25456 & ~a25454;
assign a25460 = ~a25458 & a25452;
assign a25462 = ~a25406 & l1074;
assign a25464 = a25406 & ~l1074;
assign a25466 = ~a25464 & ~a25462;
assign a25468 = ~a25466 & a25460;
assign a25470 = ~a25408 & l1078;
assign a25472 = a25408 & ~l1078;
assign a25474 = ~a25472 & ~a25470;
assign a25476 = ~a25474 & a25468;
assign a25478 = ~a25410 & l2058;
assign a25480 = a25410 & ~l2058;
assign a25482 = ~a25480 & ~a25478;
assign a25484 = ~a25482 & a25476;
assign a25486 = ~a25484 & ~a25418;
assign a25488 = a25484 & a25418;
assign a25490 = ~a25488 & ~a25486;
assign a25492 = ~a25490 & a25386;
assign a25494 = ~a25386 & l1026;
assign a25496 = ~a25494 & ~a25492;
assign a25498 = ~a25496 & ~a25350;
assign a25500 = ~a25498 & ~a25384;
assign a25502 = ~a25500 & ~a17272;
assign a25504 = ~a25502 & ~a25348;
assign a25506 = ~a25504 & ~l978;
assign a25508 = a25504 & l978;
assign a25510 = ~a25508 & ~a25506;
assign a25512 = a25280 & a17272;
assign a25514 = ~a21670 & ~i278;
assign a25516 = a21670 & i278;
assign a25518 = ~a25516 & ~a25514;
assign a25520 = ~a25518 & a25350;
assign a25522 = a25424 & a25386;
assign a25524 = ~a25386 & ~a17296;
assign a25526 = ~a25524 & ~a25522;
assign a25528 = ~a25526 & ~a25350;
assign a25530 = ~a25528 & ~a25520;
assign a25532 = ~a25530 & ~a17272;
assign a25536 = a25534 & ~a6254;
assign a25538 = ~a25292 & a25280;
assign a25540 = a25292 & ~a25280;
assign a25542 = ~a25540 & ~a25538;
assign a25544 = ~a25542 & a17272;
assign a25546 = ~a21880 & ~i284;
assign a25548 = a21880 & i284;
assign a25550 = ~a25548 & ~a25546;
assign a25552 = ~a25550 & ~a25352;
assign a25554 = a25550 & a25352;
assign a25556 = ~a25554 & ~a25552;
assign a25558 = ~a25556 & a25350;
assign a25560 = ~a25436 & a25424;
assign a25562 = a25436 & ~a25424;
assign a25564 = ~a25562 & ~a25560;
assign a25566 = ~a25564 & a25386;
assign a25568 = ~a25386 & ~a17330;
assign a25570 = ~a25568 & ~a25566;
assign a25572 = ~a25570 & ~a25350;
assign a25574 = ~a25572 & ~a25558;
assign a25576 = ~a25574 & ~a17272;
assign a25580 = a25578 & ~a6262;
assign a25582 = ~a25580 & ~a25536;
assign a25584 = ~a25578 & a6262;
assign a25586 = ~a25584 & ~a25582;
assign a25588 = ~a25306 & ~a25294;
assign a25590 = a25306 & a25294;
assign a25592 = ~a25590 & ~a25588;
assign a25594 = ~a25592 & a17272;
assign a25596 = ~a22014 & ~i300;
assign a25598 = a22014 & i300;
assign a25600 = ~a25598 & ~a25596;
assign a25602 = ~a25600 & ~a25360;
assign a25604 = a25600 & a25360;
assign a25606 = ~a25604 & ~a25602;
assign a25608 = ~a25606 & a25350;
assign a25610 = ~a25450 & ~a25438;
assign a25612 = a25450 & a25438;
assign a25614 = ~a25612 & ~a25610;
assign a25616 = ~a25614 & a25386;
assign a25618 = ~a25386 & ~a17378;
assign a25620 = ~a25618 & ~a25616;
assign a25622 = ~a25620 & ~a25350;
assign a25624 = ~a25622 & ~a25608;
assign a25626 = ~a25624 & ~a17272;
assign a25630 = a25628 & ~a6270;
assign a25632 = ~a25630 & ~a25586;
assign a25634 = ~a25628 & a6270;
assign a25636 = ~a25634 & ~a25632;
assign a25638 = ~a25314 & ~a25308;
assign a25640 = a25314 & a25308;
assign a25642 = ~a25640 & ~a25638;
assign a25644 = ~a25642 & a17272;
assign a25646 = ~a25368 & ~a22148;
assign a25648 = a25368 & a22148;
assign a25650 = ~a25648 & ~a25646;
assign a25652 = ~a25650 & a25350;
assign a25654 = ~a25458 & ~a25452;
assign a25656 = a25458 & a25452;
assign a25658 = ~a25656 & ~a25654;
assign a25660 = ~a25658 & a25386;
assign a25662 = ~a25386 & ~a17396;
assign a25664 = ~a25662 & ~a25660;
assign a25666 = ~a25664 & ~a25350;
assign a25668 = ~a25666 & ~a25652;
assign a25670 = ~a25668 & ~a17272;
assign a25674 = a25672 & ~a6278;
assign a25676 = ~a25674 & ~a25636;
assign a25678 = ~a25672 & a6278;
assign a25680 = ~a25678 & ~a25676;
assign a25682 = ~a25322 & ~a25316;
assign a25684 = a25322 & a25316;
assign a25686 = ~a25684 & ~a25682;
assign a25688 = ~a25686 & a17272;
assign a25690 = ~a25370 & ~a22282;
assign a25692 = a25370 & a22282;
assign a25694 = ~a25692 & ~a25690;
assign a25696 = ~a25694 & a25350;
assign a25698 = ~a25466 & ~a25460;
assign a25700 = a25466 & a25460;
assign a25702 = ~a25700 & ~a25698;
assign a25704 = ~a25702 & a25386;
assign a25706 = ~a25386 & l1072;
assign a25708 = ~a25706 & ~a25704;
assign a25710 = ~a25708 & ~a25350;
assign a25712 = ~a25710 & ~a25696;
assign a25714 = ~a25712 & ~a17272;
assign a25716 = ~a25714 & ~a25688;
assign a25718 = a25716 & ~a6286;
assign a25720 = ~a25718 & ~a25680;
assign a25722 = ~a25716 & a6286;
assign a25724 = ~a25722 & ~a25720;
assign a25726 = ~a25330 & ~a25324;
assign a25728 = a25330 & a25324;
assign a25730 = ~a25728 & ~a25726;
assign a25732 = ~a25730 & a17272;
assign a25734 = ~a25372 & ~a22416;
assign a25736 = a25372 & a22416;
assign a25738 = ~a25736 & ~a25734;
assign a25740 = ~a25738 & a25350;
assign a25742 = ~a25474 & ~a25468;
assign a25744 = a25474 & a25468;
assign a25746 = ~a25744 & ~a25742;
assign a25748 = ~a25746 & a25386;
assign a25750 = ~a25386 & l1076;
assign a25752 = ~a25750 & ~a25748;
assign a25754 = ~a25752 & ~a25350;
assign a25756 = ~a25754 & ~a25740;
assign a25758 = ~a25756 & ~a17272;
assign a25760 = ~a25758 & ~a25732;
assign a25762 = a25760 & l1054;
assign a25764 = ~a25762 & ~a25724;
assign a25766 = ~a25760 & ~l1054;
assign a25768 = ~a25766 & ~a25764;
assign a25770 = ~a25338 & ~a25332;
assign a25772 = a25338 & a25332;
assign a25774 = ~a25772 & ~a25770;
assign a25776 = ~a25774 & a17272;
assign a25778 = ~a25374 & ~a22550;
assign a25780 = a25374 & a22550;
assign a25782 = ~a25780 & ~a25778;
assign a25784 = ~a25782 & a25350;
assign a25786 = ~a25482 & ~a25476;
assign a25788 = a25482 & a25476;
assign a25790 = ~a25788 & ~a25786;
assign a25792 = ~a25790 & a25386;
assign a25794 = ~a25386 & l1028;
assign a25796 = ~a25794 & ~a25792;
assign a25798 = ~a25796 & ~a25350;
assign a25800 = ~a25798 & ~a25784;
assign a25802 = ~a25800 & ~a17272;
assign a25804 = ~a25802 & ~a25776;
assign a25806 = a25804 & l1058;
assign a25808 = ~a25806 & ~a25768;
assign a25810 = ~a25804 & ~l1058;
assign a25812 = ~a25810 & ~a25808;
assign a25814 = a25812 & a25510;
assign a25816 = ~a25812 & ~a25510;
assign a25818 = ~a25816 & ~a25814;
assign a25820 = a16252 & ~l910;
assign a25822 = a25820 & a14378;
assign a25824 = a25822 & i250;
assign a25826 = ~a25824 & a16208;
assign a25828 = ~a25826 & a16220;
assign a25830 = ~a16208 & l990;
assign a25832 = a16208 & ~l990;
assign a25834 = ~a25832 & ~a25830;
assign a25836 = ~a25834 & ~a16220;
assign a25840 = a25832 & ~l986;
assign a25842 = ~a25832 & l986;
assign a25844 = ~a25842 & ~a25840;
assign a25848 = ~a25840 & ~a16214;
assign a25854 = ~a5408 & l994;
assign a25856 = ~a21594 & l996;
assign a25858 = a21594 & ~l996;
assign a25860 = ~a25858 & ~a25856;
assign a25862 = a21644 & ~a16236;
assign a25864 = a21642 & ~a16594;
assign a25866 = ~a25864 & ~a25862;
assign a25868 = ~a21642 & a16594;
assign a25870 = ~a25868 & ~a25866;
assign a25872 = a21634 & ~a16698;
assign a25874 = ~a25872 & ~a25870;
assign a25876 = ~a21634 & a16698;
assign a25878 = ~a25876 & ~a25874;
assign a25880 = a21626 & ~a16802;
assign a25882 = ~a25880 & ~a25878;
assign a25884 = ~a21626 & a16802;
assign a25886 = ~a25884 & ~a25882;
assign a25888 = a21618 & ~a16906;
assign a25890 = ~a25888 & ~a25886;
assign a25892 = ~a21618 & a16906;
assign a25894 = ~a25892 & ~a25890;
assign a25896 = a21610 & l1136;
assign a25898 = ~a25896 & ~a25894;
assign a25900 = ~a21610 & ~l1136;
assign a25902 = ~a25900 & ~a25898;
assign a25904 = a21602 & l1144;
assign a25906 = ~a25904 & ~a25902;
assign a25908 = ~a21602 & ~l1144;
assign a25910 = ~a25908 & ~a25906;
assign a25912 = ~a25910 & ~a25860;
assign a25914 = a25910 & a25860;
assign a25916 = ~a25914 & ~a25912;
assign a25918 = ~a25916 & l1100;
assign a25920 = ~a9044 & a9038;
assign a25922 = a25920 & a16188;
assign a25924 = ~a25922 & ~a14362;
assign a25926 = a25924 & a5562;
assign a25928 = a25926 & ~l946;
assign a25930 = ~a21594 & l994;
assign a25932 = a21594 & ~l994;
assign a25934 = ~a25932 & ~a25930;
assign a25936 = a21644 & ~a14354;
assign a25938 = a21642 & ~a14340;
assign a25940 = ~a25938 & ~a25936;
assign a25942 = ~a21642 & a14340;
assign a25944 = ~a25942 & ~a25940;
assign a25946 = a21634 & ~a14326;
assign a25948 = ~a25946 & ~a25944;
assign a25950 = ~a21634 & a14326;
assign a25952 = ~a25950 & ~a25948;
assign a25954 = a21626 & ~a14312;
assign a25956 = ~a25954 & ~a25952;
assign a25958 = ~a21626 & a14312;
assign a25960 = ~a25958 & ~a25956;
assign a25962 = a21618 & ~a14298;
assign a25964 = ~a25962 & ~a25960;
assign a25966 = ~a21618 & a14298;
assign a25968 = ~a25966 & ~a25964;
assign a25970 = a21610 & l1134;
assign a25972 = ~a25970 & ~a25968;
assign a25974 = ~a21610 & ~l1134;
assign a25976 = ~a25974 & ~a25972;
assign a25978 = a21602 & l1142;
assign a25980 = ~a25978 & ~a25976;
assign a25982 = ~a21602 & ~l1142;
assign a25984 = ~a25982 & ~a25980;
assign a25986 = ~a25984 & ~a25934;
assign a25988 = a25984 & a25934;
assign a25990 = ~a25988 & ~a25986;
assign a25992 = ~a25990 & ~a25928;
assign a25994 = ~a21594 & l992;
assign a25996 = a21594 & ~l992;
assign a25998 = ~a25996 & ~a25994;
assign a26000 = a21644 & ~a10646;
assign a26002 = a21642 & ~a10622;
assign a26004 = ~a26002 & ~a26000;
assign a26006 = ~a21642 & a10622;
assign a26008 = ~a26006 & ~a26004;
assign a26010 = a21634 & ~a10586;
assign a26012 = ~a26010 & ~a26008;
assign a26014 = ~a21634 & a10586;
assign a26016 = ~a26014 & ~a26012;
assign a26018 = a21626 & ~a10550;
assign a26020 = ~a26018 & ~a26016;
assign a26022 = ~a21626 & a10550;
assign a26024 = ~a26022 & ~a26020;
assign a26026 = a21618 & ~a10514;
assign a26028 = ~a26026 & ~a26024;
assign a26030 = ~a21618 & a10514;
assign a26032 = ~a26030 & ~a26028;
assign a26034 = a21610 & ~a10478;
assign a26036 = ~a26034 & ~a26032;
assign a26038 = ~a21610 & a10478;
assign a26040 = ~a26038 & ~a26036;
assign a26042 = a21602 & l1140;
assign a26044 = ~a26042 & ~a26040;
assign a26046 = ~a21602 & ~l1140;
assign a26048 = ~a26046 & ~a26044;
assign a26050 = ~a26048 & ~a25998;
assign a26052 = a26048 & a25998;
assign a26054 = ~a26052 & ~a26050;
assign a26056 = ~a26054 & a14378;
assign a26058 = ~a14378 & l992;
assign a26060 = ~a26058 & ~a26056;
assign a26062 = ~a26060 & a25928;
assign a26064 = ~a26062 & ~a25992;
assign a26066 = ~a26064 & ~l1100;
assign a26068 = ~a26066 & ~a25918;
assign a26070 = ~a26068 & a5408;
assign a26072 = ~a26070 & ~a25854;
assign a26074 = a25828 & l992;
assign a26076 = ~a25828 & l996;
assign a26078 = ~a26076 & ~a26074;
assign a26080 = ~a22670 & a22544;
assign a26082 = ~a26080 & ~a22928;
assign a26084 = a26080 & a22928;
assign a26086 = ~a26084 & ~a26082;
assign a26088 = ~a26086 & ~a12380;
assign a26090 = a23720 & ~a13958;
assign a26092 = ~a26090 & l998;
assign a26094 = a26090 & ~l998;
assign a26096 = ~a26094 & ~a26092;
assign a26098 = ~a26096 & ~a23678;
assign a26100 = a23678 & l998;
assign a26102 = ~a26100 & ~a26098;
assign a26104 = ~a26102 & a12380;
assign a26106 = ~a26104 & ~a26088;
assign a26108 = ~a8870 & l946;
assign a26110 = ~a11996 & a8970;
assign a26112 = a11996 & ~a8970;
assign a26114 = ~a11974 & a9006;
assign a26116 = a11974 & ~a9006;
assign a26118 = a8946 & l1308;
assign a26120 = ~a8946 & ~l1308;
assign a26122 = a8906 & l1000;
assign a26124 = ~a8906 & ~l1000;
assign a26126 = ~a11996 & a8954;
assign a26128 = a11996 & ~a8954;
assign a26130 = ~a11974 & a8986;
assign a26132 = a11974 & ~a8986;
assign a26134 = a8924 & l1308;
assign a26136 = ~a8924 & ~l1308;
assign a26138 = a8870 & l1000;
assign a26140 = ~a8870 & ~l1000;
assign a26142 = ~a26140 & ~a26138;
assign a26144 = a26142 & ~a26136;
assign a26146 = a26144 & ~a26134;
assign a26148 = a26146 & ~a26132;
assign a26150 = a26148 & ~a26130;
assign a26152 = a26150 & ~a26128;
assign a26154 = a26152 & ~a26126;
assign a26156 = a26154 & ~a26124;
assign a26158 = a26156 & ~a26122;
assign a26160 = a26158 & ~a26120;
assign a26162 = a26160 & ~a26118;
assign a26164 = a26162 & ~a26116;
assign a26166 = a26164 & ~a26114;
assign a26168 = a26166 & ~a26112;
assign a26170 = a26168 & ~a26110;
assign a26172 = a26106 & l1060;
assign a26174 = ~a26106 & ~l1060;
assign a26176 = ~a26174 & ~a26172;
assign a26178 = a21872 & ~a21862;
assign a26180 = ~a21872 & a21862;
assign a26182 = ~a26180 & ~a26178;
assign a26184 = ~a26182 & ~a12380;
assign a26186 = a21872 & a12836;
assign a26188 = ~a21872 & ~a12836;
assign a26190 = ~a26188 & ~a26186;
assign a26192 = ~a26190 & ~a23678;
assign a26194 = a23678 & a12836;
assign a26196 = ~a26194 & ~a26192;
assign a26198 = ~a26196 & a12380;
assign a26200 = ~a26198 & ~a26184;
assign a26202 = ~a26200 & ~l972;
assign a26204 = ~a22000 & i348;
assign a26206 = a22000 & ~i348;
assign a26208 = ~a26206 & ~a26204;
assign a26210 = ~a26208 & ~a21874;
assign a26212 = a26208 & a21874;
assign a26214 = ~a26212 & ~a26210;
assign a26216 = ~a26214 & ~a12380;
assign a26218 = a13020 & i348;
assign a26220 = ~a13020 & ~i348;
assign a26222 = ~a26220 & ~a26218;
assign a26224 = ~a26222 & ~a23680;
assign a26226 = a26222 & a23680;
assign a26228 = ~a26226 & ~a26224;
assign a26230 = ~a26228 & ~a23678;
assign a26232 = a23678 & a13020;
assign a26234 = ~a26232 & ~a26230;
assign a26236 = ~a26234 & a12380;
assign a26238 = ~a26236 & ~a26216;
assign a26240 = ~a26238 & ~l1024;
assign a26242 = ~a26240 & ~a26202;
assign a26244 = a26238 & l1024;
assign a26246 = ~a26244 & ~a26242;
assign a26248 = ~a22134 & i350;
assign a26250 = a22134 & ~i350;
assign a26252 = ~a26250 & ~a26248;
assign a26254 = ~a26252 & ~a22008;
assign a26256 = a26252 & a22008;
assign a26258 = ~a26256 & ~a26254;
assign a26260 = ~a26258 & ~a12380;
assign a26262 = a13210 & i350;
assign a26264 = ~a13210 & ~i350;
assign a26266 = ~a26264 & ~a26262;
assign a26268 = ~a26266 & ~a23688;
assign a26270 = a26266 & a23688;
assign a26272 = ~a26270 & ~a26268;
assign a26274 = ~a26272 & ~a23678;
assign a26276 = a23678 & a13210;
assign a26278 = ~a26276 & ~a26274;
assign a26280 = ~a26278 & a12380;
assign a26282 = ~a26280 & ~a26260;
assign a26284 = ~a26282 & ~l1092;
assign a26286 = ~a26284 & ~a26246;
assign a26288 = a26282 & l1092;
assign a26290 = ~a26288 & ~a26286;
assign a26292 = ~a22268 & i352;
assign a26294 = a22268 & ~i352;
assign a26296 = ~a26294 & ~a26292;
assign a26298 = ~a26296 & ~a22142;
assign a26300 = a26296 & a22142;
assign a26302 = ~a26300 & ~a26298;
assign a26304 = ~a26302 & ~a12380;
assign a26306 = a13400 & i352;
assign a26308 = ~a13400 & ~i352;
assign a26310 = ~a26308 & ~a26306;
assign a26312 = ~a26310 & ~a23696;
assign a26314 = a26310 & a23696;
assign a26316 = ~a26314 & ~a26312;
assign a26318 = ~a26316 & ~a23678;
assign a26320 = a23678 & a13400;
assign a26322 = ~a26320 & ~a26318;
assign a26324 = ~a26322 & a12380;
assign a26326 = ~a26324 & ~a26304;
assign a26328 = ~a26326 & ~l1090;
assign a26330 = ~a26328 & ~a26290;
assign a26332 = a26326 & l1090;
assign a26334 = ~a26332 & ~a26330;
assign a26336 = ~a22402 & i356;
assign a26338 = a22402 & ~i356;
assign a26340 = ~a26338 & ~a26336;
assign a26342 = ~a26340 & ~a22276;
assign a26344 = a26340 & a22276;
assign a26346 = ~a26344 & ~a26342;
assign a26348 = ~a26346 & ~a12380;
assign a26350 = a13590 & i356;
assign a26352 = ~a13590 & ~i356;
assign a26354 = ~a26352 & ~a26350;
assign a26356 = ~a26354 & ~a23704;
assign a26358 = a26354 & a23704;
assign a26360 = ~a26358 & ~a26356;
assign a26362 = ~a26360 & ~a23678;
assign a26364 = a23678 & a13590;
assign a26366 = ~a26364 & ~a26362;
assign a26368 = ~a26366 & a12380;
assign a26370 = ~a26368 & ~a26348;
assign a26372 = ~a26370 & ~l1088;
assign a26374 = ~a26372 & ~a26334;
assign a26376 = a26370 & l1088;
assign a26378 = ~a26376 & ~a26374;
assign a26380 = ~a22536 & ~i354;
assign a26382 = a22536 & i354;
assign a26384 = ~a26382 & ~a26380;
assign a26386 = ~a26384 & ~a22410;
assign a26388 = a26384 & a22410;
assign a26390 = ~a26388 & ~a26386;
assign a26392 = ~a26390 & ~a12380;
assign a26394 = a13780 & ~i354;
assign a26396 = ~a13780 & i354;
assign a26398 = ~a26396 & ~a26394;
assign a26400 = ~a26398 & ~a23712;
assign a26402 = a26398 & a23712;
assign a26404 = ~a26402 & ~a26400;
assign a26406 = ~a26404 & ~a23678;
assign a26408 = a23678 & a13780;
assign a26410 = ~a26408 & ~a26406;
assign a26412 = ~a26410 & a12380;
assign a26414 = ~a26412 & ~a26392;
assign a26416 = ~a26414 & ~l1086;
assign a26418 = ~a26416 & ~a26378;
assign a26420 = a26414 & l1086;
assign a26422 = ~a26420 & ~a26418;
assign a26424 = ~a23736 & ~l1084;
assign a26426 = ~a26424 & ~a26422;
assign a26428 = a23736 & l1084;
assign a26430 = ~a26428 & ~a26426;
assign a26432 = a26430 & ~a26176;
assign a26434 = ~a26430 & a26176;
assign a26436 = a26200 & ~a21862;
assign a26438 = a26238 & ~a22000;
assign a26440 = ~a26438 & ~a26436;
assign a26442 = ~a26238 & a22000;
assign a26444 = ~a26442 & ~a26440;
assign a26446 = a26282 & ~a22134;
assign a26448 = ~a26446 & ~a26444;
assign a26450 = ~a26282 & a22134;
assign a26452 = ~a26450 & ~a26448;
assign a26454 = a26326 & ~a22268;
assign a26456 = ~a26454 & ~a26452;
assign a26458 = ~a26326 & a22268;
assign a26460 = ~a26458 & ~a26456;
assign a26462 = a26370 & ~a22402;
assign a26464 = ~a26462 & ~a26460;
assign a26466 = ~a26370 & a22402;
assign a26468 = ~a26466 & ~a26464;
assign a26470 = a26414 & ~a22536;
assign a26472 = ~a26470 & ~a26468;
assign a26474 = ~a26414 & a22536;
assign a26476 = ~a26474 & ~a26472;
assign a26478 = a23736 & ~a22670;
assign a26480 = ~a26478 & ~a26476;
assign a26482 = ~a23736 & a22670;
assign a26484 = ~a26482 & ~a26480;
assign a26486 = a26106 & ~a22928;
assign a26488 = ~a26106 & a22928;
assign a26490 = ~a26488 & ~a26486;
assign a26492 = a26490 & ~a26484;
assign a26494 = a26200 & ~a23114;
assign a26496 = a26238 & ~a23182;
assign a26498 = ~a26496 & ~a26494;
assign a26500 = ~a26238 & a23182;
assign a26502 = ~a26500 & ~a26498;
assign a26504 = a26282 & ~a23256;
assign a26506 = ~a26504 & ~a26502;
assign a26508 = ~a26282 & a23256;
assign a26510 = ~a26508 & ~a26506;
assign a26512 = a26326 & ~a23330;
assign a26514 = ~a26512 & ~a26510;
assign a26516 = ~a26326 & a23330;
assign a26518 = ~a26516 & ~a26514;
assign a26520 = a26370 & ~a23404;
assign a26522 = ~a26520 & ~a26518;
assign a26524 = ~a26370 & a23404;
assign a26526 = ~a26524 & ~a26522;
assign a26528 = a26414 & ~a23478;
assign a26530 = ~a26528 & ~a26526;
assign a26532 = ~a26414 & a23478;
assign a26534 = ~a26532 & ~a26530;
assign a26536 = a23736 & ~a23552;
assign a26538 = ~a26536 & ~a26534;
assign a26540 = ~a23736 & a23552;
assign a26542 = ~a26540 & ~a26538;
assign a26544 = a26542 & a23632;
assign a26546 = a26544 & a26492;
assign a26548 = a26106 & ~a23626;
assign a26550 = ~a26106 & a23626;
assign a26552 = ~a26550 & ~a26548;
assign a26554 = a26552 & a26542;
assign a26556 = ~a26554 & ~a26492;
assign a26558 = ~a26556 & ~a23632;
assign a26560 = ~a26558 & ~a26546;
assign a26562 = ~a26560 & ~a26434;
assign a26564 = a26562 & ~a26432;
assign a26566 = ~a26564 & ~a22966;
assign a26568 = a26566 & a12380;
assign a26570 = a26568 & ~a26170;
assign a26572 = a26570 & ~a23030;
assign a26574 = a26572 & i336;
assign a26576 = a26574 & ~a23040;
assign a26578 = a26570 & a23030;
assign a26580 = a26578 & i372;
assign a26582 = ~a26580 & ~a26574;
assign a26584 = a26582 & l1000;
assign a26586 = ~a26584 & ~a26576;
assign a26588 = ~a26586 & ~l946;
assign a26590 = ~a26588 & ~a26108;
assign a26592 = ~a26590 & ~l886;
assign a26594 = ~a26592 & ~a5626;
assign a26596 = a2752 & a2516;
assign a26598 = a26596 & a2536;
assign a26600 = a26598 & a2504;
assign a26602 = ~a2516 & ~a2504;
assign a26604 = ~a26602 & ~a26600;
assign a26606 = ~a26604 & l1010;
assign a26608 = a2780 & ~l1010;
assign a26610 = a26608 & ~a2516;
assign a26612 = ~a26610 & ~a26606;
assign a26614 = a2536 & l1932;
assign a26616 = a26614 & ~a2504;
assign a26618 = a26616 & a26596;
assign a26620 = a26600 & l1936;
assign a26622 = ~a26620 & ~a26618;
assign a26624 = ~a2752 & a2504;
assign a26626 = a2536 & a2516;
assign a26628 = a26626 & l1938;
assign a26630 = a26628 & a26624;
assign a26632 = ~a26630 & a26622;
assign a26634 = a26626 & l1940;
assign a26636 = a26634 & ~a2504;
assign a26638 = a26636 & ~a2752;
assign a26640 = ~a26638 & a26632;
assign a26642 = a2752 & ~a2536;
assign a26644 = a26642 & a2504;
assign a26646 = a26644 & l1942;
assign a26648 = ~a26646 & a26640;
assign a26650 = a2752 & ~a2504;
assign a26652 = a2516 & l1944;
assign a26654 = a26652 & ~a2536;
assign a26656 = a26654 & a26650;
assign a26658 = ~a26656 & a26648;
assign a26660 = ~a2536 & a2516;
assign a26662 = a26660 & l1946;
assign a26664 = a26662 & ~a2752;
assign a26666 = a26664 & a2504;
assign a26668 = ~a26666 & a26658;
assign a26670 = a26660 & l1948;
assign a26672 = a26670 & ~a2752;
assign a26674 = a26672 & ~a2504;
assign a26676 = ~a26674 & a26668;
assign a26678 = a2536 & ~a2516;
assign a26680 = a26678 & l1950;
assign a26682 = a26680 & a2504;
assign a26684 = ~a26682 & a26676;
assign a26686 = a26602 & a2536;
assign a26688 = a26686 & l1952;
assign a26690 = ~a26688 & a26684;
assign a26692 = ~a26690 & a26608;
assign a26694 = a26628 & ~a2504;
assign a26696 = a26694 & a2752;
assign a26698 = a26600 & l1932;
assign a26700 = ~a26698 & ~a26696;
assign a26702 = a26634 & a26624;
assign a26704 = ~a26702 & a26700;
assign a26706 = ~a2752 & a2536;
assign a26708 = a2516 & l1942;
assign a26710 = a26708 & ~a2504;
assign a26712 = a26710 & a26706;
assign a26714 = ~a26712 & a26704;
assign a26716 = a26644 & l1944;
assign a26718 = ~a26716 & a26714;
assign a26720 = a26662 & a26650;
assign a26722 = ~a26720 & a26718;
assign a26724 = a26672 & a2504;
assign a26726 = ~a26724 & a26722;
assign a26728 = ~a2752 & ~a2536;
assign a26730 = a26728 & a2516;
assign a26732 = a26730 & l1950;
assign a26734 = a26732 & ~a2504;
assign a26736 = ~a26734 & a26726;
assign a26738 = ~a2516 & a2504;
assign a26740 = a26738 & a2536;
assign a26742 = a26740 & l1952;
assign a26744 = ~a26742 & a26736;
assign a26746 = a2536 & l1936;
assign a26748 = a26746 & ~a2516;
assign a26750 = a26748 & ~a2504;
assign a26752 = ~a26750 & a26744;
assign a26754 = ~a26752 & ~a2780;
assign a26756 = ~a26754 & ~a26692;
assign a26758 = a26650 & a2516;
assign a26760 = a26758 & a26746;
assign a26762 = a26600 & l1952;
assign a26764 = ~a26762 & ~a26760;
assign a26766 = ~a2752 & a2516;
assign a26768 = a26766 & a2504;
assign a26770 = a26768 & a26614;
assign a26772 = ~a26770 & a26764;
assign a26774 = a26694 & ~a2752;
assign a26776 = ~a26774 & a26772;
assign a26778 = a26644 & l1940;
assign a26780 = ~a26778 & a26776;
assign a26782 = a26710 & a26642;
assign a26784 = ~a26782 & a26780;
assign a26786 = a26654 & a26624;
assign a26788 = ~a26786 & a26784;
assign a26790 = a26664 & ~a2504;
assign a26792 = ~a26790 & a26788;
assign a26794 = a26740 & l1948;
assign a26796 = ~a26794 & a26792;
assign a26798 = a26680 & ~a2504;
assign a26800 = ~a26798 & a26796;
assign a26802 = ~a26800 & l1010;
assign a26804 = ~a26802 & a26756;
assign a26806 = a26804 & ~a19408;
assign a26808 = ~a26804 & a19408;
assign a26810 = ~a26808 & ~a26806;
assign a26812 = ~a18856 & a2536;
assign a26814 = a26812 & ~a2504;
assign a26816 = a26814 & a26596;
assign a26818 = a26600 & l1784;
assign a26820 = ~a26818 & ~a26816;
assign a26822 = a26626 & ~a18872;
assign a26824 = a26822 & a26624;
assign a26826 = ~a26824 & a26820;
assign a26828 = a26626 & l1786;
assign a26830 = a26828 & ~a2504;
assign a26832 = a26830 & ~a2752;
assign a26834 = ~a26832 & a26826;
assign a26836 = a26644 & l1788;
assign a26838 = ~a26836 & a26834;
assign a26840 = a2516 & l1790;
assign a26842 = a26840 & ~a2536;
assign a26844 = a26842 & a26650;
assign a26846 = ~a26844 & a26838;
assign a26848 = a26660 & l1792;
assign a26850 = a26848 & ~a2752;
assign a26852 = a26850 & a2504;
assign a26854 = ~a26852 & a26846;
assign a26856 = a26660 & l1794;
assign a26858 = a26856 & ~a2752;
assign a26860 = a26858 & ~a2504;
assign a26862 = ~a26860 & a26854;
assign a26864 = a26678 & l1796;
assign a26866 = a26864 & a2504;
assign a26868 = ~a26866 & a26862;
assign a26870 = a26686 & l1798;
assign a26872 = ~a26870 & a26868;
assign a26874 = ~a26872 & a26608;
assign a26876 = a26822 & ~a2504;
assign a26878 = a26876 & a2752;
assign a26880 = a26600 & ~a18856;
assign a26882 = ~a26880 & ~a26878;
assign a26884 = a26828 & a26624;
assign a26886 = ~a26884 & a26882;
assign a26888 = a2516 & l1788;
assign a26890 = a26888 & ~a2504;
assign a26892 = a26890 & a26706;
assign a26894 = ~a26892 & a26886;
assign a26896 = a26644 & l1790;
assign a26898 = ~a26896 & a26894;
assign a26900 = a26848 & a26650;
assign a26902 = ~a26900 & a26898;
assign a26904 = a26858 & a2504;
assign a26906 = ~a26904 & a26902;
assign a26908 = a26730 & l1796;
assign a26910 = a26908 & ~a2504;
assign a26912 = ~a26910 & a26906;
assign a26914 = a26740 & l1798;
assign a26916 = ~a26914 & a26912;
assign a26918 = a2536 & l1784;
assign a26920 = a26918 & ~a2516;
assign a26922 = a26920 & ~a2504;
assign a26924 = ~a26922 & a26916;
assign a26926 = ~a26924 & ~a2780;
assign a26928 = ~a26926 & ~a26874;
assign a26930 = a26918 & a26758;
assign a26932 = a26600 & l1798;
assign a26934 = ~a26932 & ~a26930;
assign a26936 = a26812 & a26768;
assign a26938 = ~a26936 & a26934;
assign a26940 = a26876 & ~a2752;
assign a26942 = ~a26940 & a26938;
assign a26944 = a26644 & l1786;
assign a26946 = ~a26944 & a26942;
assign a26948 = a26890 & a26642;
assign a26950 = ~a26948 & a26946;
assign a26952 = a26842 & a26624;
assign a26954 = ~a26952 & a26950;
assign a26956 = a26850 & ~a2504;
assign a26958 = ~a26956 & a26954;
assign a26960 = a26740 & l1794;
assign a26962 = ~a26960 & a26958;
assign a26964 = a26864 & ~a2504;
assign a26966 = ~a26964 & a26962;
assign a26968 = ~a26966 & l1010;
assign a26970 = ~a26968 & a26928;
assign a26972 = ~a26970 & a18850;
assign a26974 = ~a18930 & a2536;
assign a26976 = a26974 & ~a2504;
assign a26978 = a26976 & a26596;
assign a26980 = a26600 & l1804;
assign a26982 = ~a26980 & ~a26978;
assign a26984 = a26626 & ~a18946;
assign a26986 = a26984 & a26624;
assign a26988 = ~a26986 & a26982;
assign a26990 = a26626 & l1808;
assign a26992 = a26990 & ~a2504;
assign a26994 = a26992 & ~a2752;
assign a26996 = ~a26994 & a26988;
assign a26998 = a26644 & l1810;
assign a27000 = ~a26998 & a26996;
assign a27002 = a2516 & l1812;
assign a27004 = a27002 & ~a2536;
assign a27006 = a27004 & a26650;
assign a27008 = ~a27006 & a27000;
assign a27010 = a26660 & l1814;
assign a27012 = a27010 & ~a2752;
assign a27014 = a27012 & a2504;
assign a27016 = ~a27014 & a27008;
assign a27018 = a26660 & l1816;
assign a27020 = a27018 & ~a2752;
assign a27022 = a27020 & ~a2504;
assign a27024 = ~a27022 & a27016;
assign a27026 = a26678 & l1818;
assign a27028 = a27026 & a2504;
assign a27030 = ~a27028 & a27024;
assign a27032 = a26686 & l1820;
assign a27034 = ~a27032 & a27030;
assign a27036 = ~a27034 & a26608;
assign a27038 = a26984 & ~a2504;
assign a27040 = a27038 & a2752;
assign a27042 = a26600 & ~a18930;
assign a27044 = ~a27042 & ~a27040;
assign a27046 = a26990 & a26624;
assign a27048 = ~a27046 & a27044;
assign a27050 = a2516 & l1810;
assign a27052 = a27050 & ~a2504;
assign a27054 = a27052 & a26706;
assign a27056 = ~a27054 & a27048;
assign a27058 = a26644 & l1812;
assign a27060 = ~a27058 & a27056;
assign a27062 = a27010 & a26650;
assign a27064 = ~a27062 & a27060;
assign a27066 = a27020 & a2504;
assign a27068 = ~a27066 & a27064;
assign a27070 = a26730 & l1818;
assign a27072 = a27070 & ~a2504;
assign a27074 = ~a27072 & a27068;
assign a27076 = a26740 & l1820;
assign a27078 = ~a27076 & a27074;
assign a27080 = a2536 & l1804;
assign a27082 = a27080 & ~a2516;
assign a27084 = a27082 & ~a2504;
assign a27086 = ~a27084 & a27078;
assign a27088 = ~a27086 & ~a2780;
assign a27090 = ~a27088 & ~a27036;
assign a27092 = a27080 & a26758;
assign a27094 = a26600 & l1820;
assign a27096 = ~a27094 & ~a27092;
assign a27098 = a26974 & a26768;
assign a27100 = ~a27098 & a27096;
assign a27102 = a27038 & ~a2752;
assign a27104 = ~a27102 & a27100;
assign a27106 = a26644 & l1808;
assign a27108 = ~a27106 & a27104;
assign a27110 = a27052 & a26642;
assign a27112 = ~a27110 & a27108;
assign a27114 = a27004 & a26624;
assign a27116 = ~a27114 & a27112;
assign a27118 = a27012 & ~a2504;
assign a27120 = ~a27118 & a27116;
assign a27122 = a26740 & l1816;
assign a27124 = ~a27122 & a27120;
assign a27126 = a27026 & ~a2504;
assign a27128 = ~a27126 & a27124;
assign a27130 = ~a27128 & l1010;
assign a27132 = ~a27130 & a27090;
assign a27134 = ~a27132 & a18924;
assign a27136 = ~a27134 & ~a26972;
assign a27138 = a27132 & ~a18924;
assign a27140 = ~a27138 & ~a27136;
assign a27142 = ~a19010 & a2536;
assign a27144 = a27142 & ~a2504;
assign a27146 = a27144 & a26596;
assign a27148 = a26600 & l1826;
assign a27150 = ~a27148 & ~a27146;
assign a27152 = a26626 & ~a19026;
assign a27154 = a27152 & a26624;
assign a27156 = ~a27154 & a27150;
assign a27158 = a26626 & l1830;
assign a27160 = a27158 & ~a2504;
assign a27162 = a27160 & ~a2752;
assign a27164 = ~a27162 & a27156;
assign a27166 = a26644 & l1832;
assign a27168 = ~a27166 & a27164;
assign a27170 = a2516 & l1834;
assign a27172 = a27170 & ~a2536;
assign a27174 = a27172 & a26650;
assign a27176 = ~a27174 & a27168;
assign a27178 = a26660 & l1836;
assign a27180 = a27178 & ~a2752;
assign a27182 = a27180 & a2504;
assign a27184 = ~a27182 & a27176;
assign a27186 = a26660 & l1838;
assign a27188 = a27186 & ~a2752;
assign a27190 = a27188 & ~a2504;
assign a27192 = ~a27190 & a27184;
assign a27194 = a26678 & l1840;
assign a27196 = a27194 & a2504;
assign a27198 = ~a27196 & a27192;
assign a27200 = a26678 & l1842;
assign a27202 = a27200 & ~a2504;
assign a27204 = ~a27202 & a27198;
assign a27206 = ~a27204 & a26608;
assign a27208 = a27152 & ~a2504;
assign a27210 = a27208 & a2752;
assign a27212 = a26600 & ~a19010;
assign a27214 = ~a27212 & ~a27210;
assign a27216 = a27158 & a26624;
assign a27218 = ~a27216 & a27214;
assign a27220 = a2516 & l1832;
assign a27222 = a27220 & ~a2504;
assign a27224 = a27222 & a26706;
assign a27226 = ~a27224 & a27218;
assign a27228 = a26644 & l1834;
assign a27230 = ~a27228 & a27226;
assign a27232 = a27178 & a26650;
assign a27234 = ~a27232 & a27230;
assign a27236 = a27188 & a2504;
assign a27238 = ~a27236 & a27234;
assign a27240 = a26730 & l1840;
assign a27242 = a27240 & ~a2504;
assign a27244 = ~a27242 & a27238;
assign a27246 = a27200 & a2504;
assign a27248 = ~a27246 & a27244;
assign a27250 = a2536 & l1826;
assign a27252 = a27250 & ~a2516;
assign a27254 = a27252 & ~a2504;
assign a27256 = ~a27254 & a27248;
assign a27258 = ~a27256 & ~a2780;
assign a27260 = ~a27258 & ~a27206;
assign a27262 = a27250 & a26758;
assign a27264 = a26600 & l1842;
assign a27266 = ~a27264 & ~a27262;
assign a27268 = a27142 & a26768;
assign a27270 = ~a27268 & a27266;
assign a27272 = a27208 & ~a2752;
assign a27274 = ~a27272 & a27270;
assign a27276 = a26644 & l1830;
assign a27278 = ~a27276 & a27274;
assign a27280 = a27222 & a26642;
assign a27282 = ~a27280 & a27278;
assign a27284 = a27172 & a26624;
assign a27286 = ~a27284 & a27282;
assign a27288 = a27180 & ~a2504;
assign a27290 = ~a27288 & a27286;
assign a27292 = a26740 & l1838;
assign a27294 = ~a27292 & a27290;
assign a27296 = a27194 & ~a2504;
assign a27298 = ~a27296 & a27294;
assign a27300 = ~a27298 & l1010;
assign a27302 = ~a27300 & a27260;
assign a27304 = ~a27302 & a19004;
assign a27306 = ~a27304 & ~a27140;
assign a27308 = a27302 & ~a19004;
assign a27310 = ~a27308 & ~a27306;
assign a27312 = ~a19092 & a2536;
assign a27314 = a27312 & ~a2504;
assign a27316 = a27314 & a26596;
assign a27318 = a26600 & l1848;
assign a27320 = ~a27318 & ~a27316;
assign a27322 = a26626 & ~a19108;
assign a27324 = a27322 & a26624;
assign a27326 = ~a27324 & a27320;
assign a27328 = a26626 & l1852;
assign a27330 = a27328 & ~a2504;
assign a27332 = a27330 & ~a2752;
assign a27334 = ~a27332 & a27326;
assign a27336 = a26644 & l1854;
assign a27338 = ~a27336 & a27334;
assign a27340 = a2516 & l1856;
assign a27342 = a27340 & ~a2536;
assign a27344 = a27342 & a26650;
assign a27346 = ~a27344 & a27338;
assign a27348 = a26660 & l1858;
assign a27350 = a27348 & ~a2752;
assign a27352 = a27350 & a2504;
assign a27354 = ~a27352 & a27346;
assign a27356 = a26660 & l1860;
assign a27358 = a27356 & ~a2752;
assign a27360 = a27358 & ~a2504;
assign a27362 = ~a27360 & a27354;
assign a27364 = a26678 & l1862;
assign a27366 = a27364 & a2504;
assign a27368 = ~a27366 & a27362;
assign a27370 = a26678 & l1864;
assign a27372 = a27370 & ~a2504;
assign a27374 = ~a27372 & a27368;
assign a27376 = ~a27374 & a26608;
assign a27378 = a27322 & ~a2504;
assign a27380 = a27378 & a2752;
assign a27382 = a26600 & ~a19092;
assign a27384 = ~a27382 & ~a27380;
assign a27386 = a27328 & a26624;
assign a27388 = ~a27386 & a27384;
assign a27390 = a2516 & l1854;
assign a27392 = a27390 & ~a2504;
assign a27394 = a27392 & a26706;
assign a27396 = ~a27394 & a27388;
assign a27398 = a26644 & l1856;
assign a27400 = ~a27398 & a27396;
assign a27402 = a27348 & a26650;
assign a27404 = ~a27402 & a27400;
assign a27406 = a27358 & a2504;
assign a27408 = ~a27406 & a27404;
assign a27410 = a26730 & l1862;
assign a27412 = a27410 & ~a2504;
assign a27414 = ~a27412 & a27408;
assign a27416 = a27370 & a2504;
assign a27418 = ~a27416 & a27414;
assign a27420 = a2536 & l1848;
assign a27422 = a27420 & ~a2516;
assign a27424 = a27422 & ~a2504;
assign a27426 = ~a27424 & a27418;
assign a27428 = ~a27426 & ~a2780;
assign a27430 = ~a27428 & ~a27376;
assign a27432 = a27420 & a26758;
assign a27434 = a26600 & l1864;
assign a27436 = ~a27434 & ~a27432;
assign a27438 = a27312 & a26768;
assign a27440 = ~a27438 & a27436;
assign a27442 = a27378 & ~a2752;
assign a27444 = ~a27442 & a27440;
assign a27446 = a26644 & l1852;
assign a27448 = ~a27446 & a27444;
assign a27450 = a27392 & a26642;
assign a27452 = ~a27450 & a27448;
assign a27454 = a27342 & a26624;
assign a27456 = ~a27454 & a27452;
assign a27458 = a27350 & ~a2504;
assign a27460 = ~a27458 & a27456;
assign a27462 = a26740 & l1860;
assign a27464 = ~a27462 & a27460;
assign a27466 = a27364 & ~a2504;
assign a27468 = ~a27466 & a27464;
assign a27470 = ~a27468 & l1010;
assign a27472 = ~a27470 & a27430;
assign a27474 = ~a27472 & a19086;
assign a27476 = ~a27474 & ~a27310;
assign a27478 = a27472 & ~a19086;
assign a27480 = ~a27478 & ~a27476;
assign a27482 = ~a19174 & a2536;
assign a27484 = a27482 & ~a2504;
assign a27486 = a27484 & a26596;
assign a27488 = a26600 & l1870;
assign a27490 = ~a27488 & ~a27486;
assign a27492 = a26626 & ~a19190;
assign a27494 = a27492 & a26624;
assign a27496 = ~a27494 & a27490;
assign a27498 = a26626 & l1874;
assign a27500 = a27498 & ~a2504;
assign a27502 = a27500 & ~a2752;
assign a27504 = ~a27502 & a27496;
assign a27506 = a26644 & l1876;
assign a27508 = ~a27506 & a27504;
assign a27510 = a2516 & l1878;
assign a27512 = a27510 & ~a2536;
assign a27514 = a27512 & a26650;
assign a27516 = ~a27514 & a27508;
assign a27518 = a26660 & l1880;
assign a27520 = a27518 & ~a2752;
assign a27522 = a27520 & a2504;
assign a27524 = ~a27522 & a27516;
assign a27526 = a26660 & l1882;
assign a27528 = a27526 & ~a2752;
assign a27530 = a27528 & ~a2504;
assign a27532 = ~a27530 & a27524;
assign a27534 = a26678 & l1884;
assign a27536 = a27534 & a2504;
assign a27538 = ~a27536 & a27532;
assign a27540 = a26678 & l1886;
assign a27542 = a27540 & ~a2504;
assign a27544 = ~a27542 & a27538;
assign a27546 = ~a27544 & a26608;
assign a27548 = a27492 & ~a2504;
assign a27550 = a27548 & a2752;
assign a27552 = a26600 & ~a19174;
assign a27554 = ~a27552 & ~a27550;
assign a27556 = a27498 & a26624;
assign a27558 = ~a27556 & a27554;
assign a27560 = a2516 & l1876;
assign a27562 = a27560 & ~a2504;
assign a27564 = a27562 & a26706;
assign a27566 = ~a27564 & a27558;
assign a27568 = a26644 & l1878;
assign a27570 = ~a27568 & a27566;
assign a27572 = a27518 & a26650;
assign a27574 = ~a27572 & a27570;
assign a27576 = a27528 & a2504;
assign a27578 = ~a27576 & a27574;
assign a27580 = a26730 & l1884;
assign a27582 = a27580 & ~a2504;
assign a27584 = ~a27582 & a27578;
assign a27586 = a27540 & a2504;
assign a27588 = ~a27586 & a27584;
assign a27590 = a2536 & l1870;
assign a27592 = a27590 & ~a2516;
assign a27594 = a27592 & ~a2504;
assign a27596 = ~a27594 & a27588;
assign a27598 = ~a27596 & ~a2780;
assign a27600 = ~a27598 & ~a27546;
assign a27602 = a27590 & a26758;
assign a27604 = a26600 & l1886;
assign a27606 = ~a27604 & ~a27602;
assign a27608 = a27482 & a26768;
assign a27610 = ~a27608 & a27606;
assign a27612 = a27548 & ~a2752;
assign a27614 = ~a27612 & a27610;
assign a27616 = a26644 & l1874;
assign a27618 = ~a27616 & a27614;
assign a27620 = a27562 & a26642;
assign a27622 = ~a27620 & a27618;
assign a27624 = a27512 & a26624;
assign a27626 = ~a27624 & a27622;
assign a27628 = a27520 & ~a2504;
assign a27630 = ~a27628 & a27626;
assign a27632 = a26740 & l1882;
assign a27634 = ~a27632 & a27630;
assign a27636 = a27534 & ~a2504;
assign a27638 = ~a27636 & a27634;
assign a27640 = ~a27638 & l1010;
assign a27642 = ~a27640 & a27600;
assign a27644 = ~a27642 & a19168;
assign a27646 = ~a27644 & ~a27480;
assign a27648 = a27642 & ~a19168;
assign a27650 = ~a27648 & ~a27646;
assign a27652 = ~a19256 & a2536;
assign a27654 = a27652 & ~a2504;
assign a27656 = a27654 & a26596;
assign a27658 = a26600 & l1892;
assign a27660 = ~a27658 & ~a27656;
assign a27662 = a26626 & ~a19272;
assign a27664 = a27662 & a26624;
assign a27666 = ~a27664 & a27660;
assign a27668 = a26626 & l1896;
assign a27670 = a27668 & ~a2504;
assign a27672 = a27670 & ~a2752;
assign a27674 = ~a27672 & a27666;
assign a27676 = a26644 & l1898;
assign a27678 = ~a27676 & a27674;
assign a27680 = a2516 & l1900;
assign a27682 = a27680 & ~a2536;
assign a27684 = a27682 & a26650;
assign a27686 = ~a27684 & a27678;
assign a27688 = a26660 & l1902;
assign a27690 = a27688 & ~a2752;
assign a27692 = a27690 & a2504;
assign a27694 = ~a27692 & a27686;
assign a27696 = a26660 & l1904;
assign a27698 = a27696 & ~a2752;
assign a27700 = a27698 & ~a2504;
assign a27702 = ~a27700 & a27694;
assign a27704 = a26678 & l1906;
assign a27706 = a27704 & a2504;
assign a27708 = ~a27706 & a27702;
assign a27710 = a26678 & l1908;
assign a27712 = a27710 & ~a2504;
assign a27714 = ~a27712 & a27708;
assign a27716 = ~a27714 & a26608;
assign a27718 = a27662 & ~a2504;
assign a27720 = a27718 & a2752;
assign a27722 = a26600 & ~a19256;
assign a27724 = ~a27722 & ~a27720;
assign a27726 = a27668 & a26624;
assign a27728 = ~a27726 & a27724;
assign a27730 = a2516 & l1898;
assign a27732 = a27730 & ~a2504;
assign a27734 = a27732 & a26706;
assign a27736 = ~a27734 & a27728;
assign a27738 = a26644 & l1900;
assign a27740 = ~a27738 & a27736;
assign a27742 = a27688 & a26650;
assign a27744 = ~a27742 & a27740;
assign a27746 = a27698 & a2504;
assign a27748 = ~a27746 & a27744;
assign a27750 = a26730 & l1906;
assign a27752 = a27750 & ~a2504;
assign a27754 = ~a27752 & a27748;
assign a27756 = a27710 & a2504;
assign a27758 = ~a27756 & a27754;
assign a27760 = a2536 & l1892;
assign a27762 = a27760 & ~a2516;
assign a27764 = a27762 & ~a2504;
assign a27766 = ~a27764 & a27758;
assign a27768 = ~a27766 & ~a2780;
assign a27770 = ~a27768 & ~a27716;
assign a27772 = a27760 & a26758;
assign a27774 = a26600 & l1908;
assign a27776 = ~a27774 & ~a27772;
assign a27778 = a27652 & a26768;
assign a27780 = ~a27778 & a27776;
assign a27782 = a27718 & ~a2752;
assign a27784 = ~a27782 & a27780;
assign a27786 = a26644 & l1896;
assign a27788 = ~a27786 & a27784;
assign a27790 = a27732 & a26642;
assign a27792 = ~a27790 & a27788;
assign a27794 = a27682 & a26624;
assign a27796 = ~a27794 & a27792;
assign a27798 = a27690 & ~a2504;
assign a27800 = ~a27798 & a27796;
assign a27802 = a26740 & l1904;
assign a27804 = ~a27802 & a27800;
assign a27806 = a27704 & ~a2504;
assign a27808 = ~a27806 & a27804;
assign a27810 = ~a27808 & l1010;
assign a27812 = ~a27810 & a27770;
assign a27814 = ~a27812 & a19250;
assign a27816 = ~a27814 & ~a27650;
assign a27818 = a27812 & ~a19250;
assign a27820 = ~a27818 & ~a27816;
assign a27822 = a2536 & l1910;
assign a27824 = a27822 & ~a2504;
assign a27826 = a27824 & a26596;
assign a27828 = a26600 & l1914;
assign a27830 = ~a27828 & ~a27826;
assign a27832 = a26626 & ~a19348;
assign a27834 = a27832 & a26624;
assign a27836 = ~a27834 & a27830;
assign a27838 = a26626 & l1918;
assign a27840 = a27838 & ~a2504;
assign a27842 = a27840 & ~a2752;
assign a27844 = ~a27842 & a27836;
assign a27846 = a26644 & l1920;
assign a27848 = ~a27846 & a27844;
assign a27850 = a2516 & l1922;
assign a27852 = a27850 & ~a2536;
assign a27854 = a27852 & a26650;
assign a27856 = ~a27854 & a27848;
assign a27858 = a26660 & l1924;
assign a27860 = a27858 & ~a2752;
assign a27862 = a27860 & a2504;
assign a27864 = ~a27862 & a27856;
assign a27866 = a26660 & l1926;
assign a27868 = a27866 & ~a2752;
assign a27870 = a27868 & ~a2504;
assign a27872 = ~a27870 & a27864;
assign a27874 = a26678 & l1928;
assign a27876 = a27874 & a2504;
assign a27878 = ~a27876 & a27872;
assign a27880 = a26678 & l1930;
assign a27882 = a27880 & ~a2504;
assign a27884 = ~a27882 & a27878;
assign a27886 = ~a27884 & a26608;
assign a27888 = a27832 & ~a2504;
assign a27890 = a27888 & a2752;
assign a27892 = a26600 & l1910;
assign a27894 = ~a27892 & ~a27890;
assign a27896 = a27838 & a26624;
assign a27898 = ~a27896 & a27894;
assign a27900 = a2516 & l1920;
assign a27902 = a27900 & ~a2504;
assign a27904 = a27902 & a26706;
assign a27906 = ~a27904 & a27898;
assign a27908 = a26644 & l1922;
assign a27910 = ~a27908 & a27906;
assign a27912 = a27858 & a26650;
assign a27914 = ~a27912 & a27910;
assign a27916 = a27868 & a2504;
assign a27918 = ~a27916 & a27914;
assign a27920 = a26730 & l1928;
assign a27922 = a27920 & ~a2504;
assign a27924 = ~a27922 & a27918;
assign a27926 = a27880 & a2504;
assign a27928 = ~a27926 & a27924;
assign a27930 = a2536 & l1914;
assign a27932 = a27930 & ~a2516;
assign a27934 = a27932 & ~a2504;
assign a27936 = ~a27934 & a27928;
assign a27938 = ~a27936 & ~a2780;
assign a27940 = ~a27938 & ~a27886;
assign a27942 = a27930 & a26758;
assign a27944 = a26600 & l1930;
assign a27946 = ~a27944 & ~a27942;
assign a27948 = a27822 & a26768;
assign a27950 = ~a27948 & a27946;
assign a27952 = a27888 & ~a2752;
assign a27954 = ~a27952 & a27950;
assign a27956 = a26644 & l1918;
assign a27958 = ~a27956 & a27954;
assign a27960 = a27902 & a26642;
assign a27962 = ~a27960 & a27958;
assign a27964 = a27852 & a26624;
assign a27966 = ~a27964 & a27962;
assign a27968 = a27860 & ~a2504;
assign a27970 = ~a27968 & a27966;
assign a27972 = a26740 & l1926;
assign a27974 = ~a27972 & a27970;
assign a27976 = a27874 & ~a2504;
assign a27978 = ~a27976 & a27974;
assign a27980 = ~a27978 & l1010;
assign a27982 = ~a27980 & a27940;
assign a27984 = ~a27982 & a19332;
assign a27986 = ~a27984 & ~a27820;
assign a27988 = a27982 & ~a19332;
assign a27990 = ~a27988 & ~a27986;
assign a27992 = a27990 & a26810;
assign a27994 = a26970 & ~a18850;
assign a27996 = ~a27994 & ~a27138;
assign a27998 = ~a27996 & ~a27134;
assign a28000 = ~a27998 & ~a27308;
assign a28002 = ~a28000 & ~a27304;
assign a28004 = ~a28002 & ~a27478;
assign a28006 = ~a28004 & ~a27474;
assign a28008 = ~a28006 & ~a27648;
assign a28010 = ~a28008 & ~a27644;
assign a28012 = ~a28010 & ~a27818;
assign a28014 = ~a28012 & ~a27814;
assign a28016 = ~a28014 & ~a27988;
assign a28018 = ~a27984 & ~a26810;
assign a28020 = a28018 & ~a28016;
assign a28022 = ~a28020 & ~a27992;
assign a28024 = a26626 & a18596;
assign a28026 = a28024 & ~a2504;
assign a28028 = a28026 & a2752;
assign a28030 = a26600 & a18568;
assign a28032 = ~a28030 & ~a28028;
assign a28034 = a26626 & l1974;
assign a28036 = a28034 & a26624;
assign a28038 = ~a28036 & a28032;
assign a28040 = a2516 & l1976;
assign a28042 = a28040 & ~a2504;
assign a28044 = a28042 & a26706;
assign a28046 = ~a28044 & a28038;
assign a28048 = a26644 & l1978;
assign a28050 = ~a28048 & a28046;
assign a28052 = a26660 & l1980;
assign a28054 = a28052 & a26650;
assign a28056 = ~a28054 & a28050;
assign a28058 = a26660 & l1982;
assign a28060 = a28058 & ~a2752;
assign a28062 = a28060 & a2504;
assign a28064 = ~a28062 & a28056;
assign a28066 = a26730 & a18646;
assign a28068 = a28066 & ~a2504;
assign a28070 = ~a28068 & a28064;
assign a28072 = a26678 & l1986;
assign a28074 = a28072 & a2504;
assign a28076 = ~a28074 & a28070;
assign a28078 = a18582 & a2536;
assign a28080 = a28078 & ~a2516;
assign a28082 = a28080 & ~a2504;
assign a28084 = ~a28082 & a28076;
assign a28086 = ~a28084 & ~a2780;
assign a28088 = a18568 & a2536;
assign a28090 = a28088 & ~a2504;
assign a28092 = a28090 & a26596;
assign a28094 = a26600 & a18582;
assign a28096 = ~a28094 & ~a28092;
assign a28098 = a28024 & a26624;
assign a28100 = ~a28098 & a28096;
assign a28102 = a28034 & ~a2504;
assign a28104 = a28102 & ~a2752;
assign a28106 = ~a28104 & a28100;
assign a28108 = a26644 & l1976;
assign a28110 = ~a28108 & a28106;
assign a28112 = a2516 & l1978;
assign a28114 = a28112 & ~a2536;
assign a28116 = a28114 & a26650;
assign a28118 = ~a28116 & a28110;
assign a28120 = a28052 & ~a2752;
assign a28122 = a28120 & a2504;
assign a28124 = ~a28122 & a28118;
assign a28126 = a28060 & ~a2504;
assign a28128 = ~a28126 & a28124;
assign a28130 = a26678 & a18646;
assign a28132 = a28130 & a2504;
assign a28134 = ~a28132 & a28128;
assign a28136 = a28072 & ~a2504;
assign a28138 = ~a28136 & a28134;
assign a28140 = ~a28138 & a26608;
assign a28142 = ~a28140 & ~a28086;
assign a28144 = a28078 & a26758;
assign a28146 = a26600 & l1986;
assign a28148 = ~a28146 & ~a28144;
assign a28150 = a28088 & a26768;
assign a28152 = ~a28150 & a28148;
assign a28154 = a28026 & ~a2752;
assign a28156 = ~a28154 & a28152;
assign a28158 = a26644 & l1974;
assign a28160 = ~a28158 & a28156;
assign a28162 = a28042 & a26642;
assign a28164 = ~a28162 & a28160;
assign a28166 = a28114 & a26624;
assign a28168 = ~a28166 & a28164;
assign a28170 = a28120 & ~a2504;
assign a28172 = ~a28170 & a28168;
assign a28174 = a26740 & l1982;
assign a28176 = ~a28174 & a28172;
assign a28178 = a28130 & ~a2504;
assign a28180 = ~a28178 & a28176;
assign a28182 = ~a28180 & l1010;
assign a28184 = ~a28182 & a28142;
assign a28186 = ~a28184 & ~l886;
assign a28190 = a25828 & ~a10646;
assign a28192 = ~a25828 & ~a16236;
assign a28196 = ~a14354 & ~a5408;
assign a28198 = ~a21644 & ~a16236;
assign a28200 = a21644 & a16236;
assign a28202 = ~a28200 & ~a28198;
assign a28204 = ~a28202 & l1100;
assign a28206 = ~a21644 & ~a14354;
assign a28208 = a21644 & a14354;
assign a28210 = ~a28208 & ~a28206;
assign a28212 = ~a28210 & ~a25928;
assign a28214 = ~a21644 & ~a10646;
assign a28216 = a21644 & a10646;
assign a28218 = ~a28216 & ~a28214;
assign a28220 = ~a28218 & a14378;
assign a28222 = ~a14378 & ~a10646;
assign a28224 = ~a28222 & ~a28220;
assign a28226 = ~a28224 & a25928;
assign a28228 = ~a28226 & ~a28212;
assign a28230 = ~a28228 & ~l1100;
assign a28232 = ~a28230 & ~a28204;
assign a28234 = ~a28232 & a5408;
assign a28238 = ~a5624 & l948;
assign a28240 = a28238 & a7226;
assign a28242 = ~a8430 & a8150;
assign a28244 = ~a8802 & a8434;
assign a28246 = ~a28244 & ~a28242;
assign a28248 = ~a28246 & a5568;
assign a28250 = ~a28246 & ~a5568;
assign a28252 = a28250 & a5594;
assign a28254 = ~a28252 & ~a28248;
assign a28256 = a28250 & ~a5594;
assign a28258 = a28256 & a5600;
assign a28260 = ~a28258 & a28254;
assign a28262 = a28256 & ~a5600;
assign a28264 = a28262 & a5606;
assign a28266 = ~a28264 & a28260;
assign a28268 = a28262 & ~a5606;
assign a28270 = a28268 & l960;
assign a28272 = ~a28270 & a28266;
assign a28274 = a28268 & ~l960;
assign a28276 = a28274 & l962;
assign a28278 = ~a28276 & a28272;
assign a28280 = a28274 & ~l962;
assign a28282 = a28280 & l964;
assign a28284 = ~a28282 & a28278;
assign a28286 = a28280 & ~l964;
assign a28288 = a28286 & l966;
assign a28290 = ~a28288 & a28284;
assign a28292 = a28286 & ~l966;
assign a28294 = a28292 & l968;
assign a28296 = ~a28294 & a28290;
assign a28298 = a28292 & ~l968;
assign a28300 = a28298 & l970;
assign a28302 = ~a28300 & a28296;
assign a28304 = ~a28302 & ~l886;
assign a28306 = a28304 & ~l948;
assign a28308 = a8802 & a8434;
assign a28310 = a28308 & a5568;
assign a28312 = a28308 & ~a5568;
assign a28314 = a28312 & a5594;
assign a28316 = ~a28314 & ~a28310;
assign a28318 = a28312 & ~a5594;
assign a28320 = a28318 & a5600;
assign a28322 = ~a28320 & a28316;
assign a28324 = a28318 & ~a5600;
assign a28326 = a28324 & a5606;
assign a28328 = ~a28326 & a28322;
assign a28330 = a28324 & ~a5606;
assign a28332 = a28330 & l960;
assign a28334 = ~a28332 & a28328;
assign a28336 = a28330 & ~l960;
assign a28338 = a28336 & l962;
assign a28340 = ~a28338 & a28334;
assign a28342 = a28336 & ~l962;
assign a28344 = a28342 & l964;
assign a28346 = ~a28344 & a28340;
assign a28348 = a28342 & ~l964;
assign a28350 = a28348 & l966;
assign a28352 = ~a28350 & a28346;
assign a28354 = a28348 & ~l966;
assign a28356 = a28354 & l968;
assign a28358 = ~a28356 & a28352;
assign a28360 = a28354 & ~l968;
assign a28362 = a28360 & l970;
assign a28364 = ~a28362 & a28358;
assign a28366 = ~a28364 & ~l886;
assign a28368 = a28366 & ~l948;
assign a28370 = ~a28368 & ~a28306;
assign a28372 = ~a28370 & a5748;
assign a28374 = ~a7780 & l972;
assign a28376 = ~a7858 & ~a7782;
assign a28378 = ~a28376 & ~l972;
assign a28380 = ~a28378 & ~a28374;
assign a28382 = a28380 & a28372;
assign a28384 = a28298 & ~l970;
assign a28386 = a28360 & ~l970;
assign a28388 = ~a28386 & ~a28384;
assign a28390 = ~a28388 & ~l886;
assign a28392 = a28390 & a5748;
assign a28394 = ~a6166 & l972;
assign a28396 = ~a6232 & ~a6168;
assign a28398 = ~a28396 & ~l972;
assign a28400 = ~a28398 & ~a28394;
assign a28402 = a28400 & a28392;
assign a28404 = ~a28402 & ~a28382;
assign a28406 = ~a28376 & l972;
assign a28408 = ~a7856 & ~l972;
assign a28410 = ~a28408 & ~a28406;
assign a28412 = a28410 & a28372;
assign a28414 = ~a28396 & l972;
assign a28416 = ~a6230 & ~l972;
assign a28418 = ~a28416 & ~a28414;
assign a28420 = a28418 & a28392;
assign a28422 = ~a28420 & ~a28412;
assign a28424 = a28422 & a28404;
assign a28426 = a28424 & i532;
assign a28428 = ~a28426 & a28404;
assign a28430 = a28428 & ~a5760;
assign a28432 = ~a28428 & a5760;
assign a28434 = ~a28432 & ~a28430;
assign a28436 = a28434 & a5748;
assign a28438 = ~a5760 & ~a5748;
assign a28440 = ~a28438 & ~a28436;
assign a28442 = ~a28440 & ~a28238;
assign a28444 = ~a28442 & ~a28240;
assign a28446 = ~a28444 & ~l886;
assign a28450 = ~a17436 & l1024;
assign a28452 = ~a28450 & ~a17486;
assign a28454 = a25350 & ~a21670;
assign a28456 = ~a25350 & l1032;
assign a28458 = ~a28456 & ~a28454;
assign a28460 = ~a28458 & ~a17272;
assign a28462 = ~a28460 & ~a17462;
assign a28464 = a7226 & ~a6426;
assign a28466 = ~a7226 & a6426;
assign a28468 = ~a28466 & ~a28464;
assign a28470 = ~a28468 & a28238;
assign a28472 = ~a28428 & ~a5760;
assign a28474 = ~a28428 & a28392;
assign a28476 = a28474 & l972;
assign a28478 = a28428 & a28392;
assign a28480 = a28478 & ~l972;
assign a28482 = ~a28480 & ~a28476;
assign a28484 = ~a28482 & a5760;
assign a28486 = a28478 & l972;
assign a28488 = ~a28486 & ~a28484;
assign a28490 = ~a6148 & ~a5796;
assign a28492 = ~a6134 & ~a5814;
assign a28494 = ~a6120 & ~a5832;
assign a28496 = ~a6046 & ~l1088;
assign a28498 = ~a28496 & ~a5922;
assign a28500 = ~a28498 & a5832;
assign a28502 = ~a28500 & ~a28494;
assign a28504 = ~a28502 & l1090;
assign a28506 = ~a6064 & ~l1090;
assign a28508 = ~a28506 & ~a28504;
assign a28510 = ~a28508 & a5814;
assign a28512 = ~a28510 & ~a28492;
assign a28514 = ~a28512 & l1092;
assign a28516 = ~a6082 & ~l1092;
assign a28518 = ~a28516 & ~a28514;
assign a28520 = ~a28518 & a5796;
assign a28522 = ~a28520 & ~a28490;
assign a28524 = ~a28522 & a5778;
assign a28526 = ~a28524 & ~a6154;
assign a28528 = ~a28526 & l1024;
assign a28530 = ~a6152 & ~l1024;
assign a28532 = ~a28530 & ~a28528;
assign a28534 = a28532 & ~a28488;
assign a28536 = a28474 & ~l972;
assign a28538 = ~a28482 & ~a5760;
assign a28540 = ~a28538 & ~a28536;
assign a28542 = ~a6152 & l1024;
assign a28544 = ~a6222 & ~a6160;
assign a28546 = ~a28544 & ~l1024;
assign a28548 = ~a28546 & ~a28542;
assign a28550 = a28548 & ~a28540;
assign a28552 = ~a28428 & a28372;
assign a28554 = a28552 & ~l972;
assign a28556 = a28552 & l972;
assign a28558 = a28428 & a28372;
assign a28560 = a28558 & ~l972;
assign a28562 = ~a28560 & ~a28556;
assign a28564 = ~a28562 & ~a5760;
assign a28566 = ~a28564 & ~a28554;
assign a28568 = ~a7766 & l1024;
assign a28570 = ~a7848 & ~a7774;
assign a28572 = ~a28570 & ~l1024;
assign a28574 = ~a28572 & ~a28568;
assign a28576 = a28574 & ~a28566;
assign a28578 = ~a28562 & a5760;
assign a28580 = a28558 & l972;
assign a28582 = ~a28580 & ~a28578;
assign a28584 = ~a7762 & ~a5796;
assign a28586 = ~a7748 & ~a5814;
assign a28588 = ~a7734 & ~a5832;
assign a28590 = a7720 & ~a5850;
assign a28592 = ~a7640 & a5850;
assign a28594 = ~a28592 & ~a28590;
assign a28596 = a28594 & l1088;
assign a28598 = ~a7650 & ~l1088;
assign a28600 = ~a28598 & ~a28596;
assign a28602 = ~a28600 & a5832;
assign a28604 = ~a28602 & ~a28588;
assign a28606 = ~a28604 & l1090;
assign a28608 = ~a7668 & ~l1090;
assign a28610 = ~a28608 & ~a28606;
assign a28612 = ~a28610 & a5814;
assign a28614 = ~a28612 & ~a28586;
assign a28616 = ~a28614 & l1092;
assign a28618 = ~a7686 & ~l1092;
assign a28620 = ~a28618 & ~a28616;
assign a28622 = ~a28620 & a5796;
assign a28624 = ~a28622 & ~a28584;
assign a28626 = ~a28624 & a5778;
assign a28628 = ~a28626 & ~a7768;
assign a28630 = ~a28628 & l1024;
assign a28632 = ~a7766 & ~l1024;
assign a28634 = ~a28632 & ~a28630;
assign a28636 = a28634 & ~a28582;
assign a28638 = ~a28636 & ~a28576;
assign a28640 = a28638 & ~a28550;
assign a28642 = a28640 & ~a28534;
assign a28644 = a28548 & ~a28488;
assign a28646 = ~a28544 & l1024;
assign a28648 = ~a6220 & ~l1024;
assign a28650 = ~a28648 & ~a28646;
assign a28652 = a28650 & ~a28540;
assign a28654 = ~a28570 & l1024;
assign a28656 = ~a7846 & ~l1024;
assign a28658 = ~a28656 & ~a28654;
assign a28660 = a28658 & ~a28566;
assign a28662 = ~a28582 & a28574;
assign a28664 = ~a28662 & ~a28660;
assign a28666 = a28664 & ~a28652;
assign a28668 = a28666 & ~a28644;
assign a28670 = a28668 & a28642;
assign a28672 = a28670 & i534;
assign a28674 = ~a28672 & a28642;
assign a28676 = a28674 & ~a5778;
assign a28678 = ~a28674 & a5778;
assign a28680 = ~a28678 & ~a28676;
assign a28682 = ~a28680 & ~a28472;
assign a28684 = a28680 & a28472;
assign a28686 = ~a28684 & ~a28682;
assign a28688 = ~a28686 & a28434;
assign a28690 = a28686 & ~a28434;
assign a28692 = ~a28690 & ~a28688;
assign a28694 = ~a28692 & a5748;
assign a28696 = ~a5778 & ~a5748;
assign a28698 = ~a28696 & ~a28694;
assign a28700 = ~a28698 & ~a28238;
assign a28702 = ~a28700 & ~a28470;
assign a28704 = ~a28702 & ~l886;
assign a28708 = ~a7226 & ~a6426;
assign a28710 = ~a28708 & ~a6434;
assign a28712 = a28708 & a6434;
assign a28714 = ~a28712 & ~a28710;
assign a28716 = ~a28714 & a28238;
assign a28718 = ~a28686 & ~a28434;
assign a28720 = ~a28674 & ~a5778;
assign a28722 = ~a28720 & ~a28472;
assign a28724 = a28674 & a5778;
assign a28726 = ~a28724 & ~a28722;
assign a28728 = a28674 & ~a28488;
assign a28730 = a28728 & l1024;
assign a28732 = a28730 & a5778;
assign a28734 = ~a28514 & ~a6146;
assign a28736 = ~a28734 & ~a5796;
assign a28738 = ~a28512 & a5796;
assign a28740 = ~a28738 & ~a28736;
assign a28742 = a28740 & a28732;
assign a28744 = ~a28674 & ~a28540;
assign a28746 = a28744 & l1024;
assign a28748 = a28674 & ~a28540;
assign a28750 = ~a28674 & ~a28488;
assign a28752 = ~a28750 & ~a28748;
assign a28754 = ~a28752 & ~l1024;
assign a28756 = ~a28754 & ~a28746;
assign a28758 = ~a28756 & a5778;
assign a28760 = ~a28752 & l1024;
assign a28762 = ~a28760 & ~a28758;
assign a28764 = a28728 & ~l1024;
assign a28766 = ~a28764 & a28762;
assign a28768 = a28730 & ~a5778;
assign a28770 = ~a28768 & a28766;
assign a28772 = ~a6138 & ~a5796;
assign a28774 = ~a28734 & a5796;
assign a28776 = ~a28774 & ~a28772;
assign a28778 = a28776 & ~a28770;
assign a28780 = a28744 & ~l1024;
assign a28782 = ~a28756 & ~a5778;
assign a28784 = ~a28782 & ~a28780;
assign a28786 = ~a6212 & ~a6140;
assign a28788 = ~a28786 & ~a5796;
assign a28790 = ~a6138 & a5796;
assign a28792 = ~a28790 & ~a28788;
assign a28794 = a28792 & ~a28784;
assign a28796 = a28674 & ~a28582;
assign a28798 = a28796 & l1024;
assign a28800 = a28798 & a5778;
assign a28802 = ~a28616 & ~a7760;
assign a28804 = ~a28802 & ~a5796;
assign a28806 = ~a28614 & a5796;
assign a28808 = ~a28806 & ~a28804;
assign a28810 = a28808 & a28800;
assign a28812 = ~a28674 & ~a28566;
assign a28814 = a28812 & ~l1024;
assign a28816 = a28812 & l1024;
assign a28818 = a28674 & ~a28566;
assign a28820 = ~a28674 & ~a28582;
assign a28822 = ~a28820 & ~a28818;
assign a28824 = ~a28822 & ~l1024;
assign a28826 = ~a28824 & ~a28816;
assign a28828 = ~a28826 & ~a5778;
assign a28830 = ~a28828 & ~a28814;
assign a28832 = ~a7838 & ~a7754;
assign a28834 = ~a28832 & ~a5796;
assign a28836 = ~a7752 & a5796;
assign a28838 = ~a28836 & ~a28834;
assign a28840 = a28838 & ~a28830;
assign a28842 = ~a28826 & a5778;
assign a28844 = ~a28822 & l1024;
assign a28846 = ~a28844 & ~a28842;
assign a28848 = a28796 & ~l1024;
assign a28850 = ~a28848 & a28846;
assign a28852 = a28798 & ~a5778;
assign a28854 = ~a28852 & a28850;
assign a28856 = ~a7752 & ~a5796;
assign a28858 = ~a28802 & a5796;
assign a28860 = ~a28858 & ~a28856;
assign a28862 = a28860 & ~a28854;
assign a28864 = ~a28862 & ~a28840;
assign a28866 = a28864 & ~a28810;
assign a28868 = a28866 & ~a28794;
assign a28870 = a28868 & ~a28778;
assign a28872 = a28870 & ~a28742;
assign a28874 = a28776 & a28732;
assign a28876 = a28792 & ~a28770;
assign a28878 = ~a6210 & ~a5796;
assign a28880 = ~a28786 & a5796;
assign a28882 = ~a28880 & ~a28878;
assign a28884 = a28882 & ~a28784;
assign a28886 = a28860 & a28800;
assign a28888 = ~a7836 & ~a5796;
assign a28890 = ~a28832 & a5796;
assign a28892 = ~a28890 & ~a28888;
assign a28894 = a28892 & ~a28830;
assign a28896 = ~a28854 & a28838;
assign a28898 = ~a28896 & ~a28894;
assign a28900 = a28898 & ~a28886;
assign a28902 = a28900 & ~a28884;
assign a28904 = a28902 & ~a28876;
assign a28906 = a28904 & ~a28874;
assign a28908 = a28906 & a28872;
assign a28910 = a28908 & i536;
assign a28912 = ~a28910 & a28872;
assign a28914 = a28912 & ~a5796;
assign a28916 = ~a28912 & a5796;
assign a28918 = ~a28916 & ~a28914;
assign a28920 = ~a28918 & ~a28726;
assign a28922 = a28918 & a28726;
assign a28924 = ~a28922 & ~a28920;
assign a28926 = ~a28924 & ~a28718;
assign a28928 = a28924 & a28718;
assign a28930 = ~a28928 & ~a28926;
assign a28932 = ~a28930 & a5748;
assign a28934 = ~a5796 & ~a5748;
assign a28936 = ~a28934 & ~a28932;
assign a28938 = ~a28936 & ~a28238;
assign a28940 = ~a28938 & ~a28716;
assign a28942 = ~a28940 & ~l886;
assign a28946 = a28708 & ~a6434;
assign a28948 = ~a28946 & ~a6442;
assign a28950 = a28946 & a6442;
assign a28952 = ~a28950 & ~a28948;
assign a28954 = ~a28952 & a28238;
assign a28956 = ~a28924 & a28718;
assign a28958 = ~a28912 & ~a5796;
assign a28960 = ~a28958 & ~a28726;
assign a28962 = a28912 & a5796;
assign a28964 = ~a28962 & ~a28960;
assign a28966 = a28912 & ~a28770;
assign a28968 = ~a28912 & a28732;
assign a28970 = ~a28968 & ~a28966;
assign a28972 = ~a28970 & a5796;
assign a28974 = a28912 & a28732;
assign a28976 = a28974 & ~a5796;
assign a28978 = ~a28976 & ~a28972;
assign a28980 = ~a28978 & l1092;
assign a28982 = a28974 & a5796;
assign a28984 = ~a28982 & ~a28980;
assign a28986 = ~a28504 & ~a6132;
assign a28988 = ~a28986 & ~a5814;
assign a28990 = ~a28502 & a5814;
assign a28992 = ~a28990 & ~a28988;
assign a28994 = a28992 & ~a28984;
assign a28996 = ~a28912 & ~a28784;
assign a28998 = a28996 & a5796;
assign a29000 = a28912 & ~a28784;
assign a29002 = ~a28912 & ~a28770;
assign a29004 = ~a29002 & ~a29000;
assign a29006 = ~a29004 & ~a5796;
assign a29008 = ~a29006 & ~a28998;
assign a29010 = ~a29008 & l1092;
assign a29012 = ~a29004 & a5796;
assign a29014 = ~a29012 & ~a29010;
assign a29016 = ~a28978 & ~l1092;
assign a29018 = ~a29016 & a29014;
assign a29020 = ~a28970 & ~a5796;
assign a29022 = ~a29020 & a29018;
assign a29024 = ~a6124 & ~a5814;
assign a29026 = ~a28986 & a5814;
assign a29028 = ~a29026 & ~a29024;
assign a29030 = a29028 & ~a29022;
assign a29032 = ~a29008 & ~l1092;
assign a29034 = a28996 & ~a5796;
assign a29036 = ~a29034 & ~a29032;
assign a29038 = ~a6202 & ~a6126;
assign a29040 = ~a29038 & ~a5814;
assign a29042 = ~a6124 & a5814;
assign a29044 = ~a29042 & ~a29040;
assign a29046 = a29044 & ~a29036;
assign a29048 = a28912 & ~a28854;
assign a29050 = ~a28912 & a28800;
assign a29052 = ~a29050 & ~a29048;
assign a29054 = ~a29052 & a5796;
assign a29056 = a28912 & a28800;
assign a29058 = a29056 & ~a5796;
assign a29060 = ~a29058 & ~a29054;
assign a29062 = ~a29060 & l1092;
assign a29064 = a29056 & a5796;
assign a29066 = ~a29064 & ~a29062;
assign a29068 = ~a28606 & ~a7746;
assign a29070 = ~a29068 & ~a5814;
assign a29072 = ~a28604 & a5814;
assign a29074 = ~a29072 & ~a29070;
assign a29076 = a29074 & ~a29066;
assign a29078 = ~a28912 & ~a28830;
assign a29080 = a29078 & a5796;
assign a29082 = a28912 & ~a28830;
assign a29084 = ~a28912 & ~a28854;
assign a29086 = ~a29084 & ~a29082;
assign a29088 = ~a29086 & ~a5796;
assign a29090 = ~a29088 & ~a29080;
assign a29092 = ~a29090 & ~l1092;
assign a29094 = a29078 & ~a5796;
assign a29096 = ~a29094 & ~a29092;
assign a29098 = ~a7828 & ~a7740;
assign a29100 = ~a29098 & ~a5814;
assign a29102 = ~a7738 & a5814;
assign a29104 = ~a29102 & ~a29100;
assign a29106 = a29104 & ~a29096;
assign a29108 = ~a29090 & l1092;
assign a29110 = ~a29086 & a5796;
assign a29112 = ~a29110 & ~a29108;
assign a29114 = ~a29060 & ~l1092;
assign a29116 = ~a29114 & a29112;
assign a29118 = ~a29052 & ~a5796;
assign a29120 = ~a29118 & a29116;
assign a29122 = ~a7738 & ~a5814;
assign a29124 = ~a29068 & a5814;
assign a29126 = ~a29124 & ~a29122;
assign a29128 = a29126 & ~a29120;
assign a29130 = ~a29128 & ~a29106;
assign a29132 = a29130 & ~a29076;
assign a29134 = a29132 & ~a29046;
assign a29136 = a29134 & ~a29030;
assign a29138 = a29136 & ~a28994;
assign a29140 = a29028 & ~a28984;
assign a29142 = a29044 & ~a29022;
assign a29144 = ~a6200 & ~a5814;
assign a29146 = ~a29038 & a5814;
assign a29148 = ~a29146 & ~a29144;
assign a29150 = a29148 & ~a29036;
assign a29152 = a29126 & ~a29066;
assign a29154 = ~a7826 & ~a5814;
assign a29156 = ~a29098 & a5814;
assign a29158 = ~a29156 & ~a29154;
assign a29160 = a29158 & ~a29096;
assign a29162 = ~a29120 & a29104;
assign a29164 = ~a29162 & ~a29160;
assign a29166 = a29164 & ~a29152;
assign a29168 = a29166 & ~a29150;
assign a29170 = a29168 & ~a29142;
assign a29172 = a29170 & ~a29140;
assign a29174 = a29172 & a29138;
assign a29176 = a29174 & i538;
assign a29178 = ~a29176 & a29138;
assign a29180 = a29178 & ~a5814;
assign a29182 = ~a29178 & a5814;
assign a29184 = ~a29182 & ~a29180;
assign a29186 = ~a29184 & ~a28964;
assign a29188 = a29184 & a28964;
assign a29190 = ~a29188 & ~a29186;
assign a29192 = ~a29190 & ~a28956;
assign a29194 = a29190 & a28956;
assign a29196 = ~a29194 & ~a29192;
assign a29198 = ~a29196 & a5748;
assign a29200 = ~a5814 & ~a5748;
assign a29202 = ~a29200 & ~a29198;
assign a29204 = ~a29202 & ~a28238;
assign a29206 = ~a29204 & ~a28954;
assign a29208 = ~a29206 & ~l886;
assign a29212 = a28946 & ~a6442;
assign a29214 = ~a29212 & ~a6450;
assign a29216 = a29212 & a6450;
assign a29218 = ~a29216 & ~a29214;
assign a29220 = ~a29218 & a28238;
assign a29222 = ~a29190 & a28956;
assign a29224 = ~a29178 & ~a5814;
assign a29226 = ~a29224 & ~a28964;
assign a29228 = a29178 & a5814;
assign a29230 = ~a29228 & ~a29226;
assign a29232 = a29178 & ~a29022;
assign a29234 = ~a29178 & ~a28984;
assign a29236 = ~a29234 & ~a29232;
assign a29238 = ~a29236 & a5814;
assign a29240 = a29178 & ~a28984;
assign a29242 = a29240 & ~a5814;
assign a29244 = ~a29242 & ~a29238;
assign a29246 = ~a29244 & l1090;
assign a29248 = a29240 & a5814;
assign a29250 = ~a29248 & ~a29246;
assign a29252 = ~a29250 & ~a5936;
assign a29254 = ~a29178 & ~a29036;
assign a29256 = a29254 & a5814;
assign a29258 = a29178 & ~a29036;
assign a29260 = ~a29178 & ~a29022;
assign a29262 = ~a29260 & ~a29258;
assign a29264 = ~a29262 & ~a5814;
assign a29266 = ~a29264 & ~a29256;
assign a29268 = ~a29266 & l1090;
assign a29270 = ~a29262 & a5814;
assign a29272 = ~a29270 & ~a29268;
assign a29274 = ~a29244 & ~l1090;
assign a29276 = ~a29274 & a29272;
assign a29278 = ~a29236 & ~a5814;
assign a29280 = ~a29278 & a29276;
assign a29282 = ~a29280 & a5928;
assign a29284 = ~a29266 & ~l1090;
assign a29286 = a29254 & ~a5814;
assign a29288 = ~a29286 & ~a29284;
assign a29290 = ~a6192 & ~a6114;
assign a29292 = ~a29290 & ~a5832;
assign a29294 = ~a5910 & a5832;
assign a29296 = ~a29294 & ~a29292;
assign a29298 = a29296 & ~a29288;
assign a29300 = a29178 & ~a29120;
assign a29302 = ~a29178 & ~a29066;
assign a29304 = ~a29302 & ~a29300;
assign a29306 = ~a29304 & a5814;
assign a29308 = a29178 & ~a29066;
assign a29310 = a29308 & ~a5814;
assign a29312 = ~a29310 & ~a29306;
assign a29314 = ~a29312 & l1090;
assign a29316 = a29308 & a5814;
assign a29318 = ~a29316 & ~a29314;
assign a29320 = ~a28596 & ~a7732;
assign a29322 = a29320 & ~a5832;
assign a29324 = ~a28594 & a5832;
assign a29326 = ~a29324 & ~a29322;
assign a29328 = ~a29326 & ~a29318;
assign a29330 = ~a29178 & ~a29096;
assign a29332 = a29330 & a5814;
assign a29334 = a29178 & ~a29096;
assign a29336 = ~a29178 & ~a29120;
assign a29338 = ~a29336 & ~a29334;
assign a29340 = ~a29338 & ~a5814;
assign a29342 = ~a29340 & ~a29332;
assign a29344 = ~a29342 & ~l1090;
assign a29346 = a29330 & ~a5814;
assign a29348 = ~a29346 & ~a29344;
assign a29350 = ~a7818 & ~a7726;
assign a29352 = ~a29350 & ~a5832;
assign a29354 = ~a7724 & a5832;
assign a29356 = ~a29354 & ~a29352;
assign a29358 = a29356 & ~a29348;
assign a29360 = ~a29342 & l1090;
assign a29362 = ~a29338 & a5814;
assign a29364 = ~a29362 & ~a29360;
assign a29366 = ~a29312 & ~l1090;
assign a29368 = ~a29366 & a29364;
assign a29370 = ~a29304 & ~a5814;
assign a29372 = ~a29370 & a29368;
assign a29374 = ~a7724 & ~a5832;
assign a29376 = ~a29320 & a5832;
assign a29378 = ~a29376 & ~a29374;
assign a29380 = a29378 & ~a29372;
assign a29382 = ~a29380 & ~a29358;
assign a29384 = a29382 & ~a29328;
assign a29386 = a29384 & ~a29298;
assign a29388 = a29386 & ~a29282;
assign a29390 = a29388 & ~a29252;
assign a29392 = ~a29250 & a5928;
assign a29394 = a29296 & ~a29280;
assign a29396 = ~a6190 & ~a5832;
assign a29398 = ~a29290 & a5832;
assign a29400 = ~a29398 & ~a29396;
assign a29402 = a29400 & ~a29288;
assign a29404 = a29378 & ~a29318;
assign a29406 = ~a7816 & ~a5832;
assign a29408 = ~a29350 & a5832;
assign a29410 = ~a29408 & ~a29406;
assign a29412 = a29410 & ~a29348;
assign a29414 = ~a29372 & a29356;
assign a29416 = ~a29414 & ~a29412;
assign a29418 = a29416 & ~a29404;
assign a29420 = a29418 & ~a29402;
assign a29422 = a29420 & ~a29394;
assign a29424 = a29422 & ~a29392;
assign a29426 = a29424 & a29390;
assign a29428 = a29426 & i540;
assign a29430 = ~a29428 & a29390;
assign a29432 = a29430 & ~a5832;
assign a29434 = ~a29430 & a5832;
assign a29436 = ~a29434 & ~a29432;
assign a29438 = ~a29436 & ~a29230;
assign a29440 = a29436 & a29230;
assign a29442 = ~a29440 & ~a29438;
assign a29444 = ~a29442 & ~a29222;
assign a29446 = a29442 & a29222;
assign a29448 = ~a29446 & ~a29444;
assign a29450 = ~a29448 & a5748;
assign a29452 = ~a5832 & ~a5748;
assign a29454 = ~a29452 & ~a29450;
assign a29456 = ~a29454 & ~a28238;
assign a29458 = ~a29456 & ~a29220;
assign a29460 = ~a29458 & ~l886;
assign a29464 = a29212 & ~a6450;
assign a29466 = ~a29464 & l1130;
assign a29468 = a29464 & ~l1130;
assign a29470 = ~a29468 & ~a29466;
assign a29472 = ~a29470 & a28238;
assign a29474 = ~a29442 & a29222;
assign a29476 = ~a29430 & ~a5832;
assign a29478 = ~a29476 & ~a29230;
assign a29480 = a29430 & a5832;
assign a29482 = ~a29480 & ~a29478;
assign a29484 = ~a29482 & ~a5850;
assign a29486 = a29482 & a5850;
assign a29488 = ~a29486 & ~a29484;
assign a29490 = ~a29488 & ~a29474;
assign a29492 = a29488 & a29474;
assign a29494 = ~a29492 & ~a29490;
assign a29496 = ~a29494 & a5748;
assign a29498 = ~a5850 & ~a5748;
assign a29500 = ~a29498 & ~a29496;
assign a29502 = ~a29500 & ~a28238;
assign a29504 = ~a29502 & ~a29472;
assign a29506 = ~a29504 & ~l886;
assign a29510 = a29464 & l1130;
assign a29512 = ~a29510 & l1138;
assign a29514 = a29510 & ~l1138;
assign a29516 = ~a29514 & ~a29512;
assign a29518 = ~a29516 & a28238;
assign a29520 = ~a29488 & a29474;
assign a29522 = a29482 & ~a5850;
assign a29524 = ~a29522 & ~a5868;
assign a29526 = a29522 & a5868;
assign a29528 = ~a29526 & ~a29524;
assign a29530 = ~a29528 & ~a29520;
assign a29532 = a29528 & a29520;
assign a29534 = ~a29532 & ~a29530;
assign a29536 = ~a29534 & a5748;
assign a29538 = ~a5868 & ~a5748;
assign a29540 = ~a29538 & ~a29536;
assign a29542 = ~a29540 & ~a28238;
assign a29544 = ~a29542 & ~a29518;
assign a29546 = ~a29544 & ~l886;
assign a29550 = ~a17436 & l1060;
assign a29552 = ~a29550 & ~a17444;
assign a29554 = a25350 & ~a21880;
assign a29556 = ~a25350 & l1064;
assign a29558 = ~a29556 & ~a29554;
assign a29560 = ~a29558 & ~a17272;
assign a29562 = ~a29560 & ~a17480;
assign a29564 = a25350 & ~a22014;
assign a29566 = ~a25350 & l1066;
assign a29568 = ~a29566 & ~a29564;
assign a29570 = ~a29568 & ~a17272;
assign a29572 = ~a29570 & ~a17504;
assign a29574 = a25350 & ~a22148;
assign a29576 = ~a25350 & l1070;
assign a29578 = ~a29576 & ~a29574;
assign a29580 = ~a29578 & ~a17272;
assign a29582 = ~a29580 & ~a17528;
assign a29584 = a25350 & ~a22282;
assign a29586 = ~a25350 & l1074;
assign a29588 = ~a29586 & ~a29584;
assign a29590 = ~a29588 & ~a17272;
assign a29592 = ~a29590 & ~a17552;
assign a29594 = a25350 & ~a22416;
assign a29596 = ~a25350 & l1078;
assign a29598 = ~a29596 & ~a29594;
assign a29600 = ~a29598 & ~a17272;
assign a29602 = ~a29600 & ~a17576;
assign a29604 = a29510 & l1138;
assign a29606 = ~a29604 & l1082;
assign a29608 = a29604 & ~l1082;
assign a29610 = ~a29608 & ~a29606;
assign a29612 = ~a29610 & a28238;
assign a29614 = a29522 & ~a5868;
assign a29616 = ~a29614 & ~a5874;
assign a29618 = a29614 & a5874;
assign a29620 = ~a29618 & ~a29616;
assign a29622 = ~a29528 & a29520;
assign a29624 = ~a29622 & ~a29620;
assign a29626 = a29622 & a29620;
assign a29628 = ~a29626 & ~a29624;
assign a29630 = ~a29628 & a5748;
assign a29632 = ~a5874 & ~a5748;
assign a29634 = ~a29632 & ~a29630;
assign a29636 = ~a29634 & ~a28238;
assign a29638 = ~a29636 & ~a29612;
assign a29640 = ~a29638 & ~l886;
assign a29644 = ~a17436 & l1084;
assign a29646 = ~a29644 & ~a17608;
assign a29648 = ~a17436 & l1086;
assign a29650 = ~a29648 & ~a17582;
assign a29652 = ~a17436 & l1088;
assign a29654 = ~a29652 & ~a17558;
assign a29656 = ~a17436 & l1090;
assign a29658 = ~a29656 & ~a17534;
assign a29660 = ~a17436 & l1092;
assign a29662 = ~a29660 & ~a17510;
assign a29664 = ~a14340 & ~a5408;
assign a29666 = ~a21642 & ~a16594;
assign a29668 = a21642 & a16594;
assign a29670 = ~a29668 & ~a29666;
assign a29672 = ~a29670 & ~a25862;
assign a29674 = a29670 & a25862;
assign a29676 = ~a29674 & ~a29672;
assign a29678 = ~a29676 & l1100;
assign a29680 = ~a21642 & ~a14340;
assign a29682 = a21642 & a14340;
assign a29684 = ~a29682 & ~a29680;
assign a29686 = ~a29684 & ~a25936;
assign a29688 = a29684 & a25936;
assign a29690 = ~a29688 & ~a29686;
assign a29692 = ~a29690 & ~a25928;
assign a29694 = ~a21642 & ~a10622;
assign a29696 = a21642 & a10622;
assign a29698 = ~a29696 & ~a29694;
assign a29700 = ~a29698 & ~a26000;
assign a29702 = a29698 & a26000;
assign a29704 = ~a29702 & ~a29700;
assign a29706 = ~a29704 & a14378;
assign a29708 = ~a14378 & ~a10622;
assign a29710 = ~a29708 & ~a29706;
assign a29712 = ~a29710 & a25928;
assign a29714 = ~a29712 & ~a29692;
assign a29716 = ~a29714 & ~l1100;
assign a29718 = ~a29716 & ~a29678;
assign a29720 = ~a29718 & a5408;
assign a29724 = a25828 & ~a10622;
assign a29726 = ~a25828 & ~a16594;
assign a29730 = ~a14326 & ~a5408;
assign a29732 = ~a21634 & ~a16698;
assign a29734 = a21634 & a16698;
assign a29736 = ~a29734 & ~a29732;
assign a29738 = ~a29736 & ~a25870;
assign a29740 = a29736 & a25870;
assign a29742 = ~a29740 & ~a29738;
assign a29744 = ~a29742 & l1100;
assign a29746 = ~a21634 & ~a14326;
assign a29748 = a21634 & a14326;
assign a29750 = ~a29748 & ~a29746;
assign a29752 = ~a29750 & ~a25944;
assign a29754 = a29750 & a25944;
assign a29756 = ~a29754 & ~a29752;
assign a29758 = ~a29756 & ~a25928;
assign a29760 = ~a21634 & ~a10586;
assign a29762 = a21634 & a10586;
assign a29764 = ~a29762 & ~a29760;
assign a29766 = ~a29764 & ~a26008;
assign a29768 = a29764 & a26008;
assign a29770 = ~a29768 & ~a29766;
assign a29772 = ~a29770 & a14378;
assign a29774 = ~a14378 & ~a10586;
assign a29776 = ~a29774 & ~a29772;
assign a29778 = ~a29776 & a25928;
assign a29780 = ~a29778 & ~a29758;
assign a29782 = ~a29780 & ~l1100;
assign a29784 = ~a29782 & ~a29744;
assign a29786 = ~a29784 & a5408;
assign a29790 = a25828 & ~a10586;
assign a29792 = ~a25828 & ~a16698;
assign a29796 = ~a14312 & ~a5408;
assign a29798 = ~a21626 & ~a16802;
assign a29800 = a21626 & a16802;
assign a29802 = ~a29800 & ~a29798;
assign a29804 = ~a29802 & ~a25878;
assign a29806 = a29802 & a25878;
assign a29808 = ~a29806 & ~a29804;
assign a29810 = ~a29808 & l1100;
assign a29812 = ~a21626 & ~a14312;
assign a29814 = a21626 & a14312;
assign a29816 = ~a29814 & ~a29812;
assign a29818 = ~a29816 & ~a25952;
assign a29820 = a29816 & a25952;
assign a29822 = ~a29820 & ~a29818;
assign a29824 = ~a29822 & ~a25928;
assign a29826 = ~a21626 & ~a10550;
assign a29828 = a21626 & a10550;
assign a29830 = ~a29828 & ~a29826;
assign a29832 = ~a29830 & ~a26016;
assign a29834 = a29830 & a26016;
assign a29836 = ~a29834 & ~a29832;
assign a29838 = ~a29836 & a14378;
assign a29840 = ~a14378 & ~a10550;
assign a29842 = ~a29840 & ~a29838;
assign a29844 = ~a29842 & a25928;
assign a29846 = ~a29844 & ~a29824;
assign a29848 = ~a29846 & ~l1100;
assign a29850 = ~a29848 & ~a29810;
assign a29852 = ~a29850 & a5408;
assign a29856 = a25828 & ~a10550;
assign a29858 = ~a25828 & ~a16802;
assign a29862 = ~a14298 & ~a5408;
assign a29864 = ~a21618 & ~a16906;
assign a29866 = a21618 & a16906;
assign a29868 = ~a29866 & ~a29864;
assign a29870 = ~a29868 & ~a25886;
assign a29872 = a29868 & a25886;
assign a29874 = ~a29872 & ~a29870;
assign a29876 = ~a29874 & l1100;
assign a29878 = ~a21618 & ~a14298;
assign a29880 = a21618 & a14298;
assign a29882 = ~a29880 & ~a29878;
assign a29884 = ~a29882 & ~a25960;
assign a29886 = a29882 & a25960;
assign a29888 = ~a29886 & ~a29884;
assign a29890 = ~a29888 & ~a25928;
assign a29892 = ~a21618 & ~a10514;
assign a29894 = a21618 & a10514;
assign a29896 = ~a29894 & ~a29892;
assign a29898 = ~a29896 & ~a26024;
assign a29900 = a29896 & a26024;
assign a29902 = ~a29900 & ~a29898;
assign a29904 = ~a29902 & a14378;
assign a29906 = ~a14378 & ~a10514;
assign a29908 = ~a29906 & ~a29904;
assign a29910 = ~a29908 & a25928;
assign a29912 = ~a29910 & ~a29890;
assign a29914 = ~a29912 & ~l1100;
assign a29916 = ~a29914 & ~a29876;
assign a29918 = ~a29916 & a5408;
assign a29922 = a25828 & ~a10514;
assign a29924 = ~a25828 & ~a16906;
assign a29928 = ~a5408 & l1134;
assign a29930 = ~a21610 & l1136;
assign a29932 = a21610 & ~l1136;
assign a29934 = ~a29932 & ~a29930;
assign a29936 = ~a29934 & ~a25894;
assign a29938 = a29934 & a25894;
assign a29940 = ~a29938 & ~a29936;
assign a29942 = ~a29940 & l1100;
assign a29944 = ~a21610 & l1134;
assign a29946 = a21610 & ~l1134;
assign a29948 = ~a29946 & ~a29944;
assign a29950 = ~a29948 & ~a25968;
assign a29952 = a29948 & a25968;
assign a29954 = ~a29952 & ~a29950;
assign a29956 = ~a29954 & ~a25928;
assign a29958 = ~a21610 & ~a10478;
assign a29960 = a21610 & a10478;
assign a29962 = ~a29960 & ~a29958;
assign a29964 = ~a29962 & ~a26032;
assign a29966 = a29962 & a26032;
assign a29968 = ~a29966 & ~a29964;
assign a29970 = ~a29968 & a14378;
assign a29972 = ~a14378 & ~a10478;
assign a29974 = ~a29972 & ~a29970;
assign a29976 = ~a29974 & a25928;
assign a29978 = ~a29976 & ~a29956;
assign a29980 = ~a29978 & ~l1100;
assign a29982 = ~a29980 & ~a29942;
assign a29984 = ~a29982 & a5408;
assign a29988 = a25828 & ~a10478;
assign a29990 = ~a25828 & l1136;
assign a29992 = ~a29990 & ~a29988;
assign a29994 = ~a5408 & l1142;
assign a29996 = ~a21602 & l1144;
assign a29998 = a21602 & ~l1144;
assign a30000 = ~a29998 & ~a29996;
assign a30002 = ~a30000 & ~a25902;
assign a30004 = a30000 & a25902;
assign a30006 = ~a30004 & ~a30002;
assign a30008 = ~a30006 & l1100;
assign a30010 = ~a21602 & l1142;
assign a30012 = a21602 & ~l1142;
assign a30014 = ~a30012 & ~a30010;
assign a30016 = ~a30014 & ~a25976;
assign a30018 = a30014 & a25976;
assign a30020 = ~a30018 & ~a30016;
assign a30022 = ~a30020 & ~a25928;
assign a30024 = ~a21602 & l1140;
assign a30026 = a21602 & ~l1140;
assign a30028 = ~a30026 & ~a30024;
assign a30030 = ~a30028 & ~a26040;
assign a30032 = a30028 & a26040;
assign a30034 = ~a30032 & ~a30030;
assign a30036 = ~a30034 & a14378;
assign a30038 = ~a14378 & l1140;
assign a30040 = ~a30038 & ~a30036;
assign a30042 = ~a30040 & a25928;
assign a30044 = ~a30042 & ~a30022;
assign a30046 = ~a30044 & ~l1100;
assign a30048 = ~a30046 & ~a30008;
assign a30050 = ~a30048 & a5408;
assign a30052 = ~a30050 & ~a29994;
assign a30054 = a25828 & l1140;
assign a30056 = ~a25828 & l1144;
assign a30058 = ~a30056 & ~a30054;
assign a30060 = l884 & ~l880;
assign a30062 = ~l1150 & ~l884;
assign a30064 = a30062 & l1148;
assign a30066 = l1150 & ~l884;
assign a30068 = a30066 & ~l1148;
assign a30070 = ~a30068 & ~a30064;
assign a30072 = a30070 & ~a30060;
assign a30074 = ~a18872 & a6538;
assign a30076 = a30074 & l1148;
assign a30078 = ~a18856 & ~l1166;
assign a30080 = a19864 & ~l1148;
assign a30082 = a30080 & a30078;
assign a30084 = ~a30082 & ~a30076;
assign a30086 = l1162 & ~l1148;
assign a30088 = l1786 & ~l1166;
assign a30090 = a30088 & a30086;
assign a30092 = ~a30090 & a30084;
assign a30094 = l1162 & l1148;
assign a30096 = a30094 & ~l1166;
assign a30098 = a30096 & l1788;
assign a30100 = ~a30098 & a30092;
assign a30102 = l1166 & ~l1162;
assign a30104 = a30102 & ~l1148;
assign a30106 = a30104 & l1790;
assign a30108 = ~a30106 & a30100;
assign a30110 = a30102 & l1792;
assign a30112 = a30110 & l1148;
assign a30114 = ~a30112 & a30108;
assign a30116 = l1166 & ~l1148;
assign a30118 = ~l1164 & l1162;
assign a30120 = a30118 & a30116;
assign a30122 = a30120 & l1794;
assign a30124 = ~a30122 & a30114;
assign a30126 = a6522 & l1796;
assign a30128 = a30126 & l1148;
assign a30130 = ~a30128 & a30124;
assign a30132 = l1164 & ~l1148;
assign a30134 = a30132 & l1798;
assign a30136 = ~a30134 & a30130;
assign a30138 = l1164 & l1148;
assign a30140 = a30138 & ~l1166;
assign a30142 = a30140 & l1784;
assign a30144 = ~a30142 & a30136;
assign a30146 = ~a30144 & ~l1150;
assign a30148 = a19864 & l1148;
assign a30150 = a30148 & a30088;
assign a30152 = a30074 & ~l1148;
assign a30154 = ~a30152 & ~a30150;
assign a30156 = a30086 & ~l1166;
assign a30158 = a30156 & l1788;
assign a30160 = ~a30158 & a30154;
assign a30162 = a30096 & l1790;
assign a30164 = ~a30162 & a30160;
assign a30166 = a30110 & ~l1148;
assign a30168 = ~a30166 & a30164;
assign a30170 = a30102 & l1148;
assign a30172 = a30170 & l1794;
assign a30174 = ~a30172 & a30168;
assign a30176 = a30126 & ~l1148;
assign a30178 = ~a30176 & a30174;
assign a30180 = a30094 & l1166;
assign a30182 = a30180 & ~l1164;
assign a30184 = a30182 & l1798;
assign a30186 = ~a30184 & a30178;
assign a30188 = a30132 & l1784;
assign a30190 = ~a30188 & a30186;
assign a30192 = a30138 & a30078;
assign a30194 = ~a30192 & a30190;
assign a30196 = ~a30194 & l1150;
assign a30198 = ~a30196 & ~a30146;
assign a30200 = a30198 & ~a17476;
assign a30202 = ~a18946 & a6538;
assign a30204 = a30202 & l1148;
assign a30206 = ~a18930 & ~l1166;
assign a30208 = a30206 & a30080;
assign a30210 = ~a30208 & ~a30204;
assign a30212 = l1808 & ~l1166;
assign a30214 = a30212 & a30086;
assign a30216 = ~a30214 & a30210;
assign a30218 = a30096 & l1810;
assign a30220 = ~a30218 & a30216;
assign a30222 = a30104 & l1812;
assign a30224 = ~a30222 & a30220;
assign a30226 = a30102 & l1814;
assign a30228 = a30226 & l1148;
assign a30230 = ~a30228 & a30224;
assign a30232 = a30120 & l1816;
assign a30234 = ~a30232 & a30230;
assign a30236 = a6522 & l1818;
assign a30238 = a30236 & l1148;
assign a30240 = ~a30238 & a30234;
assign a30242 = a30132 & l1820;
assign a30244 = ~a30242 & a30240;
assign a30246 = a30140 & l1804;
assign a30248 = ~a30246 & a30244;
assign a30250 = ~a30248 & ~l1150;
assign a30252 = a30212 & a30148;
assign a30254 = a30202 & ~l1148;
assign a30256 = ~a30254 & ~a30252;
assign a30258 = a30156 & l1810;
assign a30260 = ~a30258 & a30256;
assign a30262 = a30096 & l1812;
assign a30264 = ~a30262 & a30260;
assign a30266 = a30226 & ~l1148;
assign a30268 = ~a30266 & a30264;
assign a30270 = a30170 & l1816;
assign a30272 = ~a30270 & a30268;
assign a30274 = a30236 & ~l1148;
assign a30276 = ~a30274 & a30272;
assign a30278 = a30182 & l1820;
assign a30280 = ~a30278 & a30276;
assign a30282 = a30132 & l1804;
assign a30284 = ~a30282 & a30280;
assign a30286 = a30206 & a30138;
assign a30288 = ~a30286 & a30284;
assign a30290 = ~a30288 & l1150;
assign a30292 = ~a30290 & ~a30250;
assign a30294 = a30292 & ~a17494;
assign a30296 = ~a30294 & ~a30200;
assign a30298 = ~a30292 & a17494;
assign a30300 = ~a30298 & ~a30296;
assign a30302 = ~a19026 & a6538;
assign a30304 = a30302 & l1148;
assign a30306 = ~a19010 & ~l1166;
assign a30308 = a30306 & a30080;
assign a30310 = ~a30308 & ~a30304;
assign a30312 = l1830 & ~l1166;
assign a30314 = a30312 & a30086;
assign a30316 = ~a30314 & a30310;
assign a30318 = a30096 & l1832;
assign a30320 = ~a30318 & a30316;
assign a30322 = a30104 & l1834;
assign a30324 = ~a30322 & a30320;
assign a30326 = a30102 & l1836;
assign a30328 = a30326 & l1148;
assign a30330 = ~a30328 & a30324;
assign a30332 = a30120 & l1838;
assign a30334 = ~a30332 & a30330;
assign a30336 = a6522 & l1840;
assign a30338 = a30336 & l1148;
assign a30340 = ~a30338 & a30334;
assign a30342 = a30132 & l1842;
assign a30344 = ~a30342 & a30340;
assign a30346 = a30140 & l1826;
assign a30348 = ~a30346 & a30344;
assign a30350 = ~a30348 & ~l1150;
assign a30352 = a30312 & a30148;
assign a30354 = a30302 & ~l1148;
assign a30356 = ~a30354 & ~a30352;
assign a30358 = a30156 & l1832;
assign a30360 = ~a30358 & a30356;
assign a30362 = a30096 & l1834;
assign a30364 = ~a30362 & a30360;
assign a30366 = a30326 & ~l1148;
assign a30368 = ~a30366 & a30364;
assign a30370 = a30170 & l1838;
assign a30372 = ~a30370 & a30368;
assign a30374 = a30336 & ~l1148;
assign a30376 = ~a30374 & a30372;
assign a30378 = a30182 & l1842;
assign a30380 = ~a30378 & a30376;
assign a30382 = a30132 & l1826;
assign a30384 = ~a30382 & a30380;
assign a30386 = a30306 & a30138;
assign a30388 = ~a30386 & a30384;
assign a30390 = ~a30388 & l1150;
assign a30392 = ~a30390 & ~a30350;
assign a30394 = a30392 & ~a17518;
assign a30396 = ~a30394 & ~a30300;
assign a30398 = ~a30392 & a17518;
assign a30400 = ~a30398 & ~a30396;
assign a30402 = ~a19108 & a6538;
assign a30404 = a30402 & l1148;
assign a30406 = ~a19092 & ~l1166;
assign a30408 = a30406 & a30080;
assign a30410 = ~a30408 & ~a30404;
assign a30412 = l1852 & ~l1166;
assign a30414 = a30412 & a30086;
assign a30416 = ~a30414 & a30410;
assign a30418 = a30096 & l1854;
assign a30420 = ~a30418 & a30416;
assign a30422 = a30104 & l1856;
assign a30424 = ~a30422 & a30420;
assign a30426 = a30102 & l1858;
assign a30428 = a30426 & l1148;
assign a30430 = ~a30428 & a30424;
assign a30432 = a30120 & l1860;
assign a30434 = ~a30432 & a30430;
assign a30436 = a6522 & l1862;
assign a30438 = a30436 & l1148;
assign a30440 = ~a30438 & a30434;
assign a30442 = a30132 & l1864;
assign a30444 = ~a30442 & a30440;
assign a30446 = a30140 & l1848;
assign a30448 = ~a30446 & a30444;
assign a30450 = ~a30448 & ~l1150;
assign a30452 = a30412 & a30148;
assign a30454 = a30402 & ~l1148;
assign a30456 = ~a30454 & ~a30452;
assign a30458 = a30156 & l1854;
assign a30460 = ~a30458 & a30456;
assign a30462 = a30096 & l1856;
assign a30464 = ~a30462 & a30460;
assign a30466 = a30426 & ~l1148;
assign a30468 = ~a30466 & a30464;
assign a30470 = a30170 & l1860;
assign a30472 = ~a30470 & a30468;
assign a30474 = a30436 & ~l1148;
assign a30476 = ~a30474 & a30472;
assign a30478 = a30182 & l1864;
assign a30480 = ~a30478 & a30476;
assign a30482 = a30132 & l1848;
assign a30484 = ~a30482 & a30480;
assign a30486 = a30406 & a30138;
assign a30488 = ~a30486 & a30484;
assign a30490 = ~a30488 & l1150;
assign a30492 = ~a30490 & ~a30450;
assign a30494 = a30492 & ~a17542;
assign a30496 = ~a30494 & ~a30400;
assign a30498 = ~a30492 & a17542;
assign a30500 = ~a30498 & ~a30496;
assign a30502 = ~a19190 & a6538;
assign a30504 = a30502 & l1148;
assign a30506 = ~a19174 & ~l1166;
assign a30508 = a30506 & a30080;
assign a30510 = ~a30508 & ~a30504;
assign a30512 = l1874 & ~l1166;
assign a30514 = a30512 & a30086;
assign a30516 = ~a30514 & a30510;
assign a30518 = a30096 & l1876;
assign a30520 = ~a30518 & a30516;
assign a30522 = a30104 & l1878;
assign a30524 = ~a30522 & a30520;
assign a30526 = a30102 & l1880;
assign a30528 = a30526 & l1148;
assign a30530 = ~a30528 & a30524;
assign a30532 = a30120 & l1882;
assign a30534 = ~a30532 & a30530;
assign a30536 = a6522 & l1884;
assign a30538 = a30536 & l1148;
assign a30540 = ~a30538 & a30534;
assign a30542 = a30132 & l1886;
assign a30544 = ~a30542 & a30540;
assign a30546 = a30140 & l1870;
assign a30548 = ~a30546 & a30544;
assign a30550 = ~a30548 & ~l1150;
assign a30552 = a30512 & a30148;
assign a30554 = a30502 & ~l1148;
assign a30556 = ~a30554 & ~a30552;
assign a30558 = a30156 & l1876;
assign a30560 = ~a30558 & a30556;
assign a30562 = a30096 & l1878;
assign a30564 = ~a30562 & a30560;
assign a30566 = a30526 & ~l1148;
assign a30568 = ~a30566 & a30564;
assign a30570 = a30170 & l1882;
assign a30572 = ~a30570 & a30568;
assign a30574 = a30536 & ~l1148;
assign a30576 = ~a30574 & a30572;
assign a30578 = a30182 & l1886;
assign a30580 = ~a30578 & a30576;
assign a30582 = a30132 & l1870;
assign a30584 = ~a30582 & a30580;
assign a30586 = a30506 & a30138;
assign a30588 = ~a30586 & a30584;
assign a30590 = ~a30588 & l1150;
assign a30592 = ~a30590 & ~a30550;
assign a30594 = a30592 & ~a17566;
assign a30596 = ~a30594 & ~a30500;
assign a30598 = ~a30592 & a17566;
assign a30600 = ~a30598 & ~a30596;
assign a30602 = ~a19272 & a6538;
assign a30604 = a30602 & l1148;
assign a30606 = ~a19256 & ~l1166;
assign a30608 = a30606 & a30080;
assign a30610 = ~a30608 & ~a30604;
assign a30612 = l1896 & ~l1166;
assign a30614 = a30612 & a30086;
assign a30616 = ~a30614 & a30610;
assign a30618 = a30096 & l1898;
assign a30620 = ~a30618 & a30616;
assign a30622 = a30104 & l1900;
assign a30624 = ~a30622 & a30620;
assign a30626 = a30102 & l1902;
assign a30628 = a30626 & l1148;
assign a30630 = ~a30628 & a30624;
assign a30632 = a30120 & l1904;
assign a30634 = ~a30632 & a30630;
assign a30636 = a6522 & l1906;
assign a30638 = a30636 & l1148;
assign a30640 = ~a30638 & a30634;
assign a30642 = a30132 & l1908;
assign a30644 = ~a30642 & a30640;
assign a30646 = a30140 & l1892;
assign a30648 = ~a30646 & a30644;
assign a30650 = ~a30648 & ~l1150;
assign a30652 = a30612 & a30148;
assign a30654 = a30602 & ~l1148;
assign a30656 = ~a30654 & ~a30652;
assign a30658 = a30156 & l1898;
assign a30660 = ~a30658 & a30656;
assign a30662 = a30096 & l1900;
assign a30664 = ~a30662 & a30660;
assign a30666 = a30626 & ~l1148;
assign a30668 = ~a30666 & a30664;
assign a30670 = a30170 & l1904;
assign a30672 = ~a30670 & a30668;
assign a30674 = a30636 & ~l1148;
assign a30676 = ~a30674 & a30672;
assign a30678 = a30182 & l1908;
assign a30680 = ~a30678 & a30676;
assign a30682 = a30132 & l1892;
assign a30684 = ~a30682 & a30680;
assign a30686 = a30606 & a30138;
assign a30688 = ~a30686 & a30684;
assign a30690 = ~a30688 & l1150;
assign a30692 = ~a30690 & ~a30650;
assign a30694 = a30692 & ~a17592;
assign a30696 = ~a30694 & ~a30600;
assign a30698 = ~a30692 & a17592;
assign a30700 = ~a30698 & ~a30696;
assign a30702 = ~a19348 & a6538;
assign a30704 = a30702 & l1148;
assign a30706 = l1910 & ~l1166;
assign a30708 = a30706 & a30080;
assign a30710 = ~a30708 & ~a30704;
assign a30712 = l1918 & ~l1166;
assign a30714 = a30712 & a30086;
assign a30716 = ~a30714 & a30710;
assign a30718 = a30096 & l1920;
assign a30720 = ~a30718 & a30716;
assign a30722 = a30104 & l1922;
assign a30724 = ~a30722 & a30720;
assign a30726 = a30102 & l1924;
assign a30728 = a30726 & l1148;
assign a30730 = ~a30728 & a30724;
assign a30732 = a30120 & l1926;
assign a30734 = ~a30732 & a30730;
assign a30736 = a6522 & l1928;
assign a30738 = a30736 & l1148;
assign a30740 = ~a30738 & a30734;
assign a30742 = a30132 & l1930;
assign a30744 = ~a30742 & a30740;
assign a30746 = a30140 & l1914;
assign a30748 = ~a30746 & a30744;
assign a30750 = ~a30748 & ~l1150;
assign a30752 = a30712 & a30148;
assign a30754 = a30702 & ~l1148;
assign a30756 = ~a30754 & ~a30752;
assign a30758 = a30156 & l1920;
assign a30760 = ~a30758 & a30756;
assign a30762 = a30096 & l1922;
assign a30764 = ~a30762 & a30760;
assign a30766 = a30726 & ~l1148;
assign a30768 = ~a30766 & a30764;
assign a30770 = a30170 & l1926;
assign a30772 = ~a30770 & a30768;
assign a30774 = a30736 & ~l1148;
assign a30776 = ~a30774 & a30772;
assign a30778 = a30182 & l1930;
assign a30780 = ~a30778 & a30776;
assign a30782 = a30132 & l1914;
assign a30784 = ~a30782 & a30780;
assign a30786 = a30706 & a30138;
assign a30788 = ~a30786 & a30784;
assign a30790 = ~a30788 & l1150;
assign a30792 = ~a30790 & ~a30750;
assign a30794 = a30792 & ~a17616;
assign a30796 = ~a30794 & ~a30700;
assign a30798 = ~a30792 & a17616;
assign a30800 = a6538 & l1938;
assign a30802 = a30800 & l1148;
assign a30804 = l1932 & ~l1166;
assign a30806 = a30804 & a30080;
assign a30808 = ~a30806 & ~a30802;
assign a30810 = l1940 & ~l1166;
assign a30812 = a30810 & a30086;
assign a30814 = ~a30812 & a30808;
assign a30816 = a30096 & l1942;
assign a30818 = ~a30816 & a30814;
assign a30820 = a30104 & l1944;
assign a30822 = ~a30820 & a30818;
assign a30824 = a30102 & l1946;
assign a30826 = a30824 & l1148;
assign a30828 = ~a30826 & a30822;
assign a30830 = a30120 & l1948;
assign a30832 = ~a30830 & a30828;
assign a30834 = a6522 & l1950;
assign a30836 = a30834 & l1148;
assign a30838 = ~a30836 & a30832;
assign a30840 = a30132 & l1952;
assign a30842 = ~a30840 & a30838;
assign a30844 = a30140 & l1936;
assign a30846 = ~a30844 & a30842;
assign a30848 = ~a30846 & ~l1150;
assign a30850 = a30810 & a30148;
assign a30852 = a30800 & ~l1148;
assign a30854 = ~a30852 & ~a30850;
assign a30856 = a30156 & l1942;
assign a30858 = ~a30856 & a30854;
assign a30860 = a30096 & l1944;
assign a30862 = ~a30860 & a30858;
assign a30864 = a30824 & ~l1148;
assign a30866 = ~a30864 & a30862;
assign a30868 = a30170 & l1948;
assign a30870 = ~a30868 & a30866;
assign a30872 = a30834 & ~l1148;
assign a30874 = ~a30872 & a30870;
assign a30876 = a30182 & l1952;
assign a30878 = ~a30876 & a30874;
assign a30880 = a30132 & l1936;
assign a30882 = ~a30880 & a30878;
assign a30884 = a30804 & a30138;
assign a30886 = ~a30884 & a30882;
assign a30888 = ~a30886 & l1150;
assign a30890 = ~a30888 & ~a30848;
assign a30892 = a30890 & ~a17454;
assign a30894 = ~a30890 & a17454;
assign a30896 = ~a30894 & ~a30892;
assign a30898 = ~a30896 & ~a30798;
assign a30900 = a30898 & ~a30796;
assign a30902 = ~a30198 & a17476;
assign a30904 = ~a30902 & ~a30298;
assign a30906 = ~a30904 & ~a30294;
assign a30908 = ~a30906 & ~a30398;
assign a30910 = ~a30908 & ~a30394;
assign a30912 = ~a30910 & ~a30498;
assign a30914 = ~a30912 & ~a30494;
assign a30916 = ~a30914 & ~a30598;
assign a30918 = ~a30916 & ~a30594;
assign a30920 = ~a30918 & ~a30698;
assign a30922 = ~a30920 & ~a30694;
assign a30924 = ~a30922 & ~a30798;
assign a30926 = ~a30924 & ~a30794;
assign a30928 = a30926 & a30896;
assign a30930 = a30148 & ~l1166;
assign a30932 = a30930 & a18596;
assign a30934 = a30080 & ~l1166;
assign a30936 = a30934 & a18568;
assign a30938 = ~a30936 & ~a30932;
assign a30940 = a30156 & l1974;
assign a30942 = ~a30940 & a30938;
assign a30944 = a30096 & l1976;
assign a30946 = ~a30944 & a30942;
assign a30948 = a30104 & l1978;
assign a30950 = ~a30948 & a30946;
assign a30952 = a30170 & l1980;
assign a30954 = ~a30952 & a30950;
assign a30956 = a30120 & l1982;
assign a30958 = ~a30956 & a30954;
assign a30960 = a30182 & a18646;
assign a30962 = ~a30960 & a30958;
assign a30964 = a30132 & l1986;
assign a30966 = ~a30964 & a30962;
assign a30968 = a30140 & a18582;
assign a30970 = ~a30968 & a30966;
assign a30972 = ~a30970 & ~l1150;
assign a30974 = a30930 & l1974;
assign a30976 = a30934 & a18596;
assign a30978 = ~a30976 & ~a30974;
assign a30980 = a30156 & l1976;
assign a30982 = ~a30980 & a30978;
assign a30984 = a30096 & l1978;
assign a30986 = ~a30984 & a30982;
assign a30988 = a30104 & l1980;
assign a30990 = ~a30988 & a30986;
assign a30992 = a30170 & l1982;
assign a30994 = ~a30992 & a30990;
assign a30996 = a30120 & a18646;
assign a30998 = ~a30996 & a30994;
assign a31000 = a30182 & l1986;
assign a31002 = ~a31000 & a30998;
assign a31004 = a30132 & a18582;
assign a31006 = ~a31004 & a31002;
assign a31008 = a30140 & a18568;
assign a31010 = ~a31008 & a31006;
assign a31012 = ~a31010 & l1150;
assign a31014 = ~a31012 & ~a30972;
assign a31016 = ~a31014 & ~a30928;
assign a31022 = a19876 & a2768;
assign a31024 = a31022 & ~l1244;
assign a31026 = a31024 & ~a2740;
assign a31028 = a31026 & ~l1156;
assign a31030 = ~a31028 & ~a18872;
assign a31032 = ~l1782 & l890;
assign a31034 = ~a11250 & ~l890;
assign a31036 = ~a31034 & ~a31032;
assign a31038 = ~a31036 & a31028;
assign a31044 = ~a31042 & l1156;
assign a31046 = a31042 & ~a21682;
assign a31048 = ~a31046 & ~a31044;
assign a31050 = ~a2748 & l884;
assign a31052 = a30062 & l1162;
assign a31054 = ~a30148 & ~a30086;
assign a31056 = ~a31054 & a30066;
assign a31058 = ~a31056 & ~a31052;
assign a31060 = a31058 & ~a31050;
assign a31062 = ~a2512 & l884;
assign a31064 = a30062 & l1164;
assign a31066 = ~a30180 & ~a30132;
assign a31068 = ~a31066 & a30066;
assign a31070 = ~a31068 & ~a31064;
assign a31072 = a31070 & ~a31062;
assign a31074 = ~a2532 & l884;
assign a31076 = a30062 & l1166;
assign a31078 = ~a30116 & ~a30096;
assign a31080 = a31078 & ~a30102;
assign a31082 = ~a31080 & a30066;
assign a31084 = ~a31082 & ~a31076;
assign a31086 = a31084 & ~a31074;
assign a31090 = l1186 & ~l880;
assign a31092 = ~a31090 & ~l1188;
assign a31094 = ~l1190 & ~l884;
assign a31096 = ~a31092 & a2768;
assign a31098 = a31092 & ~a2768;
assign a31100 = ~a2748 & l1186;
assign a31102 = ~a31100 & ~l1210;
assign a31104 = ~a31102 & a2740;
assign a31106 = a31102 & ~a2740;
assign a31108 = ~a2532 & l1186;
assign a31110 = ~a31108 & ~l1226;
assign a31112 = ~a31110 & ~l1156;
assign a31114 = a31110 & l1156;
assign a31116 = ~a2512 & l1186;
assign a31118 = ~a31116 & ~l1242;
assign a31120 = ~a31118 & ~l1244;
assign a31122 = a31118 & l1244;
assign a31124 = ~a31122 & ~a31120;
assign a31126 = a31124 & ~a31114;
assign a31128 = a31126 & ~a31112;
assign a31130 = a31128 & ~a31106;
assign a31132 = a31130 & ~a31104;
assign a31134 = a31132 & ~a31098;
assign a31136 = a31134 & ~a31096;
assign a31138 = ~a31136 & l1248;
assign a31140 = ~a31138 & ~l1102;
assign a31142 = a31140 & a31094;
assign a31144 = a31142 & ~a31092;
assign a31146 = a31138 & a31094;
assign a31148 = a31146 & a31092;
assign a31150 = ~a31148 & ~l2054;
assign a31152 = a31150 & ~a31144;
assign a31154 = ~a9052 & ~a9046;
assign a31156 = ~a31154 & ~a16190;
assign a31158 = ~a31156 & ~a18552;
assign a31162 = a31142 & ~a31102;
assign a31164 = a31118 & ~a31092;
assign a31166 = a31164 & a31102;
assign a31168 = ~a31102 & a31092;
assign a31170 = ~a31168 & ~a31166;
assign a31172 = ~a31170 & a31146;
assign a31174 = ~a31172 & ~l2050;
assign a31176 = a31174 & ~a31162;
assign a31178 = ~a31042 & ~a2768;
assign a31180 = a31042 & ~a21676;
assign a31184 = a31142 & ~a31110;
assign a31186 = ~a31110 & a31102;
assign a31188 = ~a31110 & a31092;
assign a31190 = ~a31102 & ~a31092;
assign a31192 = a31190 & a31110;
assign a31194 = ~a31192 & ~a31188;
assign a31196 = a31194 & ~a31186;
assign a31198 = ~a31196 & a31146;
assign a31200 = ~a31198 & ~l2046;
assign a31202 = a31200 & ~a31184;
assign a31204 = ~a31042 & ~a2740;
assign a31206 = a31042 & ~a21688;
assign a31210 = a31142 & ~a31118;
assign a31212 = a31190 & ~a31110;
assign a31214 = ~a31118 & a31092;
assign a31216 = ~a31214 & ~a31212;
assign a31218 = ~a31216 & a31146;
assign a31220 = ~a31218 & ~l2026;
assign a31222 = a31220 & ~a31210;
assign a31224 = ~a31042 & l1244;
assign a31226 = a31042 & ~a21698;
assign a31228 = ~a31226 & ~a31224;
assign a31230 = a31110 & a31102;
assign a31232 = a31230 & l1784;
assign a31234 = a31232 & ~a31118;
assign a31236 = a31234 & ~a31092;
assign a31238 = a31230 & ~a31118;
assign a31240 = a31238 & l1798;
assign a31242 = a31240 & a31092;
assign a31244 = a31118 & ~a31110;
assign a31246 = a31244 & ~a31102;
assign a31248 = a31246 & l1796;
assign a31250 = a31248 & ~a31092;
assign a31252 = a31244 & l1794;
assign a31254 = a31252 & ~a31102;
assign a31256 = a31254 & a31092;
assign a31258 = a31244 & l1792;
assign a31260 = a31102 & ~a31092;
assign a31262 = a31260 & a31258;
assign a31264 = a31118 & l1790;
assign a31266 = a31186 & a31092;
assign a31268 = a31266 & a31264;
assign a31270 = a31110 & ~a31102;
assign a31272 = a31118 & l1788;
assign a31274 = a31272 & a31270;
assign a31276 = a31274 & ~a31092;
assign a31278 = a31118 & a31110;
assign a31280 = a31278 & l1786;
assign a31282 = a31280 & ~a31102;
assign a31284 = a31282 & a31092;
assign a31286 = a31278 & ~a18872;
assign a31288 = a31286 & a31260;
assign a31290 = a31230 & ~a18856;
assign a31292 = a31118 & a31092;
assign a31294 = a31292 & a31290;
assign a31296 = ~a31294 & ~a31288;
assign a31298 = a31296 & ~a31284;
assign a31300 = a31298 & ~a31276;
assign a31302 = a31300 & ~a31268;
assign a31304 = a31302 & ~a31262;
assign a31306 = a31304 & ~a31256;
assign a31308 = a31306 & ~a31250;
assign a31310 = a31308 & ~a31242;
assign a31312 = a31310 & ~a31236;
assign a31314 = ~a31312 & ~a31138;
assign a31316 = a31280 & a31260;
assign a31318 = a31286 & a31092;
assign a31320 = a31318 & a31102;
assign a31322 = ~a31320 & ~a31316;
assign a31324 = a31274 & a31092;
assign a31326 = ~a31324 & a31322;
assign a31328 = a31264 & ~a31092;
assign a31330 = a31328 & a31270;
assign a31332 = ~a31330 & a31326;
assign a31334 = a31258 & a31092;
assign a31336 = a31334 & a31102;
assign a31338 = ~a31336 & a31332;
assign a31340 = a31260 & a31252;
assign a31342 = ~a31340 & a31338;
assign a31344 = a31248 & a31092;
assign a31346 = ~a31344 & a31342;
assign a31348 = a31246 & ~a31092;
assign a31350 = a31348 & l1798;
assign a31352 = ~a31350 & a31346;
assign a31354 = a31234 & a31092;
assign a31356 = ~a31354 & a31352;
assign a31358 = a31290 & ~a31092;
assign a31360 = a31358 & ~a31118;
assign a31362 = ~a31360 & a31356;
assign a31364 = ~a31362 & a31138;
assign a31366 = ~a31364 & ~a31314;
assign a31368 = a31366 & ~a17856;
assign a31370 = ~a31366 & a17856;
assign a31372 = a31230 & l1804;
assign a31374 = a31372 & ~a31118;
assign a31376 = a31374 & ~a31092;
assign a31378 = a31238 & l1820;
assign a31380 = a31378 & a31092;
assign a31382 = a31246 & l1818;
assign a31384 = a31382 & ~a31092;
assign a31386 = a31244 & l1816;
assign a31388 = a31386 & ~a31102;
assign a31390 = a31388 & a31092;
assign a31392 = a31244 & l1814;
assign a31394 = a31392 & a31260;
assign a31396 = a31118 & l1812;
assign a31398 = a31396 & a31266;
assign a31400 = a31118 & l1810;
assign a31402 = a31400 & a31270;
assign a31404 = a31402 & ~a31092;
assign a31406 = a31278 & l1808;
assign a31408 = a31406 & ~a31102;
assign a31410 = a31408 & a31092;
assign a31412 = a31278 & ~a18946;
assign a31414 = a31412 & a31260;
assign a31416 = a31230 & ~a18930;
assign a31418 = a31416 & a31292;
assign a31420 = ~a31418 & ~a31414;
assign a31422 = a31420 & ~a31410;
assign a31424 = a31422 & ~a31404;
assign a31426 = a31424 & ~a31398;
assign a31428 = a31426 & ~a31394;
assign a31430 = a31428 & ~a31390;
assign a31432 = a31430 & ~a31384;
assign a31434 = a31432 & ~a31380;
assign a31436 = a31434 & ~a31376;
assign a31438 = ~a31436 & ~a31138;
assign a31440 = a31406 & a31260;
assign a31442 = a31412 & a31092;
assign a31444 = a31442 & a31102;
assign a31446 = ~a31444 & ~a31440;
assign a31448 = a31402 & a31092;
assign a31450 = ~a31448 & a31446;
assign a31452 = a31396 & ~a31092;
assign a31454 = a31452 & a31270;
assign a31456 = ~a31454 & a31450;
assign a31458 = a31392 & a31092;
assign a31460 = a31458 & a31102;
assign a31462 = ~a31460 & a31456;
assign a31464 = a31386 & a31260;
assign a31466 = ~a31464 & a31462;
assign a31468 = a31382 & a31092;
assign a31470 = ~a31468 & a31466;
assign a31472 = a31348 & l1820;
assign a31474 = ~a31472 & a31470;
assign a31476 = a31374 & a31092;
assign a31478 = ~a31476 & a31474;
assign a31480 = a31416 & ~a31092;
assign a31482 = a31480 & ~a31118;
assign a31484 = ~a31482 & a31478;
assign a31486 = ~a31484 & a31138;
assign a31488 = ~a31486 & ~a31438;
assign a31490 = a31488 & ~a17924;
assign a31492 = ~a31488 & a17924;
assign a31494 = a31230 & l1826;
assign a31496 = a31494 & ~a31118;
assign a31498 = a31496 & ~a31092;
assign a31500 = a31238 & l1842;
assign a31502 = a31500 & a31092;
assign a31504 = a31246 & l1840;
assign a31506 = a31504 & ~a31092;
assign a31508 = a31244 & l1838;
assign a31510 = a31508 & ~a31102;
assign a31512 = a31510 & a31092;
assign a31514 = a31244 & l1836;
assign a31516 = a31514 & a31260;
assign a31518 = a31118 & l1834;
assign a31520 = a31518 & a31266;
assign a31522 = a31118 & l1832;
assign a31524 = a31522 & a31270;
assign a31526 = a31524 & ~a31092;
assign a31528 = a31278 & l1830;
assign a31530 = a31528 & ~a31102;
assign a31532 = a31530 & a31092;
assign a31534 = a31278 & ~a19026;
assign a31536 = a31534 & a31260;
assign a31538 = a31230 & ~a19010;
assign a31540 = a31538 & a31292;
assign a31542 = ~a31540 & ~a31536;
assign a31544 = a31542 & ~a31532;
assign a31546 = a31544 & ~a31526;
assign a31548 = a31546 & ~a31520;
assign a31550 = a31548 & ~a31516;
assign a31552 = a31550 & ~a31512;
assign a31554 = a31552 & ~a31506;
assign a31556 = a31554 & ~a31502;
assign a31558 = a31556 & ~a31498;
assign a31560 = ~a31558 & ~a31138;
assign a31562 = a31528 & a31260;
assign a31564 = a31534 & a31092;
assign a31566 = a31564 & a31102;
assign a31568 = ~a31566 & ~a31562;
assign a31570 = a31524 & a31092;
assign a31572 = ~a31570 & a31568;
assign a31574 = a31518 & ~a31092;
assign a31576 = a31574 & a31270;
assign a31578 = ~a31576 & a31572;
assign a31580 = a31514 & a31092;
assign a31582 = a31580 & a31102;
assign a31584 = ~a31582 & a31578;
assign a31586 = a31508 & a31260;
assign a31588 = ~a31586 & a31584;
assign a31590 = a31504 & a31092;
assign a31592 = ~a31590 & a31588;
assign a31594 = a31348 & l1842;
assign a31596 = ~a31594 & a31592;
assign a31598 = a31496 & a31092;
assign a31600 = ~a31598 & a31596;
assign a31602 = a31538 & ~a31092;
assign a31604 = a31602 & ~a31118;
assign a31606 = ~a31604 & a31600;
assign a31608 = ~a31606 & a31138;
assign a31610 = ~a31608 & ~a31560;
assign a31612 = a31610 & ~a17998;
assign a31614 = ~a31610 & a17998;
assign a31616 = a31230 & l1848;
assign a31618 = a31616 & ~a31118;
assign a31620 = a31618 & ~a31092;
assign a31622 = a31238 & l1864;
assign a31624 = a31622 & a31092;
assign a31626 = a31246 & l1862;
assign a31628 = a31626 & ~a31092;
assign a31630 = a31244 & l1860;
assign a31632 = a31630 & ~a31102;
assign a31634 = a31632 & a31092;
assign a31636 = a31244 & l1858;
assign a31638 = a31636 & a31260;
assign a31640 = a31118 & l1856;
assign a31642 = a31640 & a31266;
assign a31644 = a31118 & l1854;
assign a31646 = a31644 & a31270;
assign a31648 = a31646 & ~a31092;
assign a31650 = a31278 & l1852;
assign a31652 = a31650 & ~a31102;
assign a31654 = a31652 & a31092;
assign a31656 = a31278 & ~a19108;
assign a31658 = a31656 & a31260;
assign a31660 = a31230 & ~a19092;
assign a31662 = a31660 & a31292;
assign a31664 = ~a31662 & ~a31658;
assign a31666 = a31664 & ~a31654;
assign a31668 = a31666 & ~a31648;
assign a31670 = a31668 & ~a31642;
assign a31672 = a31670 & ~a31638;
assign a31674 = a31672 & ~a31634;
assign a31676 = a31674 & ~a31628;
assign a31678 = a31676 & ~a31624;
assign a31680 = a31678 & ~a31620;
assign a31682 = ~a31680 & ~a31138;
assign a31684 = a31650 & a31260;
assign a31686 = a31656 & a31092;
assign a31688 = a31686 & a31102;
assign a31690 = ~a31688 & ~a31684;
assign a31692 = a31646 & a31092;
assign a31694 = ~a31692 & a31690;
assign a31696 = a31640 & ~a31092;
assign a31698 = a31696 & a31270;
assign a31700 = ~a31698 & a31694;
assign a31702 = a31636 & a31092;
assign a31704 = a31702 & a31102;
assign a31706 = ~a31704 & a31700;
assign a31708 = a31630 & a31260;
assign a31710 = ~a31708 & a31706;
assign a31712 = a31626 & a31092;
assign a31714 = ~a31712 & a31710;
assign a31716 = a31348 & l1864;
assign a31718 = ~a31716 & a31714;
assign a31720 = a31618 & a31092;
assign a31722 = ~a31720 & a31718;
assign a31724 = a31660 & ~a31092;
assign a31726 = a31724 & ~a31118;
assign a31728 = ~a31726 & a31722;
assign a31730 = ~a31728 & a31138;
assign a31732 = ~a31730 & ~a31682;
assign a31734 = a31732 & ~a18072;
assign a31736 = ~a31732 & a18072;
assign a31738 = a31230 & l1870;
assign a31740 = a31738 & ~a31118;
assign a31742 = a31740 & ~a31092;
assign a31744 = a31238 & l1886;
assign a31746 = a31744 & a31092;
assign a31748 = a31246 & l1884;
assign a31750 = a31748 & ~a31092;
assign a31752 = a31244 & l1882;
assign a31754 = a31752 & ~a31102;
assign a31756 = a31754 & a31092;
assign a31758 = a31244 & l1880;
assign a31760 = a31758 & a31260;
assign a31762 = a31118 & l1878;
assign a31764 = a31762 & a31266;
assign a31766 = a31118 & l1876;
assign a31768 = a31766 & a31270;
assign a31770 = a31768 & ~a31092;
assign a31772 = a31278 & l1874;
assign a31774 = a31772 & ~a31102;
assign a31776 = a31774 & a31092;
assign a31778 = a31278 & ~a19190;
assign a31780 = a31778 & a31260;
assign a31782 = a31230 & ~a19174;
assign a31784 = a31782 & a31292;
assign a31786 = ~a31784 & ~a31780;
assign a31788 = a31786 & ~a31776;
assign a31790 = a31788 & ~a31770;
assign a31792 = a31790 & ~a31764;
assign a31794 = a31792 & ~a31760;
assign a31796 = a31794 & ~a31756;
assign a31798 = a31796 & ~a31750;
assign a31800 = a31798 & ~a31746;
assign a31802 = a31800 & ~a31742;
assign a31804 = ~a31802 & ~a31138;
assign a31806 = a31772 & a31260;
assign a31808 = a31778 & a31092;
assign a31810 = a31808 & a31102;
assign a31812 = ~a31810 & ~a31806;
assign a31814 = a31768 & a31092;
assign a31816 = ~a31814 & a31812;
assign a31818 = a31762 & ~a31092;
assign a31820 = a31818 & a31270;
assign a31822 = ~a31820 & a31816;
assign a31824 = a31758 & a31092;
assign a31826 = a31824 & a31102;
assign a31828 = ~a31826 & a31822;
assign a31830 = a31752 & a31260;
assign a31832 = ~a31830 & a31828;
assign a31834 = a31748 & a31092;
assign a31836 = ~a31834 & a31832;
assign a31838 = a31348 & l1886;
assign a31840 = ~a31838 & a31836;
assign a31842 = a31740 & a31092;
assign a31844 = ~a31842 & a31840;
assign a31846 = a31782 & ~a31092;
assign a31848 = a31846 & ~a31118;
assign a31850 = ~a31848 & a31844;
assign a31852 = ~a31850 & a31138;
assign a31854 = ~a31852 & ~a31804;
assign a31856 = a31854 & ~a18146;
assign a31858 = ~a31854 & a18146;
assign a31860 = a31230 & l1892;
assign a31862 = a31860 & ~a31118;
assign a31864 = a31862 & ~a31092;
assign a31866 = a31238 & l1908;
assign a31868 = a31866 & a31092;
assign a31870 = a31246 & l1906;
assign a31872 = a31870 & ~a31092;
assign a31874 = a31244 & l1904;
assign a31876 = a31874 & ~a31102;
assign a31878 = a31876 & a31092;
assign a31880 = a31244 & l1902;
assign a31882 = a31880 & a31260;
assign a31884 = a31118 & l1900;
assign a31886 = a31884 & a31266;
assign a31888 = a31118 & l1898;
assign a31890 = a31888 & a31270;
assign a31892 = a31890 & ~a31092;
assign a31894 = a31278 & l1896;
assign a31896 = a31894 & ~a31102;
assign a31898 = a31896 & a31092;
assign a31900 = a31278 & ~a19272;
assign a31902 = a31900 & a31260;
assign a31904 = a31230 & ~a19256;
assign a31906 = a31904 & a31292;
assign a31908 = ~a31906 & ~a31902;
assign a31910 = a31908 & ~a31898;
assign a31912 = a31910 & ~a31892;
assign a31914 = a31912 & ~a31886;
assign a31916 = a31914 & ~a31882;
assign a31918 = a31916 & ~a31878;
assign a31920 = a31918 & ~a31872;
assign a31922 = a31920 & ~a31868;
assign a31924 = a31922 & ~a31864;
assign a31926 = ~a31924 & ~a31138;
assign a31928 = a31894 & a31260;
assign a31930 = a31900 & a31092;
assign a31932 = a31930 & a31102;
assign a31934 = ~a31932 & ~a31928;
assign a31936 = a31890 & a31092;
assign a31938 = ~a31936 & a31934;
assign a31940 = a31884 & ~a31092;
assign a31942 = a31940 & a31270;
assign a31944 = ~a31942 & a31938;
assign a31946 = a31880 & a31092;
assign a31948 = a31946 & a31102;
assign a31950 = ~a31948 & a31944;
assign a31952 = a31874 & a31260;
assign a31954 = ~a31952 & a31950;
assign a31956 = a31870 & a31092;
assign a31958 = ~a31956 & a31954;
assign a31960 = a31348 & l1908;
assign a31962 = ~a31960 & a31958;
assign a31964 = a31862 & a31092;
assign a31966 = ~a31964 & a31962;
assign a31968 = a31904 & ~a31092;
assign a31970 = a31968 & ~a31118;
assign a31972 = ~a31970 & a31966;
assign a31974 = ~a31972 & a31138;
assign a31976 = ~a31974 & ~a31926;
assign a31978 = a31976 & ~a18220;
assign a31980 = ~a31976 & a18220;
assign a31982 = a31230 & l1914;
assign a31984 = a31982 & ~a31118;
assign a31986 = a31984 & ~a31092;
assign a31988 = a31238 & l1930;
assign a31990 = a31988 & a31092;
assign a31992 = a31246 & l1928;
assign a31994 = a31992 & ~a31092;
assign a31996 = a31244 & l1926;
assign a31998 = a31996 & ~a31102;
assign a32000 = a31998 & a31092;
assign a32002 = a31244 & l1924;
assign a32004 = a32002 & a31260;
assign a32006 = a31118 & l1922;
assign a32008 = a32006 & a31266;
assign a32010 = a31118 & l1920;
assign a32012 = a32010 & a31270;
assign a32014 = a32012 & ~a31092;
assign a32016 = a31278 & l1918;
assign a32018 = a32016 & ~a31102;
assign a32020 = a32018 & a31092;
assign a32022 = a31278 & ~a19348;
assign a32024 = a32022 & a31260;
assign a32026 = a31230 & l1910;
assign a32028 = a32026 & a31292;
assign a32030 = ~a32028 & ~a32024;
assign a32032 = a32030 & ~a32020;
assign a32034 = a32032 & ~a32014;
assign a32036 = a32034 & ~a32008;
assign a32038 = a32036 & ~a32004;
assign a32040 = a32038 & ~a32000;
assign a32042 = a32040 & ~a31994;
assign a32044 = a32042 & ~a31990;
assign a32046 = a32044 & ~a31986;
assign a32048 = ~a32046 & ~a31138;
assign a32050 = a32016 & a31260;
assign a32052 = a32022 & a31092;
assign a32054 = a32052 & a31102;
assign a32056 = ~a32054 & ~a32050;
assign a32058 = a32012 & a31092;
assign a32060 = ~a32058 & a32056;
assign a32062 = a32006 & ~a31092;
assign a32064 = a32062 & a31270;
assign a32066 = ~a32064 & a32060;
assign a32068 = a32002 & a31092;
assign a32070 = a32068 & a31102;
assign a32072 = ~a32070 & a32066;
assign a32074 = a31996 & a31260;
assign a32076 = ~a32074 & a32072;
assign a32078 = a31992 & a31092;
assign a32080 = ~a32078 & a32076;
assign a32082 = a31348 & l1930;
assign a32084 = ~a32082 & a32080;
assign a32086 = a31984 & a31092;
assign a32088 = ~a32086 & a32084;
assign a32090 = a32026 & ~a31092;
assign a32092 = a32090 & ~a31118;
assign a32094 = ~a32092 & a32088;
assign a32096 = ~a32094 & a31138;
assign a32098 = ~a32096 & ~a32048;
assign a32100 = a32098 & ~a18294;
assign a32102 = ~a32098 & a18294;
assign a32104 = a31230 & l1936;
assign a32106 = a32104 & ~a31118;
assign a32108 = a32106 & ~a31092;
assign a32110 = a31238 & l1952;
assign a32112 = a32110 & a31092;
assign a32114 = a31246 & l1950;
assign a32116 = a32114 & ~a31092;
assign a32118 = a31244 & l1948;
assign a32120 = a32118 & ~a31102;
assign a32122 = a32120 & a31092;
assign a32124 = a31244 & l1946;
assign a32126 = a32124 & a31260;
assign a32128 = a31118 & l1944;
assign a32130 = a32128 & a31266;
assign a32132 = a31118 & l1942;
assign a32134 = a32132 & a31270;
assign a32136 = a32134 & ~a31092;
assign a32138 = a31278 & l1940;
assign a32140 = a32138 & ~a31102;
assign a32142 = a32140 & a31092;
assign a32144 = a31278 & l1938;
assign a32146 = a32144 & a31260;
assign a32148 = a31230 & l1932;
assign a32150 = a32148 & a31292;
assign a32152 = ~a32150 & ~a32146;
assign a32154 = a32152 & ~a32142;
assign a32156 = a32154 & ~a32136;
assign a32158 = a32156 & ~a32130;
assign a32160 = a32158 & ~a32126;
assign a32162 = a32160 & ~a32122;
assign a32164 = a32162 & ~a32116;
assign a32166 = a32164 & ~a32112;
assign a32168 = a32166 & ~a32108;
assign a32170 = ~a32168 & ~a31138;
assign a32172 = a32138 & a31260;
assign a32174 = a32144 & a31092;
assign a32176 = a32174 & a31102;
assign a32178 = ~a32176 & ~a32172;
assign a32180 = a32134 & a31092;
assign a32182 = ~a32180 & a32178;
assign a32184 = a32128 & ~a31092;
assign a32186 = a32184 & a31270;
assign a32188 = ~a32186 & a32182;
assign a32190 = a32124 & a31092;
assign a32192 = a32190 & a31102;
assign a32194 = ~a32192 & a32188;
assign a32196 = a32118 & a31260;
assign a32198 = ~a32196 & a32194;
assign a32200 = a32114 & a31092;
assign a32202 = ~a32200 & a32198;
assign a32204 = a31348 & l1952;
assign a32206 = ~a32204 & a32202;
assign a32208 = a32106 & a31092;
assign a32210 = ~a32208 & a32206;
assign a32212 = a32148 & ~a31092;
assign a32214 = a32212 & ~a31118;
assign a32216 = ~a32214 & a32210;
assign a32218 = ~a32216 & a31138;
assign a32220 = ~a32218 & ~a32170;
assign a32222 = a32220 & ~a17728;
assign a32224 = ~a32220 & a17728;
assign a32226 = a31238 & a18582;
assign a32228 = a32226 & ~a31092;
assign a32230 = a31238 & a31092;
assign a32232 = a32230 & l1986;
assign a32234 = a31246 & a18646;
assign a32236 = a32234 & ~a31092;
assign a32238 = a31246 & a31092;
assign a32240 = a32238 & l1982;
assign a32242 = a31244 & a31102;
assign a32244 = a32242 & ~a31092;
assign a32246 = a32244 & l1980;
assign a32248 = a32242 & a31092;
assign a32250 = a32248 & l1978;
assign a32252 = a31270 & a31118;
assign a32254 = a32252 & l1976;
assign a32256 = a32254 & ~a31092;
assign a32258 = a32252 & a31092;
assign a32260 = a32258 & l1974;
assign a32262 = a31278 & a31102;
assign a32264 = a32262 & ~a31092;
assign a32266 = a32264 & a18596;
assign a32268 = a32262 & a31092;
assign a32270 = a32268 & a18568;
assign a32272 = ~a32270 & ~a32266;
assign a32274 = a32272 & ~a32260;
assign a32276 = a32274 & ~a32256;
assign a32278 = a32276 & ~a32250;
assign a32280 = a32278 & ~a32246;
assign a32282 = a32280 & ~a32240;
assign a32284 = a32282 & ~a32236;
assign a32286 = a32284 & ~a32232;
assign a32288 = a32286 & ~a32228;
assign a32290 = ~a32288 & ~a31138;
assign a32292 = a31238 & ~a31092;
assign a32294 = a32292 & a18568;
assign a32296 = a32226 & a31092;
assign a32298 = a31348 & l1986;
assign a32300 = a32234 & a31092;
assign a32302 = a32244 & l1982;
assign a32304 = a32248 & l1980;
assign a32306 = a32252 & ~a31092;
assign a32308 = a32306 & l1978;
assign a32310 = a32254 & a31092;
assign a32312 = a32264 & l1974;
assign a32314 = a32268 & a18596;
assign a32316 = ~a32314 & ~a32312;
assign a32318 = a32316 & ~a32310;
assign a32320 = a32318 & ~a32308;
assign a32322 = a32320 & ~a32304;
assign a32324 = a32322 & ~a32302;
assign a32326 = a32324 & ~a32300;
assign a32328 = a32326 & ~a32298;
assign a32330 = a32328 & ~a32296;
assign a32332 = a32330 & ~a32294;
assign a32334 = ~a32332 & a31138;
assign a32336 = ~a32334 & ~a32290;
assign a32338 = ~a32336 & ~a32224;
assign a32340 = a32338 & ~a32222;
assign a32342 = a32340 & ~a32102;
assign a32344 = a32342 & ~a32100;
assign a32346 = a32344 & ~a31980;
assign a32348 = a32346 & ~a31978;
assign a32350 = a32348 & ~a31858;
assign a32352 = a32350 & ~a31856;
assign a32354 = a32352 & ~a31736;
assign a32356 = a32354 & ~a31734;
assign a32358 = a32356 & ~a31614;
assign a32360 = a32358 & ~a31612;
assign a32362 = a32360 & ~a31492;
assign a32364 = a32362 & ~a31490;
assign a32366 = a32364 & ~a31370;
assign a32368 = a32366 & ~a31368;
assign a32372 = a9046 & ~l1250;
assign a32374 = ~a9046 & l1250;
assign a32376 = ~a32374 & ~a32372;
assign a32378 = ~a32376 & ~a16190;
assign a32382 = ~a32372 & a9058;
assign a32384 = ~a32382 & ~a18552;
assign a32388 = a32386 & a31160;
assign a32390 = a32388 & a18556;
assign a32392 = a32390 & ~a12354;
assign a32394 = ~a32390 & l1254;
assign a32396 = ~a32394 & ~a32392;
assign a32398 = a25828 & ~a12354;
assign a32400 = ~a25828 & l1258;
assign a32402 = ~a32400 & ~a32398;
assign a32404 = a32390 & ~a12300;
assign a32406 = ~a32390 & l1262;
assign a32408 = ~a32406 & ~a32404;
assign a32410 = a25828 & ~a12300;
assign a32412 = ~a25828 & l1264;
assign a32414 = ~a32412 & ~a32410;
assign a32416 = a32390 & ~a12238;
assign a32418 = ~a32390 & l1268;
assign a32420 = ~a32418 & ~a32416;
assign a32422 = a25828 & ~a12238;
assign a32424 = ~a25828 & l1270;
assign a32426 = ~a32424 & ~a32422;
assign a32428 = a32390 & ~a12178;
assign a32430 = ~a32390 & l1274;
assign a32432 = ~a32430 & ~a32428;
assign a32434 = a25828 & ~a12178;
assign a32436 = ~a25828 & l1276;
assign a32438 = ~a32436 & ~a32434;
assign a32440 = ~a8924 & l946;
assign a32442 = a26574 & ~a23054;
assign a32444 = ~a26574 & l1308;
assign a32446 = ~a32444 & ~a32442;
assign a32448 = ~a32446 & ~l946;
assign a32450 = ~a32448 & ~a32440;
assign a32452 = ~a32450 & ~l886;
assign a32454 = ~a32452 & ~a8908;
assign a32456 = ~a8986 & l946;
assign a32458 = a26574 & ~a23058;
assign a32460 = ~a26574 & ~a11974;
assign a32462 = ~a32460 & ~a32458;
assign a32464 = ~a32462 & ~l946;
assign a32466 = ~a32464 & ~a32456;
assign a32468 = ~a32466 & ~l886;
assign a32472 = ~a8954 & l946;
assign a32474 = a26574 & a11996;
assign a32476 = a26582 & ~a11996;
assign a32478 = ~a32476 & ~a32474;
assign a32480 = ~a32478 & ~l946;
assign a32482 = ~a32480 & ~a32472;
assign a32484 = ~a32482 & ~l886;
assign a32488 = a23666 & ~i370;
assign a32490 = ~l1490 & l890;
assign a32492 = a11964 & ~l890;
assign a32494 = ~a32492 & ~a32490;
assign a32496 = a32494 & ~l884;
assign a32498 = ~a32496 & ~a32488;
assign a32500 = ~a32488 & ~a22752;
assign a32502 = a32500 & ~a32498;
assign a32506 = a26564 & ~i368;
assign a32510 = a32454 & l1308;
assign a32512 = ~a26594 & ~l1000;
assign a32514 = a26594 & l1000;
assign a32516 = ~a32486 & a11996;
assign a32518 = a32486 & ~a11996;
assign a32520 = ~a32470 & a11974;
assign a32522 = a32470 & ~a11974;
assign a32524 = ~a32454 & ~l1308;
assign a32526 = ~a32524 & ~a32522;
assign a32528 = a32526 & ~a32520;
assign a32530 = a32528 & ~a32518;
assign a32532 = a32530 & ~a32516;
assign a32534 = a32532 & ~a32514;
assign a32536 = a32534 & ~a32512;
assign a32540 = l1496 & l886;
assign a32542 = a25350 & ~a21698;
assign a32544 = ~a12540 & ~a12526;
assign a32546 = a32544 & l1498;
assign a32548 = ~a32546 & l1494;
assign a32550 = a32546 & ~l1494;
assign a32552 = ~a32550 & ~a32548;
assign a32554 = a14410 & l1622;
assign a32556 = ~a32554 & ~a15512;
assign a32558 = a32556 & a15510;
assign a32560 = ~a15520 & ~a15516;
assign a32562 = ~a15528 & ~a15524;
assign a32564 = ~a15536 & ~a15532;
assign a32566 = ~a15544 & ~a15540;
assign a32568 = ~a15552 & ~a15548;
assign a32570 = a32568 & a15504;
assign a32572 = a32570 & a32566;
assign a32574 = a32572 & a32564;
assign a32576 = a32574 & a32562;
assign a32578 = a32576 & a32560;
assign a32580 = a32578 & a32558;
assign a32582 = ~a32580 & a14378;
assign a32584 = a14378 & l1542;
assign a32586 = a32584 & a32580;
assign a32588 = ~a32586 & ~l2006;
assign a32590 = ~a32588 & ~a32582;
assign a32594 = a32592 & ~a12526;
assign a32596 = a14410 & l1624;
assign a32598 = ~a32596 & ~a15346;
assign a32600 = a32598 & a15344;
assign a32602 = ~a15354 & ~a15350;
assign a32604 = ~a15362 & ~a15358;
assign a32606 = ~a15370 & ~a15366;
assign a32608 = ~a15378 & ~a15374;
assign a32610 = ~a15386 & ~a15382;
assign a32612 = a32610 & a32608;
assign a32614 = a32612 & a32606;
assign a32616 = a32614 & a32604;
assign a32618 = a32616 & a32602;
assign a32620 = a32618 & a32600;
assign a32622 = a32620 & a15338;
assign a32624 = ~a32622 & a14378;
assign a32626 = a14378 & l1584;
assign a32628 = a32626 & a32622;
assign a32630 = ~a32628 & ~l2008;
assign a32632 = ~a32630 & ~a32624;
assign a32636 = a32634 & a12526;
assign a32638 = ~a32636 & ~a32594;
assign a32640 = ~a32638 & ~a12540;
assign a32642 = a14410 & l1626;
assign a32644 = ~a32642 & ~a15180;
assign a32646 = a32644 & a15178;
assign a32648 = ~a15188 & ~a15184;
assign a32650 = ~a15196 & ~a15192;
assign a32652 = ~a15204 & ~a15200;
assign a32654 = ~a15212 & ~a15208;
assign a32656 = ~a15220 & ~a15216;
assign a32658 = a32656 & a32654;
assign a32660 = a32658 & a32652;
assign a32662 = a32660 & a32650;
assign a32664 = a32662 & a32648;
assign a32666 = a32664 & a32646;
assign a32668 = a32666 & a15172;
assign a32670 = ~a32668 & a14378;
assign a32672 = a14378 & l1586;
assign a32674 = a32672 & a32668;
assign a32676 = ~a32674 & ~l2010;
assign a32678 = ~a32676 & ~a32670;
assign a32682 = a32680 & ~a12526;
assign a32684 = a14410 & l1628;
assign a32686 = ~a32684 & ~a15010;
assign a32688 = a32686 & a15008;
assign a32690 = ~a15018 & ~a15014;
assign a32692 = ~a15026 & ~a15022;
assign a32694 = ~a15034 & ~a15030;
assign a32696 = ~a15042 & ~a15038;
assign a32698 = ~a15050 & ~a15046;
assign a32700 = a32698 & a32696;
assign a32702 = a32700 & a32694;
assign a32704 = a32702 & a32692;
assign a32706 = a32704 & a32690;
assign a32708 = a32706 & a32688;
assign a32710 = a32708 & a15002;
assign a32712 = ~a32710 & a14378;
assign a32714 = a14378 & l1588;
assign a32716 = a32714 & a32710;
assign a32718 = ~a32716 & ~l2012;
assign a32720 = ~a32718 & ~a32712;
assign a32724 = a32722 & a12526;
assign a32726 = ~a32724 & ~a32682;
assign a32728 = ~a32726 & a12540;
assign a32730 = ~a32728 & ~a32640;
assign a32732 = ~a32730 & l1498;
assign a32734 = a14410 & l1630;
assign a32736 = ~a32734 & ~a14842;
assign a32738 = a32736 & a14840;
assign a32740 = ~a14850 & ~a14846;
assign a32742 = ~a14858 & ~a14854;
assign a32744 = ~a14866 & ~a14862;
assign a32746 = ~a14874 & ~a14870;
assign a32748 = ~a14882 & ~a14878;
assign a32750 = a32748 & a32746;
assign a32752 = a32750 & a32744;
assign a32754 = a32752 & a32742;
assign a32756 = a32754 & a32740;
assign a32758 = a32756 & a32738;
assign a32760 = a32758 & a14834;
assign a32762 = ~a32760 & a14378;
assign a32764 = a14378 & l1590;
assign a32766 = a32764 & a32760;
assign a32768 = ~a32766 & ~l2014;
assign a32770 = ~a32768 & ~a32762;
assign a32774 = a32772 & ~a12526;
assign a32776 = a14410 & l1632;
assign a32778 = ~a32776 & ~a14672;
assign a32780 = a32778 & a14670;
assign a32782 = ~a14680 & ~a14676;
assign a32784 = ~a14688 & ~a14684;
assign a32786 = ~a14696 & ~a14692;
assign a32788 = ~a14704 & ~a14700;
assign a32790 = ~a14712 & ~a14708;
assign a32792 = a32790 & a32788;
assign a32794 = a32792 & a32786;
assign a32796 = a32794 & a32784;
assign a32798 = a32796 & a32782;
assign a32800 = a32798 & a32780;
assign a32802 = a32800 & a14664;
assign a32804 = ~a32802 & a14378;
assign a32806 = a14378 & l1592;
assign a32808 = a32806 & a32802;
assign a32810 = ~a32808 & ~l2016;
assign a32812 = ~a32810 & ~a32804;
assign a32816 = a32814 & a12526;
assign a32818 = ~a32816 & ~a32774;
assign a32820 = ~a32818 & ~a12540;
assign a32822 = a14410 & ~a12888;
assign a32824 = ~a32822 & ~a14430;
assign a32826 = a32824 & a14428;
assign a32828 = ~a14450 & ~a14446;
assign a32830 = ~a14470 & ~a14466;
assign a32832 = ~a14490 & ~a14486;
assign a32834 = ~a14510 & ~a14506;
assign a32836 = ~a14530 & ~a14526;
assign a32838 = a32836 & a32834;
assign a32840 = a32838 & a32832;
assign a32842 = a32840 & a32830;
assign a32844 = a32842 & a32828;
assign a32846 = a32844 & a32826;
assign a32848 = a32846 & a14398;
assign a32850 = ~a32848 & a14378;
assign a32852 = a14378 & a12574;
assign a32854 = a32852 & a32848;
assign a32856 = ~a32854 & ~l2018;
assign a32858 = ~a32856 & ~a32850;
assign a32862 = a32860 & ~a12526;
assign a32864 = a14410 & ~a12902;
assign a32866 = ~a32864 & ~a16016;
assign a32868 = a32866 & a16014;
assign a32870 = ~a16024 & ~a16020;
assign a32872 = ~a16032 & ~a16028;
assign a32874 = ~a16040 & ~a16036;
assign a32876 = ~a16048 & ~a16044;
assign a32878 = ~a16056 & ~a16052;
assign a32880 = a32878 & a32876;
assign a32882 = a32880 & a32874;
assign a32884 = a32882 & a32872;
assign a32886 = a32884 & a32870;
assign a32888 = a32886 & a32868;
assign a32890 = a32888 & a16008;
assign a32892 = ~a32890 & a14378;
assign a32894 = a14378 & a12582;
assign a32896 = a32894 & a32890;
assign a32898 = ~l2020 & l890;
assign a32900 = ~a12502 & ~l890;
assign a32902 = ~a32900 & ~a32898;
assign a32904 = ~a32902 & ~a32896;
assign a32906 = ~a32904 & ~a32892;
assign a32910 = a32908 & a12526;
assign a32912 = ~a32910 & ~a32862;
assign a32914 = ~a32912 & a12540;
assign a32916 = ~a32914 & ~a32820;
assign a32918 = ~a32916 & ~l1498;
assign a32920 = ~a32918 & ~a32732;
assign a32922 = ~a32920 & ~l1494;
assign a32924 = a16380 & ~l926;
assign a32926 = a23672 & a11996;
assign a32928 = ~a23672 & i410;
assign a32930 = ~a32928 & ~a32926;
assign a32932 = a23672 & ~l1000;
assign a32934 = ~a23672 & i412;
assign a32936 = ~a32934 & ~a32932;
assign a32938 = a23672 & ~l1308;
assign a32940 = ~a23672 & i414;
assign a32942 = ~a32940 & ~a32938;
assign a32944 = a23672 & a11974;
assign a32946 = ~a23672 & i416;
assign a32948 = ~a32946 & ~a32944;
assign a32950 = ~a32948 & ~a32942;
assign a32952 = a32950 & a32936;
assign a32954 = a32952 & a23672;
assign a32956 = a32954 & a32930;
assign a32958 = a32956 & a32924;
assign a32960 = ~a32958 & ~l1510;
assign a32962 = ~a32960 & ~l886;
assign a32964 = a32962 & ~l948;
assign a32968 = a32966 & ~a12526;
assign a32970 = a32954 & ~a32930;
assign a32972 = a32970 & a32924;
assign a32974 = ~a32972 & ~l1514;
assign a32976 = ~a32974 & ~l948;
assign a32980 = a32978 & a12526;
assign a32982 = ~a32980 & ~a32968;
assign a32984 = ~a32982 & l1494;
assign a32986 = a32932 & a32930;
assign a32988 = a32986 & a32948;
assign a32990 = a32988 & a32942;
assign a32992 = a32990 & a32924;
assign a32994 = ~a32992 & ~l1542;
assign a32996 = ~a32994 & ~l948;
assign a33000 = a32998 & ~a12526;
assign a33002 = a32932 & ~a32930;
assign a33004 = a33002 & a32948;
assign a33006 = a33004 & a32942;
assign a33008 = a33006 & a32924;
assign a33010 = ~a33008 & ~l1584;
assign a33012 = ~a33010 & ~l948;
assign a33016 = a33014 & a12526;
assign a33018 = ~a33016 & ~a33000;
assign a33020 = ~a33018 & ~a12540;
assign a33022 = a32986 & ~a32948;
assign a33024 = a33022 & a32942;
assign a33026 = a33024 & a32924;
assign a33028 = ~a33026 & ~l1586;
assign a33030 = ~a33028 & ~l948;
assign a33034 = a33032 & ~a12526;
assign a33036 = a33002 & ~a32948;
assign a33038 = a33036 & a32942;
assign a33040 = a33038 & a32924;
assign a33042 = ~a33040 & ~l1588;
assign a33044 = ~a33042 & ~l948;
assign a33048 = a33046 & a12526;
assign a33050 = ~a33048 & ~a33034;
assign a33052 = ~a33050 & a12540;
assign a33054 = ~a33052 & ~a33020;
assign a33056 = ~a33054 & l1498;
assign a33058 = a32988 & ~a32942;
assign a33060 = a33058 & a32924;
assign a33062 = ~a33060 & ~l1590;
assign a33064 = ~a33062 & ~l948;
assign a33068 = a33066 & ~a12526;
assign a33070 = a33004 & ~a32942;
assign a33072 = a33070 & a32924;
assign a33074 = ~a33072 & ~l1592;
assign a33076 = ~a33074 & ~l948;
assign a33080 = a33078 & a12526;
assign a33082 = ~a33080 & ~a33068;
assign a33084 = ~a33082 & ~a12540;
assign a33086 = a33022 & ~a32942;
assign a33088 = a33086 & a32924;
assign a33090 = ~a33088 & ~a12574;
assign a33092 = ~a33090 & ~l948;
assign a33096 = a33094 & ~a12526;
assign a33098 = a33036 & ~a32942;
assign a33100 = a33098 & a32924;
assign a33102 = ~a33100 & ~a12582;
assign a33104 = ~a33102 & ~l948;
assign a33108 = a33106 & a12526;
assign a33110 = ~a33108 & ~a33096;
assign a33112 = ~a33110 & a12540;
assign a33114 = ~a33112 & ~a33084;
assign a33116 = ~a33114 & ~l1498;
assign a33118 = ~a33116 & ~a33056;
assign a33120 = ~a33118 & ~l1494;
assign a33122 = ~a33120 & ~a32984;
assign a33124 = a14410 & l1618;
assign a33126 = ~a15852 & ~a15848;
assign a33128 = a33126 & ~a15856;
assign a33130 = a33128 & ~a15860;
assign a33132 = a33130 & ~a15864;
assign a33134 = a33132 & ~a15868;
assign a33136 = a33134 & ~a15872;
assign a33138 = a33136 & ~a15876;
assign a33140 = a33138 & ~a15880;
assign a33142 = a33140 & ~a15884;
assign a33144 = a33142 & ~a15888;
assign a33146 = a33144 & ~a33124;
assign a33148 = a33146 & a15840;
assign a33150 = a33148 & a15846;
assign a33152 = a33150 & a15834;
assign a33154 = ~a33152 & ~l2022;
assign a33158 = a33156 & ~a12526;
assign a33160 = a14410 & l1620;
assign a33162 = ~a33160 & ~a15678;
assign a33164 = a33162 & a15676;
assign a33166 = ~a15686 & ~a15682;
assign a33168 = ~a15694 & ~a15690;
assign a33170 = ~a15702 & ~a15698;
assign a33172 = ~a15710 & ~a15706;
assign a33174 = ~a15718 & ~a15714;
assign a33176 = a33174 & a15670;
assign a33178 = a33176 & a33172;
assign a33180 = a33178 & a33170;
assign a33182 = a33180 & a33168;
assign a33184 = a33182 & a33166;
assign a33186 = a33184 & a33164;
assign a33188 = ~a33186 & a14378;
assign a33190 = a14378 & l1514;
assign a33192 = a33190 & a33186;
assign a33194 = ~a33192 & ~l2024;
assign a33196 = ~a33194 & ~a33188;
assign a33200 = a33198 & a12526;
assign a33202 = ~a33200 & ~a33158;
assign a33204 = ~a33202 & l1494;
assign a33206 = ~a33204 & ~a33122;
assign a33208 = a33206 & ~a32922;
assign a33210 = ~a12526 & a11996;
assign a33212 = a12526 & ~a11996;
assign a33214 = ~a12540 & a11974;
assign a33216 = a12540 & ~a11974;
assign a33218 = l1498 & ~l1308;
assign a33220 = ~l1498 & l1308;
assign a33222 = l1494 & ~l1000;
assign a33224 = ~l1494 & l1000;
assign a33226 = ~a33224 & ~a33222;
assign a33228 = a33226 & ~a33220;
assign a33230 = a33228 & ~a33218;
assign a33232 = a33230 & ~a33216;
assign a33234 = a33232 & ~a33214;
assign a33236 = a33234 & ~a33212;
assign a33238 = a33236 & ~a33210;
assign a33240 = ~a33238 & ~a33208;
assign a33242 = a12540 & ~a12526;
assign a33244 = a33242 & a12606;
assign a33246 = a12526 & ~l1550;
assign a33248 = ~a12526 & l1550;
assign a33250 = ~a12540 & a12526;
assign a33252 = ~a33250 & ~a33242;
assign a33254 = ~a33252 & ~l1552;
assign a33256 = a33252 & l1552;
assign a33258 = ~a32544 & l1498;
assign a33260 = a32544 & ~l1498;
assign a33262 = ~a33260 & ~a33258;
assign a33264 = ~a33262 & ~l1556;
assign a33266 = a33262 & l1556;
assign a33268 = ~a32552 & ~l1554;
assign a33270 = a32552 & l1554;
assign a33272 = ~a33270 & ~a33268;
assign a33274 = a33272 & ~a33266;
assign a33276 = a33274 & ~a33264;
assign a33278 = a33276 & ~a33256;
assign a33280 = a33278 & ~a33254;
assign a33282 = a33280 & ~a33248;
assign a33284 = a33282 & ~a33246;
assign a33286 = a12526 & l968;
assign a33288 = ~a12526 & l970;
assign a33290 = ~a33288 & ~a33286;
assign a33292 = ~a33290 & ~a32552;
assign a33294 = a12526 & l966;
assign a33296 = ~a12526 & l964;
assign a33298 = ~a33296 & ~a33294;
assign a33300 = ~a33298 & ~a33252;
assign a33302 = a12526 & l962;
assign a33304 = ~a12526 & l960;
assign a33306 = ~a33304 & ~a33302;
assign a33308 = ~a33306 & a33252;
assign a33310 = ~a33308 & ~a33300;
assign a33312 = ~a33310 & ~a33262;
assign a33314 = a12526 & a5606;
assign a33316 = ~a12526 & a5600;
assign a33318 = ~a33316 & ~a33314;
assign a33320 = ~a33318 & ~a33252;
assign a33322 = a12526 & a5594;
assign a33324 = ~a12526 & a5568;
assign a33326 = ~a33324 & ~a33322;
assign a33328 = ~a33326 & a33252;
assign a33330 = ~a33328 & ~a33320;
assign a33332 = ~a33330 & a33262;
assign a33334 = ~a33332 & ~a33312;
assign a33336 = ~a33334 & a32552;
assign a33338 = ~a33336 & ~a33292;
assign a33340 = ~a33338 & ~a33284;
assign a33342 = a33340 & ~a33244;
assign a33344 = a33342 & a33240;
assign a33346 = a33344 & ~a32552;
assign a33348 = ~l1552 & ~l1550;
assign a33350 = a33348 & ~l1554;
assign a33352 = a33350 & ~l1556;
assign a33354 = ~a33352 & a5568;
assign a33356 = a33354 & a33240;
assign a33358 = ~a33356 & ~a33344;
assign a33360 = a33358 & l1494;
assign a33362 = ~a33360 & ~a33346;
assign a33364 = ~a33362 & ~a25350;
assign a33366 = ~a33364 & ~a32542;
assign a33368 = ~a33366 & ~l948;
assign a33370 = ~a33368 & ~a8872;
assign a33372 = ~a33370 & ~l886;
assign a33374 = ~a33372 & ~a32540;
assign a33376 = a5360 & ~a2512;
assign a33378 = ~a5360 & l1496;
assign a33380 = ~a33378 & ~a33376;
assign a33382 = l1500 & l886;
assign a33384 = a25350 & ~a21682;
assign a33386 = a33344 & ~a33262;
assign a33388 = a33358 & l1498;
assign a33390 = ~a33388 & ~a33386;
assign a33392 = ~a33390 & ~a25350;
assign a33394 = ~a33392 & ~a33384;
assign a33396 = ~a33394 & ~l948;
assign a33398 = ~a33396 & ~a8926;
assign a33400 = ~a33398 & ~l886;
assign a33402 = ~a33400 & ~a33382;
assign a33404 = a5360 & ~a2532;
assign a33406 = ~a5360 & l1500;
assign a33408 = ~a33406 & ~a33404;
assign a33410 = l1504 & l886;
assign a33412 = a25350 & ~a21676;
assign a33414 = a33344 & a12526;
assign a33416 = a33358 & ~a12526;
assign a33418 = ~a33416 & ~a33414;
assign a33420 = ~a33418 & ~a25350;
assign a33422 = ~a33420 & ~a33412;
assign a33424 = ~a33422 & ~l948;
assign a33426 = ~a33424 & ~a8956;
assign a33428 = ~a33426 & ~l886;
assign a33432 = a5360 & ~l880;
assign a33434 = ~a5360 & l1504;
assign a33436 = ~a33434 & ~a33432;
assign a33438 = l1508 & l886;
assign a33440 = a25350 & ~a21688;
assign a33442 = a33344 & ~a33252;
assign a33444 = a33358 & ~a12540;
assign a33446 = ~a33444 & ~a33442;
assign a33448 = ~a33446 & ~a25350;
assign a33450 = ~a33448 & ~a33440;
assign a33452 = ~a33450 & ~l948;
assign a33454 = ~a33452 & ~a8988;
assign a33456 = ~a33454 & ~l886;
assign a33460 = a5360 & ~a2748;
assign a33462 = ~a5360 & l1508;
assign a33464 = ~a33462 & ~a33460;
assign a33466 = ~l946 & ~l944;
assign a33468 = a33466 & ~l948;
assign a33470 = a32292 & l1524;
assign a33472 = a32230 & l1988;
assign a33474 = a31348 & l1990;
assign a33476 = a32238 & l1992;
assign a33478 = a32244 & l1994;
assign a33480 = a32248 & l1996;
assign a33482 = a32306 & l1998;
assign a33484 = a32258 & l2000;
assign a33486 = a32264 & l2002;
assign a33488 = a32268 & l2004;
assign a33490 = ~a33488 & ~a33486;
assign a33492 = a33490 & ~a33484;
assign a33494 = a33492 & ~a33482;
assign a33496 = a33494 & ~a33480;
assign a33498 = a33496 & ~a33478;
assign a33500 = a33498 & ~a33476;
assign a33502 = a33500 & ~a33474;
assign a33504 = a33502 & ~a33472;
assign a33506 = a33504 & ~a33470;
assign a33508 = a2740 & ~l1156;
assign a33510 = a33508 & l1244;
assign a33512 = a33510 & a19878;
assign a33514 = ~a33512 & l1524;
assign a33516 = ~l1528 & l890;
assign a33518 = i418 & ~i92;
assign a33520 = ~a33518 & ~l890;
assign a33522 = ~a33520 & ~a33516;
assign a33524 = a33522 & a33512;
assign a33526 = ~a33524 & ~a33514;
assign a33528 = a2748 & l880;
assign a33530 = a33528 & a2532;
assign a33532 = a33530 & a2512;
assign a33534 = a33532 & ~l1532;
assign a33536 = ~a33532 & l1532;
assign a33538 = ~a33536 & ~a33534;
assign a33540 = ~a33538 & l886;
assign a33542 = ~a23774 & l948;
assign a33544 = a8874 & l1530;
assign a33546 = a8888 & l1246;
assign a33548 = ~a33546 & l1530;
assign a33550 = a33546 & ~l1530;
assign a33552 = ~a33550 & ~a33548;
assign a33554 = ~a33552 & ~a8882;
assign a33556 = a8882 & ~l1530;
assign a33558 = ~a33556 & ~a33554;
assign a33560 = ~a33558 & ~a8874;
assign a33562 = ~a33560 & ~a33544;
assign a33564 = ~a33562 & ~l948;
assign a33566 = ~a33564 & ~a33542;
assign a33568 = ~a33566 & ~l886;
assign a33570 = ~a33568 & ~a33540;
assign a33572 = a26686 & l1524;
assign a33574 = a26740 & l1988;
assign a33576 = a26730 & ~a2504;
assign a33578 = a33576 & l1990;
assign a33580 = a2504 & l1992;
assign a33582 = a33580 & a26730;
assign a33584 = ~a2504 & l1994;
assign a33586 = a33584 & a26642;
assign a33588 = a26644 & l1996;
assign a33590 = ~a2752 & ~a2504;
assign a33592 = a33590 & a2536;
assign a33594 = a33592 & l1998;
assign a33596 = a33594 & a2516;
assign a33598 = a26768 & l2000;
assign a33600 = a33598 & a2536;
assign a33602 = a26758 & l2002;
assign a33604 = a33602 & a2536;
assign a33606 = a26600 & l2004;
assign a33608 = ~a33606 & ~a33604;
assign a33610 = a33608 & ~a33600;
assign a33612 = a33610 & ~a33596;
assign a33614 = a33612 & ~a33588;
assign a33616 = a33614 & ~a33586;
assign a33618 = a33616 & ~a33582;
assign a33620 = a33618 & ~a33578;
assign a33622 = a33620 & ~a33574;
assign a33624 = a33622 & ~a33572;
assign a33626 = ~a2536 & ~a2504;
assign a33628 = ~a26738 & ~a26728;
assign a33630 = a33628 & ~a33626;
assign a33632 = ~a33630 & l1010;
assign a33634 = a26608 & ~a2536;
assign a33636 = ~a33634 & ~a33632;
assign a33638 = a2504 & l1010;
assign a33640 = a26608 & ~a2504;
assign a33642 = ~a33640 & ~a33638;
assign a33644 = ~a33590 & ~a26738;
assign a33646 = a33644 & ~a26644;
assign a33648 = ~a33646 & l1010;
assign a33650 = a26608 & ~a2752;
assign a33652 = ~a33650 & ~a33648;
assign a33654 = ~a26872 & l1010;
assign a33656 = ~a26924 & a26608;
assign a33658 = a26830 & a2752;
assign a33660 = a26600 & ~a18872;
assign a33662 = ~a33660 & ~a33658;
assign a33664 = a26706 & a2504;
assign a33666 = a33664 & a26888;
assign a33668 = ~a33666 & a33662;
assign a33670 = a33592 & a26840;
assign a33672 = ~a33670 & a33668;
assign a33674 = a26644 & l1792;
assign a33676 = ~a33674 & a33672;
assign a33678 = a26856 & a26650;
assign a33680 = ~a33678 & a33676;
assign a33682 = a26908 & a2504;
assign a33684 = ~a33682 & a33680;
assign a33686 = a33576 & l1798;
assign a33688 = ~a33686 & a33684;
assign a33690 = a26920 & a2504;
assign a33692 = ~a33690 & a33688;
assign a33694 = a26814 & ~a2516;
assign a33696 = ~a33694 & a33692;
assign a33698 = ~a33696 & ~a2780;
assign a33700 = ~a33698 & ~a33656;
assign a33702 = a33700 & ~a33654;
assign a33704 = a33702 & ~a18850;
assign a33706 = ~a27034 & l1010;
assign a33708 = ~a27086 & a26608;
assign a33710 = a26992 & a2752;
assign a33712 = a26600 & ~a18946;
assign a33714 = ~a33712 & ~a33710;
assign a33716 = a33664 & a27050;
assign a33718 = ~a33716 & a33714;
assign a33720 = a33592 & a27002;
assign a33722 = ~a33720 & a33718;
assign a33724 = a26644 & l1814;
assign a33726 = ~a33724 & a33722;
assign a33728 = a27018 & a26650;
assign a33730 = ~a33728 & a33726;
assign a33732 = a27070 & a2504;
assign a33734 = ~a33732 & a33730;
assign a33736 = a33576 & l1820;
assign a33738 = ~a33736 & a33734;
assign a33740 = a27082 & a2504;
assign a33742 = ~a33740 & a33738;
assign a33744 = a26976 & ~a2516;
assign a33746 = ~a33744 & a33742;
assign a33748 = ~a33746 & ~a2780;
assign a33750 = ~a33748 & ~a33708;
assign a33752 = a33750 & ~a33706;
assign a33754 = a33752 & ~a18924;
assign a33756 = ~a33754 & ~a33704;
assign a33758 = ~a33752 & a18924;
assign a33760 = ~a33758 & ~a33756;
assign a33762 = ~a27204 & l1010;
assign a33764 = ~a27256 & a26608;
assign a33766 = a27160 & a2752;
assign a33768 = a26600 & ~a19026;
assign a33770 = ~a33768 & ~a33766;
assign a33772 = a33664 & a27220;
assign a33774 = ~a33772 & a33770;
assign a33776 = a33592 & a27170;
assign a33778 = ~a33776 & a33774;
assign a33780 = a26644 & l1836;
assign a33782 = ~a33780 & a33778;
assign a33784 = a27186 & a26650;
assign a33786 = ~a33784 & a33782;
assign a33788 = a27240 & a2504;
assign a33790 = ~a33788 & a33786;
assign a33792 = a33576 & l1842;
assign a33794 = ~a33792 & a33790;
assign a33796 = a27252 & a2504;
assign a33798 = ~a33796 & a33794;
assign a33800 = a27144 & ~a2516;
assign a33802 = ~a33800 & a33798;
assign a33804 = ~a33802 & ~a2780;
assign a33806 = ~a33804 & ~a33764;
assign a33808 = a33806 & ~a33762;
assign a33810 = a33808 & ~a19004;
assign a33812 = ~a33810 & ~a33760;
assign a33814 = ~a33808 & a19004;
assign a33816 = ~a33814 & ~a33812;
assign a33818 = ~a27374 & l1010;
assign a33820 = ~a27426 & a26608;
assign a33822 = a27330 & a2752;
assign a33824 = a26600 & ~a19108;
assign a33826 = ~a33824 & ~a33822;
assign a33828 = a33664 & a27390;
assign a33830 = ~a33828 & a33826;
assign a33832 = a33592 & a27340;
assign a33834 = ~a33832 & a33830;
assign a33836 = a26644 & l1858;
assign a33838 = ~a33836 & a33834;
assign a33840 = a27356 & a26650;
assign a33842 = ~a33840 & a33838;
assign a33844 = a27410 & a2504;
assign a33846 = ~a33844 & a33842;
assign a33848 = a33576 & l1864;
assign a33850 = ~a33848 & a33846;
assign a33852 = a27422 & a2504;
assign a33854 = ~a33852 & a33850;
assign a33856 = a27314 & ~a2516;
assign a33858 = ~a33856 & a33854;
assign a33860 = ~a33858 & ~a2780;
assign a33862 = ~a33860 & ~a33820;
assign a33864 = a33862 & ~a33818;
assign a33866 = a33864 & ~a19086;
assign a33868 = ~a33866 & ~a33816;
assign a33870 = ~a33864 & a19086;
assign a33872 = ~a33870 & ~a33868;
assign a33874 = ~a27544 & l1010;
assign a33876 = ~a27596 & a26608;
assign a33878 = a27500 & a2752;
assign a33880 = a26600 & ~a19190;
assign a33882 = ~a33880 & ~a33878;
assign a33884 = a33664 & a27560;
assign a33886 = ~a33884 & a33882;
assign a33888 = a33592 & a27510;
assign a33890 = ~a33888 & a33886;
assign a33892 = a26644 & l1880;
assign a33894 = ~a33892 & a33890;
assign a33896 = a27526 & a26650;
assign a33898 = ~a33896 & a33894;
assign a33900 = a27580 & a2504;
assign a33902 = ~a33900 & a33898;
assign a33904 = a33576 & l1886;
assign a33906 = ~a33904 & a33902;
assign a33908 = a27592 & a2504;
assign a33910 = ~a33908 & a33906;
assign a33912 = a27484 & ~a2516;
assign a33914 = ~a33912 & a33910;
assign a33916 = ~a33914 & ~a2780;
assign a33918 = ~a33916 & ~a33876;
assign a33920 = a33918 & ~a33874;
assign a33922 = a33920 & ~a19168;
assign a33924 = ~a33922 & ~a33872;
assign a33926 = ~a33920 & a19168;
assign a33928 = ~a33926 & ~a33924;
assign a33930 = ~a27714 & l1010;
assign a33932 = ~a27766 & a26608;
assign a33934 = a27670 & a2752;
assign a33936 = a26600 & ~a19272;
assign a33938 = ~a33936 & ~a33934;
assign a33940 = a33664 & a27730;
assign a33942 = ~a33940 & a33938;
assign a33944 = a33592 & a27680;
assign a33946 = ~a33944 & a33942;
assign a33948 = a26644 & l1902;
assign a33950 = ~a33948 & a33946;
assign a33952 = a27696 & a26650;
assign a33954 = ~a33952 & a33950;
assign a33956 = a27750 & a2504;
assign a33958 = ~a33956 & a33954;
assign a33960 = a33576 & l1908;
assign a33962 = ~a33960 & a33958;
assign a33964 = a27762 & a2504;
assign a33966 = ~a33964 & a33962;
assign a33968 = a27654 & ~a2516;
assign a33970 = ~a33968 & a33966;
assign a33972 = ~a33970 & ~a2780;
assign a33974 = ~a33972 & ~a33932;
assign a33976 = a33974 & ~a33930;
assign a33978 = a33976 & ~a19250;
assign a33980 = ~a33978 & ~a33928;
assign a33982 = ~a33976 & a19250;
assign a33984 = ~a33982 & ~a33980;
assign a33986 = ~a27884 & l1010;
assign a33988 = ~a27936 & a26608;
assign a33990 = a27840 & a2752;
assign a33992 = a26600 & ~a19348;
assign a33994 = ~a33992 & ~a33990;
assign a33996 = a33664 & a27900;
assign a33998 = ~a33996 & a33994;
assign a34000 = a33592 & a27850;
assign a34002 = ~a34000 & a33998;
assign a34004 = a26644 & l1924;
assign a34006 = ~a34004 & a34002;
assign a34008 = a27866 & a26650;
assign a34010 = ~a34008 & a34006;
assign a34012 = a27920 & a2504;
assign a34014 = ~a34012 & a34010;
assign a34016 = a33576 & l1930;
assign a34018 = ~a34016 & a34014;
assign a34020 = a27932 & a2504;
assign a34022 = ~a34020 & a34018;
assign a34024 = a27824 & ~a2516;
assign a34026 = ~a34024 & a34022;
assign a34028 = ~a34026 & ~a2780;
assign a34030 = ~a34028 & ~a33988;
assign a34032 = a34030 & ~a33986;
assign a34034 = a34032 & ~a19332;
assign a34036 = ~a34034 & ~a33984;
assign a34038 = ~a34032 & a19332;
assign a34040 = ~a26690 & l1010;
assign a34042 = ~a26752 & a26608;
assign a34044 = a26636 & a2752;
assign a34046 = a26600 & l1938;
assign a34048 = ~a34046 & ~a34044;
assign a34050 = a33664 & a26708;
assign a34052 = ~a34050 & a34048;
assign a34054 = a33592 & a26652;
assign a34056 = ~a34054 & a34052;
assign a34058 = a26644 & l1946;
assign a34060 = ~a34058 & a34056;
assign a34062 = a26670 & a26650;
assign a34064 = ~a34062 & a34060;
assign a34066 = a26732 & a2504;
assign a34068 = ~a34066 & a34064;
assign a34070 = a33576 & l1952;
assign a34072 = ~a34070 & a34068;
assign a34074 = a26748 & a2504;
assign a34076 = ~a34074 & a34072;
assign a34078 = a26616 & ~a2516;
assign a34080 = ~a34078 & a34076;
assign a34082 = ~a34080 & ~a2780;
assign a34084 = ~a34082 & ~a34042;
assign a34086 = a34084 & ~a34040;
assign a34088 = a34086 & ~a19408;
assign a34090 = ~a34086 & a19408;
assign a34092 = ~a34090 & ~a34088;
assign a34094 = ~a34092 & ~a34038;
assign a34096 = a34094 & ~a34036;
assign a34098 = ~a33702 & a18850;
assign a34100 = ~a34098 & ~a33758;
assign a34102 = ~a34100 & ~a33754;
assign a34104 = ~a34102 & ~a33814;
assign a34106 = ~a34104 & ~a33810;
assign a34108 = ~a34106 & ~a33870;
assign a34110 = ~a34108 & ~a33866;
assign a34112 = ~a34110 & ~a33926;
assign a34114 = ~a34112 & ~a33922;
assign a34116 = ~a34114 & ~a33982;
assign a34118 = ~a34116 & ~a33978;
assign a34120 = ~a34118 & ~a34038;
assign a34122 = ~a34120 & ~a34034;
assign a34124 = a34122 & a34092;
assign a34126 = ~a28138 & l1010;
assign a34128 = a28090 & ~a2516;
assign a34130 = a28080 & a2504;
assign a34132 = a33576 & l1986;
assign a34134 = a28066 & a2504;
assign a34136 = a28058 & a26650;
assign a34138 = a26644 & l1980;
assign a34140 = a33592 & a28112;
assign a34142 = a33664 & a28040;
assign a34144 = a28102 & a2752;
assign a34146 = a26600 & a18596;
assign a34148 = ~a34146 & ~a34144;
assign a34150 = a34148 & ~a34142;
assign a34152 = a34150 & ~a34140;
assign a34154 = a34152 & ~a34138;
assign a34156 = a34154 & ~a34136;
assign a34158 = a34156 & ~a34134;
assign a34160 = a34158 & ~a34132;
assign a34162 = a34160 & ~a34130;
assign a34164 = a34162 & ~a34128;
assign a34166 = ~a34164 & ~a2780;
assign a34168 = ~a28084 & a26608;
assign a34170 = ~a34168 & ~a34166;
assign a34172 = a34170 & ~a34126;
assign a34174 = ~a34172 & ~a34124;
assign a34178 = l1504 & l884;
assign a34180 = ~l1552 & l1550;
assign a34182 = a34180 & l1554;
assign a34184 = a34182 & ~l1556;
assign a34186 = l1550 & l966;
assign a34188 = ~l1550 & l964;
assign a34190 = ~a34188 & ~a34186;
assign a34192 = ~a34190 & l1552;
assign a34194 = l1550 & l962;
assign a34196 = ~l1550 & l960;
assign a34198 = ~a34196 & ~a34194;
assign a34200 = ~a34198 & ~l1552;
assign a34202 = ~a34200 & ~a34192;
assign a34204 = ~a34202 & l1556;
assign a34206 = a5606 & l1550;
assign a34208 = a5600 & ~l1550;
assign a34210 = ~a34208 & ~a34206;
assign a34212 = ~a34210 & l1552;
assign a34214 = a5594 & l1550;
assign a34216 = a5568 & ~l1550;
assign a34218 = ~a34216 & ~a34214;
assign a34220 = ~a34218 & ~l1552;
assign a34222 = ~a34220 & ~a34212;
assign a34224 = ~a34222 & ~l1556;
assign a34226 = ~a34224 & ~a34204;
assign a34228 = ~a34226 & ~l1554;
assign a34230 = l1550 & l968;
assign a34232 = ~l1550 & l970;
assign a34234 = ~a34232 & ~a34230;
assign a34236 = ~a34234 & l1554;
assign a34238 = ~a34236 & ~a5624;
assign a34240 = a34238 & ~a34228;
assign a34242 = a34240 & ~a34184;
assign a34244 = a34242 & ~l1550;
assign a34246 = ~a34240 & l1550;
assign a34248 = ~a34246 & ~a34244;
assign a34250 = ~a34248 & ~l884;
assign a34252 = ~a34250 & ~a34178;
assign a34254 = l1508 & l884;
assign a34256 = l1552 & ~l1550;
assign a34258 = ~a34256 & ~a34180;
assign a34260 = ~a34258 & a34242;
assign a34262 = ~a34242 & l1552;
assign a34264 = ~a34262 & ~a34260;
assign a34266 = ~a34264 & ~l884;
assign a34268 = ~a34266 & ~a34254;
assign a34270 = l1496 & l884;
assign a34272 = l1552 & l1550;
assign a34274 = a34272 & l1556;
assign a34276 = ~a34274 & l1554;
assign a34278 = a34274 & ~l1554;
assign a34280 = ~a34278 & ~a34276;
assign a34282 = ~a34280 & a34242;
assign a34284 = ~a34240 & l1554;
assign a34286 = ~a34284 & ~a34282;
assign a34288 = ~a34286 & ~l884;
assign a34290 = ~a34288 & ~a34270;
assign a34292 = l1500 & l884;
assign a34294 = ~a34272 & l1556;
assign a34296 = a34272 & ~l1556;
assign a34298 = ~a34296 & ~a34294;
assign a34300 = ~a34298 & a34242;
assign a34302 = ~a34242 & l1556;
assign a34304 = ~a34302 & ~a34300;
assign a34306 = ~a34304 & ~l884;
assign a34308 = ~a34306 & ~a34292;
assign a34310 = ~a23748 & l948;
assign a34312 = ~a25108 & ~a23748;
assign a34314 = ~a34312 & a34310;
assign a34316 = ~a21692 & l1558;
assign a34318 = a23748 & l948;
assign a34320 = ~a34318 & ~a21700;
assign a34322 = a34320 & ~a34316;
assign a34324 = ~a34322 & ~a34310;
assign a34326 = ~a34324 & ~a34314;
assign a34328 = a34310 & a8954;
assign a34330 = ~a21692 & ~a14546;
assign a34332 = ~a34318 & ~a21818;
assign a34334 = a34332 & ~a34330;
assign a34336 = ~a34334 & ~a34310;
assign a34340 = ~a24458 & ~a23746;
assign a34342 = ~a34340 & a34310;
assign a34344 = ~a21692 & l1566;
assign a34346 = ~a34344 & ~a21728;
assign a34348 = ~a34346 & ~l948;
assign a34350 = ~a34348 & ~a34342;
assign a34352 = ~a24196 & ~a23744;
assign a34354 = ~a34352 & a34310;
assign a34356 = ~a21692 & ~a14552;
assign a34358 = ~a34356 & ~a21788;
assign a34360 = ~a34358 & ~l948;
assign a34364 = a23672 & ~l998;
assign a34366 = ~a23672 & i424;
assign a34368 = ~a34366 & ~a34364;
assign a34370 = a34368 & a32956;
assign a34372 = ~a32956 & l1598;
assign a34374 = ~a34372 & ~a34370;
assign a34376 = a34368 & a32970;
assign a34378 = ~a32970 & l1600;
assign a34380 = ~a34378 & ~a34376;
assign a34382 = a34368 & a32990;
assign a34384 = ~a32990 & l1602;
assign a34386 = ~a34384 & ~a34382;
assign a34388 = a34368 & a33006;
assign a34390 = ~a33006 & l1604;
assign a34392 = ~a34390 & ~a34388;
assign a34394 = a34368 & a33024;
assign a34396 = ~a33024 & l1606;
assign a34398 = ~a34396 & ~a34394;
assign a34400 = a34368 & a33038;
assign a34402 = ~a33038 & l1608;
assign a34404 = ~a34402 & ~a34400;
assign a34406 = a34368 & a33058;
assign a34408 = ~a33058 & l1610;
assign a34410 = ~a34408 & ~a34406;
assign a34412 = a34368 & a33070;
assign a34414 = ~a33070 & l1612;
assign a34416 = ~a34414 & ~a34412;
assign a34418 = a34368 & a33086;
assign a34420 = ~a33086 & l1614;
assign a34422 = ~a34420 & ~a34418;
assign a34424 = a34368 & a33098;
assign a34426 = ~a33098 & l1616;
assign a34428 = ~a34426 & ~a34424;
assign a34430 = a23672 & ~a12836;
assign a34432 = ~a23672 & i426;
assign a34434 = ~a34432 & ~a34430;
assign a34436 = a34434 & a32956;
assign a34438 = ~a32956 & l1618;
assign a34440 = ~a34438 & ~a34436;
assign a34442 = a34434 & a32970;
assign a34444 = ~a32970 & l1620;
assign a34446 = ~a34444 & ~a34442;
assign a34448 = a34434 & a32990;
assign a34450 = ~a32990 & l1622;
assign a34452 = ~a34450 & ~a34448;
assign a34454 = a34434 & a33006;
assign a34456 = ~a33006 & l1624;
assign a34458 = ~a34456 & ~a34454;
assign a34460 = a34434 & a33024;
assign a34462 = ~a33024 & l1626;
assign a34464 = ~a34462 & ~a34460;
assign a34466 = a34434 & a33038;
assign a34468 = ~a33038 & l1628;
assign a34470 = ~a34468 & ~a34466;
assign a34472 = a34434 & a33058;
assign a34474 = ~a33058 & l1630;
assign a34476 = ~a34474 & ~a34472;
assign a34478 = a34434 & a33070;
assign a34480 = ~a33070 & l1632;
assign a34482 = ~a34480 & ~a34478;
assign a34484 = a34434 & a33086;
assign a34486 = ~a33086 & ~a12888;
assign a34490 = a34434 & a33098;
assign a34492 = ~a33098 & ~a12902;
assign a34496 = a23672 & ~a13020;
assign a34498 = ~a23672 & i430;
assign a34500 = ~a34498 & ~a34496;
assign a34502 = a34500 & a32956;
assign a34504 = ~a32956 & l1638;
assign a34506 = ~a34504 & ~a34502;
assign a34508 = a34500 & a32970;
assign a34510 = ~a32970 & l1640;
assign a34512 = ~a34510 & ~a34508;
assign a34514 = a34500 & a32990;
assign a34516 = ~a32990 & l1642;
assign a34518 = ~a34516 & ~a34514;
assign a34520 = a34500 & a33006;
assign a34522 = ~a33006 & l1644;
assign a34524 = ~a34522 & ~a34520;
assign a34526 = a34500 & a33024;
assign a34528 = ~a33024 & l1646;
assign a34530 = ~a34528 & ~a34526;
assign a34532 = a34500 & a33038;
assign a34534 = ~a33038 & l1648;
assign a34536 = ~a34534 & ~a34532;
assign a34538 = a34500 & a33058;
assign a34540 = ~a33058 & l1650;
assign a34542 = ~a34540 & ~a34538;
assign a34544 = a34500 & a33070;
assign a34546 = ~a33070 & l1652;
assign a34548 = ~a34546 & ~a34544;
assign a34550 = a34500 & a33086;
assign a34552 = ~a33086 & ~a13072;
assign a34556 = a34500 & a33098;
assign a34558 = ~a33098 & ~a13086;
assign a34562 = a23672 & ~a13210;
assign a34564 = ~a23672 & i434;
assign a34566 = ~a34564 & ~a34562;
assign a34568 = a34566 & a32956;
assign a34570 = ~a32956 & l1658;
assign a34572 = ~a34570 & ~a34568;
assign a34574 = a34566 & a32970;
assign a34576 = ~a32970 & l1660;
assign a34578 = ~a34576 & ~a34574;
assign a34580 = a34566 & a32990;
assign a34582 = ~a32990 & l1662;
assign a34584 = ~a34582 & ~a34580;
assign a34586 = a34566 & a33006;
assign a34588 = ~a33006 & l1664;
assign a34590 = ~a34588 & ~a34586;
assign a34592 = a34566 & a33024;
assign a34594 = ~a33024 & l1666;
assign a34596 = ~a34594 & ~a34592;
assign a34598 = a34566 & a33038;
assign a34600 = ~a33038 & l1668;
assign a34602 = ~a34600 & ~a34598;
assign a34604 = a34566 & a33058;
assign a34606 = ~a33058 & l1670;
assign a34608 = ~a34606 & ~a34604;
assign a34610 = a34566 & a33070;
assign a34612 = ~a33070 & l1672;
assign a34614 = ~a34612 & ~a34610;
assign a34616 = a34566 & a33086;
assign a34618 = ~a33086 & ~a13262;
assign a34622 = a34566 & a33098;
assign a34624 = ~a33098 & ~a13276;
assign a34628 = a23672 & ~a13400;
assign a34630 = ~a23672 & i438;
assign a34632 = ~a34630 & ~a34628;
assign a34634 = a34632 & a32956;
assign a34636 = ~a32956 & l1678;
assign a34638 = ~a34636 & ~a34634;
assign a34640 = a34632 & a32970;
assign a34642 = ~a32970 & l1680;
assign a34644 = ~a34642 & ~a34640;
assign a34646 = a34632 & a32990;
assign a34648 = ~a32990 & l1682;
assign a34650 = ~a34648 & ~a34646;
assign a34652 = a34632 & a33006;
assign a34654 = ~a33006 & l1684;
assign a34656 = ~a34654 & ~a34652;
assign a34658 = a34632 & a33024;
assign a34660 = ~a33024 & l1686;
assign a34662 = ~a34660 & ~a34658;
assign a34664 = a34632 & a33038;
assign a34666 = ~a33038 & l1688;
assign a34668 = ~a34666 & ~a34664;
assign a34670 = a34632 & a33058;
assign a34672 = ~a33058 & l1690;
assign a34674 = ~a34672 & ~a34670;
assign a34676 = a34632 & a33070;
assign a34678 = ~a33070 & l1692;
assign a34680 = ~a34678 & ~a34676;
assign a34682 = a34632 & a33086;
assign a34684 = ~a33086 & ~a13452;
assign a34688 = a34632 & a33098;
assign a34690 = ~a33098 & ~a13466;
assign a34694 = a23672 & ~a13590;
assign a34696 = ~a23672 & i442;
assign a34698 = ~a34696 & ~a34694;
assign a34700 = a34698 & a32956;
assign a34702 = ~a32956 & l1698;
assign a34704 = ~a34702 & ~a34700;
assign a34706 = a34698 & a32970;
assign a34708 = ~a32970 & l1700;
assign a34710 = ~a34708 & ~a34706;
assign a34712 = a34698 & a32990;
assign a34714 = ~a32990 & l1702;
assign a34716 = ~a34714 & ~a34712;
assign a34718 = a34698 & a33006;
assign a34720 = ~a33006 & l1704;
assign a34722 = ~a34720 & ~a34718;
assign a34724 = a34698 & a33024;
assign a34726 = ~a33024 & l1706;
assign a34728 = ~a34726 & ~a34724;
assign a34730 = a34698 & a33038;
assign a34732 = ~a33038 & l1708;
assign a34734 = ~a34732 & ~a34730;
assign a34736 = a34698 & a33058;
assign a34738 = ~a33058 & l1710;
assign a34740 = ~a34738 & ~a34736;
assign a34742 = a34698 & a33070;
assign a34744 = ~a33070 & l1712;
assign a34746 = ~a34744 & ~a34742;
assign a34748 = a34698 & a33086;
assign a34750 = ~a33086 & ~a13642;
assign a34754 = a34698 & a33098;
assign a34756 = ~a33098 & ~a13656;
assign a34760 = a23672 & ~a13780;
assign a34762 = ~a23672 & i446;
assign a34764 = ~a34762 & ~a34760;
assign a34766 = a34764 & a32956;
assign a34768 = ~a32956 & l1718;
assign a34770 = ~a34768 & ~a34766;
assign a34772 = a34764 & a32970;
assign a34774 = ~a32970 & l1720;
assign a34776 = ~a34774 & ~a34772;
assign a34778 = a34764 & a32990;
assign a34780 = ~a32990 & l1722;
assign a34782 = ~a34780 & ~a34778;
assign a34784 = a34764 & a33006;
assign a34786 = ~a33006 & l1724;
assign a34788 = ~a34786 & ~a34784;
assign a34790 = a34764 & a33024;
assign a34792 = ~a33024 & l1726;
assign a34794 = ~a34792 & ~a34790;
assign a34796 = a34764 & a33038;
assign a34798 = ~a33038 & l1728;
assign a34800 = ~a34798 & ~a34796;
assign a34802 = a34764 & a33058;
assign a34804 = ~a33058 & l1730;
assign a34806 = ~a34804 & ~a34802;
assign a34808 = a34764 & a33070;
assign a34810 = ~a33070 & l1732;
assign a34812 = ~a34810 & ~a34808;
assign a34814 = a34764 & a33086;
assign a34816 = ~a33086 & ~a13832;
assign a34820 = a34764 & a33098;
assign a34822 = ~a33098 & l1736;
assign a34824 = ~a34822 & ~a34820;
assign a34826 = a23672 & a13958;
assign a34828 = ~a23672 & i450;
assign a34830 = ~a34828 & ~a34826;
assign a34832 = a34830 & a32956;
assign a34834 = ~a32956 & l1738;
assign a34836 = ~a34834 & ~a34832;
assign a34838 = a34830 & a32970;
assign a34840 = ~a32970 & l1740;
assign a34842 = ~a34840 & ~a34838;
assign a34844 = a34830 & a32990;
assign a34846 = ~a32990 & l1742;
assign a34848 = ~a34846 & ~a34844;
assign a34850 = a34830 & a33006;
assign a34852 = ~a33006 & l1744;
assign a34854 = ~a34852 & ~a34850;
assign a34856 = a34830 & a33024;
assign a34858 = ~a33024 & l1746;
assign a34860 = ~a34858 & ~a34856;
assign a34862 = a34830 & a33038;
assign a34864 = ~a33038 & l1748;
assign a34866 = ~a34864 & ~a34862;
assign a34868 = a34830 & a33058;
assign a34870 = ~a33058 & l1750;
assign a34872 = ~a34870 & ~a34868;
assign a34874 = a34830 & a33070;
assign a34876 = ~a33070 & l1752;
assign a34878 = ~a34876 & ~a34874;
assign a34880 = a34830 & a33086;
assign a34882 = ~a33086 & l1754;
assign a34884 = ~a34882 & ~a34880;
assign a34886 = a34830 & a33098;
assign a34888 = ~a33098 & l1756;
assign a34890 = ~a34888 & ~a34886;
assign a34892 = ~a14368 & a5408;
assign a34906 = ~a19884 & ~a18856;
assign a34908 = ~a31036 & a19884;
assign a34912 = a31024 & a2740;
assign a34914 = a34912 & ~l1156;
assign a34916 = ~a34914 & l1784;
assign a34918 = a34914 & ~a31036;
assign a34920 = ~a34918 & ~a34916;
assign a34922 = a19882 & ~a2740;
assign a34924 = ~a34922 & l1786;
assign a34926 = a34922 & ~a31036;
assign a34928 = ~a34926 & ~a34924;
assign a34930 = a34912 & l1156;
assign a34932 = ~a34930 & l1788;
assign a34934 = a34930 & ~a31036;
assign a34936 = ~a34934 & ~a34932;
assign a34938 = a19880 & l1156;
assign a34940 = a34938 & a2740;
assign a34942 = ~a34940 & l1790;
assign a34944 = a34940 & ~a31036;
assign a34946 = ~a34944 & ~a34942;
assign a34948 = a31026 & l1156;
assign a34950 = ~a34948 & l1792;
assign a34952 = a34948 & ~a31036;
assign a34954 = ~a34952 & ~a34950;
assign a34956 = a34938 & ~a2740;
assign a34958 = ~a34956 & l1794;
assign a34960 = a34956 & ~a31036;
assign a34962 = ~a34960 & ~a34958;
assign a34964 = a33510 & a31022;
assign a34966 = ~a34964 & l1796;
assign a34968 = a34964 & ~a31036;
assign a34970 = ~a34968 & ~a34966;
assign a34972 = ~a33512 & l1798;
assign a34974 = a33512 & ~a31036;
assign a34976 = ~a34974 & ~a34972;
assign a34978 = ~a19884 & ~a18930;
assign a34980 = ~l1802 & l890;
assign a34982 = ~a11330 & ~l890;
assign a34984 = ~a34982 & ~a34980;
assign a34986 = ~a34984 & a19884;
assign a34990 = ~a34914 & l1804;
assign a34992 = ~a34984 & a34914;
assign a34994 = ~a34992 & ~a34990;
assign a34996 = ~a31028 & ~a18946;
assign a34998 = ~a34984 & a31028;
assign a35002 = ~a34922 & l1808;
assign a35004 = ~a34984 & a34922;
assign a35006 = ~a35004 & ~a35002;
assign a35008 = ~a34930 & l1810;
assign a35010 = ~a34984 & a34930;
assign a35012 = ~a35010 & ~a35008;
assign a35014 = ~a34940 & l1812;
assign a35016 = ~a34984 & a34940;
assign a35018 = ~a35016 & ~a35014;
assign a35020 = ~a34948 & l1814;
assign a35022 = ~a34984 & a34948;
assign a35024 = ~a35022 & ~a35020;
assign a35026 = ~a34956 & l1816;
assign a35028 = ~a34984 & a34956;
assign a35030 = ~a35028 & ~a35026;
assign a35032 = ~a34964 & l1818;
assign a35034 = ~a34984 & a34964;
assign a35036 = ~a35034 & ~a35032;
assign a35038 = ~a33512 & l1820;
assign a35040 = ~a34984 & a33512;
assign a35042 = ~a35040 & ~a35038;
assign a35044 = ~a19884 & ~a19010;
assign a35046 = ~l1824 & l890;
assign a35048 = ~a11372 & ~l890;
assign a35050 = ~a35048 & ~a35046;
assign a35052 = ~a35050 & a19884;
assign a35056 = ~a34914 & l1826;
assign a35058 = ~a35050 & a34914;
assign a35060 = ~a35058 & ~a35056;
assign a35062 = ~a31028 & ~a19026;
assign a35064 = ~a35050 & a31028;
assign a35068 = ~a34922 & l1830;
assign a35070 = ~a35050 & a34922;
assign a35072 = ~a35070 & ~a35068;
assign a35074 = ~a34930 & l1832;
assign a35076 = ~a35050 & a34930;
assign a35078 = ~a35076 & ~a35074;
assign a35080 = ~a34940 & l1834;
assign a35082 = ~a35050 & a34940;
assign a35084 = ~a35082 & ~a35080;
assign a35086 = ~a34948 & l1836;
assign a35088 = ~a35050 & a34948;
assign a35090 = ~a35088 & ~a35086;
assign a35092 = ~a34956 & l1838;
assign a35094 = ~a35050 & a34956;
assign a35096 = ~a35094 & ~a35092;
assign a35098 = ~a34964 & l1840;
assign a35100 = ~a35050 & a34964;
assign a35102 = ~a35100 & ~a35098;
assign a35104 = ~a33512 & l1842;
assign a35106 = ~a35050 & a33512;
assign a35108 = ~a35106 & ~a35104;
assign a35110 = ~a19884 & ~a19092;
assign a35112 = ~l1846 & l890;
assign a35114 = ~a11414 & ~l890;
assign a35116 = ~a35114 & ~a35112;
assign a35118 = ~a35116 & a19884;
assign a35122 = ~a34914 & l1848;
assign a35124 = ~a35116 & a34914;
assign a35126 = ~a35124 & ~a35122;
assign a35128 = ~a31028 & ~a19108;
assign a35130 = ~a35116 & a31028;
assign a35134 = ~a34922 & l1852;
assign a35136 = ~a35116 & a34922;
assign a35138 = ~a35136 & ~a35134;
assign a35140 = ~a34930 & l1854;
assign a35142 = ~a35116 & a34930;
assign a35144 = ~a35142 & ~a35140;
assign a35146 = ~a34940 & l1856;
assign a35148 = ~a35116 & a34940;
assign a35150 = ~a35148 & ~a35146;
assign a35152 = ~a34948 & l1858;
assign a35154 = ~a35116 & a34948;
assign a35156 = ~a35154 & ~a35152;
assign a35158 = ~a34956 & l1860;
assign a35160 = ~a35116 & a34956;
assign a35162 = ~a35160 & ~a35158;
assign a35164 = ~a34964 & l1862;
assign a35166 = ~a35116 & a34964;
assign a35168 = ~a35166 & ~a35164;
assign a35170 = ~a33512 & l1864;
assign a35172 = ~a35116 & a33512;
assign a35174 = ~a35172 & ~a35170;
assign a35176 = ~a19884 & ~a19174;
assign a35178 = ~l1868 & l890;
assign a35180 = ~a11456 & ~l890;
assign a35182 = ~a35180 & ~a35178;
assign a35184 = ~a35182 & a19884;
assign a35188 = ~a34914 & l1870;
assign a35190 = ~a35182 & a34914;
assign a35192 = ~a35190 & ~a35188;
assign a35194 = ~a31028 & ~a19190;
assign a35196 = ~a35182 & a31028;
assign a35200 = ~a34922 & l1874;
assign a35202 = ~a35182 & a34922;
assign a35204 = ~a35202 & ~a35200;
assign a35206 = ~a34930 & l1876;
assign a35208 = ~a35182 & a34930;
assign a35210 = ~a35208 & ~a35206;
assign a35212 = ~a34940 & l1878;
assign a35214 = ~a35182 & a34940;
assign a35216 = ~a35214 & ~a35212;
assign a35218 = ~a34948 & l1880;
assign a35220 = ~a35182 & a34948;
assign a35222 = ~a35220 & ~a35218;
assign a35224 = ~a34956 & l1882;
assign a35226 = ~a35182 & a34956;
assign a35228 = ~a35226 & ~a35224;
assign a35230 = ~a34964 & l1884;
assign a35232 = ~a35182 & a34964;
assign a35234 = ~a35232 & ~a35230;
assign a35236 = ~a33512 & l1886;
assign a35238 = ~a35182 & a33512;
assign a35240 = ~a35238 & ~a35236;
assign a35242 = ~a19884 & ~a19256;
assign a35244 = ~l1890 & l890;
assign a35246 = ~a11498 & ~l890;
assign a35248 = ~a35246 & ~a35244;
assign a35250 = ~a35248 & a19884;
assign a35254 = ~a34914 & l1892;
assign a35256 = ~a35248 & a34914;
assign a35258 = ~a35256 & ~a35254;
assign a35260 = ~a31028 & ~a19272;
assign a35262 = ~a35248 & a31028;
assign a35266 = ~a34922 & l1896;
assign a35268 = ~a35248 & a34922;
assign a35270 = ~a35268 & ~a35266;
assign a35272 = ~a34930 & l1898;
assign a35274 = ~a35248 & a34930;
assign a35276 = ~a35274 & ~a35272;
assign a35278 = ~a34940 & l1900;
assign a35280 = ~a35248 & a34940;
assign a35282 = ~a35280 & ~a35278;
assign a35284 = ~a34948 & l1902;
assign a35286 = ~a35248 & a34948;
assign a35288 = ~a35286 & ~a35284;
assign a35290 = ~a34956 & l1904;
assign a35292 = ~a35248 & a34956;
assign a35294 = ~a35292 & ~a35290;
assign a35296 = ~a34964 & l1906;
assign a35298 = ~a35248 & a34964;
assign a35300 = ~a35298 & ~a35296;
assign a35302 = ~a33512 & l1908;
assign a35304 = ~a35248 & a33512;
assign a35306 = ~a35304 & ~a35302;
assign a35308 = ~a19884 & l1910;
assign a35310 = ~l1912 & l890;
assign a35312 = ~a11540 & ~l890;
assign a35314 = ~a35312 & ~a35310;
assign a35316 = ~a35314 & a19884;
assign a35318 = ~a35316 & ~a35308;
assign a35320 = ~a34914 & l1914;
assign a35322 = ~a35314 & a34914;
assign a35324 = ~a35322 & ~a35320;
assign a35326 = ~a31028 & ~a19348;
assign a35328 = ~a35314 & a31028;
assign a35332 = ~a34922 & l1918;
assign a35334 = ~a35314 & a34922;
assign a35336 = ~a35334 & ~a35332;
assign a35338 = ~a34930 & l1920;
assign a35340 = ~a35314 & a34930;
assign a35342 = ~a35340 & ~a35338;
assign a35344 = ~a34940 & l1922;
assign a35346 = ~a35314 & a34940;
assign a35348 = ~a35346 & ~a35344;
assign a35350 = ~a34948 & l1924;
assign a35352 = ~a35314 & a34948;
assign a35354 = ~a35352 & ~a35350;
assign a35356 = ~a34956 & l1926;
assign a35358 = ~a35314 & a34956;
assign a35360 = ~a35358 & ~a35356;
assign a35362 = ~a34964 & l1928;
assign a35364 = ~a35314 & a34964;
assign a35366 = ~a35364 & ~a35362;
assign a35368 = ~a33512 & l1930;
assign a35370 = ~a35314 & a33512;
assign a35372 = ~a35370 & ~a35368;
assign a35374 = ~a19884 & l1932;
assign a35376 = ~l1934 & l890;
assign a35378 = i486 & ~i92;
assign a35380 = a35378 & ~l890;
assign a35382 = ~a35380 & ~a35376;
assign a35384 = ~a35382 & a19884;
assign a35386 = ~a35384 & ~a35374;
assign a35388 = ~a34914 & l1936;
assign a35390 = ~a35382 & a34914;
assign a35392 = ~a35390 & ~a35388;
assign a35394 = ~a31028 & l1938;
assign a35396 = ~a35382 & a31028;
assign a35398 = ~a35396 & ~a35394;
assign a35400 = ~a34922 & l1940;
assign a35402 = ~a35382 & a34922;
assign a35404 = ~a35402 & ~a35400;
assign a35406 = ~a34930 & l1942;
assign a35408 = ~a35382 & a34930;
assign a35410 = ~a35408 & ~a35406;
assign a35412 = ~a34940 & l1944;
assign a35414 = ~a35382 & a34940;
assign a35416 = ~a35414 & ~a35412;
assign a35418 = ~a34948 & l1946;
assign a35420 = ~a35382 & a34948;
assign a35422 = ~a35420 & ~a35418;
assign a35424 = ~a34956 & l1948;
assign a35426 = ~a35382 & a34956;
assign a35428 = ~a35426 & ~a35424;
assign a35430 = ~a34964 & l1950;
assign a35432 = ~a35382 & a34964;
assign a35434 = ~a35432 & ~a35430;
assign a35436 = ~a33512 & l1952;
assign a35438 = ~a35382 & a33512;
assign a35440 = ~a35438 & ~a35436;
assign a35442 = a2740 & ~l1964;
assign a35444 = a35442 & a19758;
assign a35446 = a35444 & ~l1156;
assign a35448 = a35446 & ~l1244;
assign a35450 = ~a35448 & ~a19838;
assign a35452 = ~a19830 & a19802;
assign a35454 = a35452 & a35450;
assign a35456 = ~a19816 & ~a19762;
assign a35458 = a35456 & a35454;
assign a35460 = ~a35458 & l924;
assign a35462 = l1150 & ~l1148;
assign a35464 = a35462 & a6538;
assign a35466 = ~a34914 & ~a18582;
assign a35468 = ~a35466 & ~l886;
assign a35470 = a35468 & ~a35464;
assign a35474 = ~l1968 & ~l1956;
assign a35476 = a35474 & l1156;
assign a35478 = a19774 & a19766;
assign a35480 = a35478 & a2740;
assign a35482 = ~a35480 & ~a35476;
assign a35484 = a35474 & ~l1964;
assign a35486 = ~a2768 & l1244;
assign a35488 = a35486 & a35484;
assign a35490 = ~a2740 & ~l1956;
assign a35492 = a35490 & ~l1156;
assign a35494 = ~a35492 & ~a35488;
assign a35496 = a35494 & a35482;
assign a35498 = a35496 & a19810;
assign a35500 = ~a35498 & l924;
assign a35502 = l1162 & l1150;
assign a35504 = a35502 & ~l1166;
assign a35506 = a35504 & ~l1148;
assign a35508 = ~a31028 & ~a18596;
assign a35510 = ~a35508 & ~l886;
assign a35512 = a35510 & ~a35506;
assign a35516 = a19836 & a19764;
assign a35518 = ~a35516 & ~a35488;
assign a35520 = a35518 & a19772;
assign a35522 = a35492 & ~a2768;
assign a35524 = ~a2768 & ~l1960;
assign a35526 = a35524 & ~a2740;
assign a35528 = a35526 & ~l1156;
assign a35530 = a19806 & ~a2768;
assign a35532 = ~a35530 & ~a19826;
assign a35534 = a35532 & ~a35528;
assign a35536 = a35534 & ~a35522;
assign a35538 = a35536 & a35482;
assign a35540 = a35538 & a19800;
assign a35542 = a35540 & a35520;
assign a35544 = ~a35542 & l924;
assign a35546 = a30096 & l1150;
assign a35548 = ~a34922 & ~l1974;
assign a35550 = ~a35548 & ~l886;
assign a35552 = a35550 & ~a35546;
assign a35556 = a35442 & a19776;
assign a35558 = ~a35556 & ~a19780;
assign a35560 = a35558 & a35520;
assign a35562 = a35560 & ~a19788;
assign a35564 = a35562 & a19798;
assign a35566 = ~l1968 & l1956;
assign a35568 = a33508 & ~a2768;
assign a35570 = a35568 & a35566;
assign a35572 = ~l1968 & l1156;
assign a35574 = ~a35572 & ~a35570;
assign a35576 = a35574 & a35564;
assign a35578 = ~a35576 & l924;
assign a35580 = a35462 & a30102;
assign a35582 = ~a34930 & ~l1976;
assign a35584 = ~a35582 & ~l886;
assign a35586 = a35584 & ~a35580;
assign a35590 = a35572 & ~a2740;
assign a35592 = ~a35590 & ~a35570;
assign a35594 = a35592 & ~a19796;
assign a35596 = a35594 & a35560;
assign a35598 = a35572 & ~a2768;
assign a35600 = l1968 & ~l1960;
assign a35602 = a35600 & ~l1156;
assign a35604 = a35602 & ~l1956;
assign a35606 = ~a2740 & l1156;
assign a35608 = a35606 & a19820;
assign a35610 = a35524 & a19792;
assign a35612 = ~a2768 & l1156;
assign a35614 = a35612 & a19834;
assign a35616 = ~a35614 & ~a35610;
assign a35618 = a35616 & ~a35608;
assign a35620 = a35618 & ~a35604;
assign a35622 = a35620 & ~a35598;
assign a35624 = a35622 & a35596;
assign a35626 = ~a35624 & l924;
assign a35628 = a30102 & a19866;
assign a35630 = ~a34940 & ~l1978;
assign a35632 = ~a35630 & ~l886;
assign a35634 = a35632 & ~a35628;
assign a35638 = l1968 & ~l1956;
assign a35640 = a35638 & ~l1156;
assign a35642 = a35490 & l1156;
assign a35644 = ~a35642 & ~a35640;
assign a35646 = a35644 & ~a19788;
assign a35648 = a35646 & a35596;
assign a35650 = ~a35648 & l924;
assign a35652 = a35502 & l1166;
assign a35654 = a35652 & ~l1164;
assign a35656 = a35654 & ~l1148;
assign a35658 = ~a34948 & ~l1980;
assign a35660 = ~a35658 & ~l886;
assign a35662 = a35660 & ~a35656;
assign a35666 = a35642 & ~a2768;
assign a35668 = a35590 & ~a2768;
assign a35670 = ~a2768 & ~a2740;
assign a35672 = a35670 & a35600;
assign a35674 = a35600 & a19834;
assign a35676 = ~a35640 & ~a35602;
assign a35678 = a35676 & ~a35570;
assign a35680 = a35678 & ~a35674;
assign a35682 = a35680 & ~a35672;
assign a35684 = a35682 & ~a35668;
assign a35686 = a35684 & ~a35666;
assign a35688 = a35686 & a35562;
assign a35690 = ~a35688 & l924;
assign a35692 = a35654 & l1148;
assign a35694 = ~a34956 & ~l1982;
assign a35696 = ~a35694 & ~l886;
assign a35698 = a35696 & ~a35692;
assign a35702 = l1956 & l1244;
assign a35704 = ~a35640 & ~a19840;
assign a35706 = a35704 & ~a19830;
assign a35708 = a35706 & ~a35702;
assign a35710 = a35708 & a35564;
assign a35712 = ~a35710 & l924;
assign a35714 = a30132 & l1150;
assign a35716 = ~a34964 & ~a18646;
assign a35718 = ~a35716 & ~a35714;
assign a35722 = a19804 & ~a2768;
assign a35724 = a35524 & l1244;
assign a35726 = a19816 & ~l1960;
assign a35728 = ~a35570 & ~a35488;
assign a35730 = a35728 & ~a35726;
assign a35732 = a35730 & ~a35724;
assign a35734 = a35732 & ~a35722;
assign a35736 = a35734 & a35454;
assign a35738 = ~a35736 & l924;
assign a35740 = a19868 & l1164;
assign a35742 = ~a33512 & ~l1986;
assign a35744 = ~a35742 & ~l886;
assign a35746 = a35744 & ~a35740;
assign a35750 = ~a34964 & l1988;
assign a35752 = a34964 & a33522;
assign a35754 = ~a35752 & ~a35750;
assign a35756 = ~a34956 & l1990;
assign a35758 = a34956 & a33522;
assign a35760 = ~a35758 & ~a35756;
assign a35762 = ~a34948 & l1992;
assign a35764 = a34948 & a33522;
assign a35766 = ~a35764 & ~a35762;
assign a35768 = ~a34940 & l1994;
assign a35770 = a34940 & a33522;
assign a35772 = ~a35770 & ~a35768;
assign a35774 = ~a34930 & l1996;
assign a35776 = a34930 & a33522;
assign a35778 = ~a35776 & ~a35774;
assign a35780 = ~a34922 & l1998;
assign a35782 = a34922 & a33522;
assign a35784 = ~a35782 & ~a35780;
assign a35786 = ~a31028 & l2000;
assign a35788 = a33522 & a31028;
assign a35790 = ~a35788 & ~a35786;
assign a35792 = ~a19884 & l2002;
assign a35794 = a33522 & a19884;
assign a35796 = ~a35794 & ~a35792;
assign a35798 = ~a34914 & l2004;
assign a35800 = a34914 & a33522;
assign a35802 = ~a35800 & ~a35798;
assign a35804 = ~l908 & l892;
assign a35806 = l2036 & l2032;
assign a35808 = a35806 & l2028;
assign a35810 = l2040 & ~l2036;
assign a35812 = ~a35810 & ~a35808;
assign a35814 = ~a35812 & a35804;
assign a35816 = l2044 & l908;
assign a35818 = ~l908 & ~l886;
assign a35820 = a35818 & ~a18526;
assign a35822 = a35820 & ~l892;
assign a35824 = a35822 & l2040;
assign a35826 = ~a35824 & ~a35816;
assign a35828 = a35826 & ~a35814;
assign a35830 = a25830 & a16216;
assign a35832 = a35830 & l2040;
assign a35834 = ~a35830 & l2044;
assign a35836 = ~a35834 & ~a35832;
assign a35838 = ~l2032 & l2028;
assign a35840 = ~l2036 & l2028;
assign a35842 = a35806 & ~l2028;
assign a35844 = ~a35842 & ~a35840;
assign a35846 = a35844 & ~a35838;
assign a35848 = ~a35846 & a35804;
assign a35850 = l2048 & l908;
assign a35852 = a35822 & l2028;
assign a35854 = ~a35852 & ~a35850;
assign a35856 = a35854 & ~a35848;
assign a35858 = a35830 & l2028;
assign a35860 = ~a35830 & l2048;
assign a35862 = ~a35860 & ~a35858;
assign a35864 = ~l2040 & l2036;
assign a35866 = a35864 & ~l2032;
assign a35868 = ~l2036 & l2032;
assign a35870 = ~a35868 & ~a35866;
assign a35872 = ~a35870 & a35804;
assign a35874 = l2052 & l908;
assign a35876 = a35822 & l2032;
assign a35878 = ~a35876 & ~a35874;
assign a35880 = a35878 & ~a35872;
assign a35882 = a35830 & l2032;
assign a35884 = ~a35830 & l2052;
assign a35886 = ~a35884 & ~a35882;
assign a35888 = a35804 & ~l2036;
assign a35890 = l2056 & l908;
assign a35892 = a35822 & l2036;
assign a35894 = ~a35892 & ~a35890;
assign a35896 = a35894 & ~a35888;
assign a35898 = a35830 & l2036;
assign a35900 = ~a35830 & l2056;
assign a35902 = ~a35900 & ~a35898;
assign a35904 = a25350 & ~a22550;
assign a35906 = ~a25350 & l2058;
assign a35908 = ~a35906 & ~a35904;
assign a35910 = ~a35908 & ~a17272;
assign a35912 = ~a35910 & ~a17602;
assign a35914 = a25350 & ~a22808;
assign a35916 = ~a25350 & l2060;
assign a35918 = ~a35916 & ~a35914;
assign a35920 = ~a35918 & ~a17272;
assign a35922 = ~a35920 & ~a17438;
assign a35924 = a21692 & a16198;
assign a35926 = ~a35924 & ~a18532;
assign a35928 = ~a35926 & ~l886;
assign a35932 = ~l2070 & l890;
assign a35934 = ~a5346 & i546;
assign a35936 = a35934 & ~a5178;
assign a35938 = ~a35936 & ~l890;
assign a35940 = ~a35938 & ~a35932;
assign a35942 = a35940 & ~a17658;
assign a35944 = a35942 & ~a19756;
assign a35948 = ~l2072 & l890;
assign a35950 = ~a5346 & ~a5178;
assign a35952 = a35950 & i548;
assign a35954 = ~a35952 & ~l890;
assign a35956 = ~a35954 & ~a35948;
assign a35958 = a35956 & ~a17658;
assign a35962 = ~a17658 & ~a14378;
assign a35964 = a35962 & i550;
assign a35966 = a35964 & ~a5352;
assign a35970 = l2076 & ~l2074;
assign a35972 = ~l2084 & l2078;
assign a35974 = ~a35972 & ~a35970;
assign a35976 = l2084 & ~l2078;
assign a35978 = ~a35976 & ~a35974;
assign a35980 = ~l2086 & l2082;
assign a35982 = ~a35980 & ~a35978;
assign a35984 = l2086 & ~l2082;
assign a35986 = ~a35984 & ~a35982;
assign a35988 = ~l2088 & l2080;
assign a35990 = ~a35988 & ~a35986;
assign a35992 = l2088 & ~l2080;
assign a35994 = ~a35992 & ~a35990;
assign a35996 = ~l2092 & l2090;
assign a35998 = l2092 & ~l2090;
assign a36000 = ~a35998 & ~a35996;
assign a36002 = a36000 & a35994;
assign a36004 = ~l2076 & l2074;
assign a36006 = ~a36004 & ~a35976;
assign a36008 = ~a36006 & ~a35972;
assign a36010 = ~a36008 & ~a35984;
assign a36012 = ~a36010 & ~a35980;
assign a36014 = ~a36012 & ~a35992;
assign a36016 = ~a36014 & ~a35988;
assign a36018 = a36016 & ~a36000;
assign a36020 = ~a36018 & ~a36002;
assign a36022 = ~l2084 & l2074;
assign a36024 = a36022 & l2088;
assign a36026 = ~a36024 & ~a36020;
assign a36028 = a36026 & ~l2074;
assign a36030 = ~a36000 & a35994;
assign a36032 = a36016 & a36000;
assign a36034 = ~a36032 & ~a36030;
assign a36036 = ~l2084 & ~l2074;
assign a36038 = a36036 & ~l2086;
assign a36040 = a36038 & ~l2088;
assign a36042 = ~a36040 & ~a36034;
assign a36044 = a36042 & ~l2074;
assign a36046 = a36040 & ~a36034;
assign a36048 = ~a36046 & ~l2074;
assign a36050 = ~a36048 & ~a36042;
assign a36052 = ~a36050 & ~a36044;
assign a36054 = ~a36052 & a36020;
assign a36056 = ~a36054 & ~a36028;
assign a36058 = ~l1332 & l978;
assign a36060 = l1332 & ~l978;
assign a36062 = ~a36060 & ~a36058;
assign a36064 = a6254 & l1352;
assign a36066 = a6262 & l1372;
assign a36068 = ~a36066 & ~a36064;
assign a36070 = ~a6262 & ~l1372;
assign a36072 = ~a36070 & ~a36068;
assign a36074 = a6270 & l1392;
assign a36076 = ~a36074 & ~a36072;
assign a36078 = ~a6270 & ~l1392;
assign a36080 = ~a36078 & ~a36076;
assign a36082 = a6278 & l1412;
assign a36084 = ~a36082 & ~a36080;
assign a36086 = ~a6278 & ~l1412;
assign a36088 = ~a36086 & ~a36084;
assign a36090 = a6286 & l1432;
assign a36092 = ~a36090 & ~a36088;
assign a36094 = ~a6286 & ~l1432;
assign a36096 = ~a36094 & ~a36092;
assign a36098 = l1452 & ~l1054;
assign a36100 = ~a36098 & ~a36096;
assign a36102 = ~l1452 & l1054;
assign a36104 = ~a36102 & ~a36100;
assign a36106 = l1472 & ~l1058;
assign a36108 = ~a36106 & ~a36104;
assign a36110 = ~l1472 & l1058;
assign a36112 = ~a36110 & ~a36108;
assign a36114 = ~a36112 & a36062;
assign a36116 = ~a6254 & ~l1352;
assign a36118 = ~a36116 & ~a36070;
assign a36120 = ~a36118 & ~a36066;
assign a36122 = ~a36120 & ~a36078;
assign a36124 = ~a36122 & ~a36074;
assign a36126 = ~a36124 & ~a36086;
assign a36128 = ~a36126 & ~a36082;
assign a36130 = ~a36128 & ~a36094;
assign a36132 = ~a36130 & ~a36090;
assign a36134 = ~a36132 & ~a36102;
assign a36136 = ~a36134 & ~a36098;
assign a36138 = ~a36136 & ~a36110;
assign a36140 = ~a36138 & ~a36106;
assign a36142 = ~a36140 & ~a36062;
assign a36144 = ~a36142 & ~a36114;
assign a36146 = a36144 & a5568;
assign a36148 = ~a36146 & ~a15902;
assign a36150 = ~l1314 & l978;
assign a36152 = l1314 & ~l978;
assign a36154 = ~a36152 & ~a36150;
assign a36156 = a6254 & l1334;
assign a36158 = a6262 & l1354;
assign a36160 = ~a36158 & ~a36156;
assign a36162 = ~a6262 & ~l1354;
assign a36164 = ~a36162 & ~a36160;
assign a36166 = a6270 & l1374;
assign a36168 = ~a36166 & ~a36164;
assign a36170 = ~a6270 & ~l1374;
assign a36172 = ~a36170 & ~a36168;
assign a36174 = a6278 & l1394;
assign a36176 = ~a36174 & ~a36172;
assign a36178 = ~a6278 & ~l1394;
assign a36180 = ~a36178 & ~a36176;
assign a36182 = a6286 & l1414;
assign a36184 = ~a36182 & ~a36180;
assign a36186 = ~a6286 & ~l1414;
assign a36188 = ~a36186 & ~a36184;
assign a36190 = l1434 & ~l1054;
assign a36192 = ~a36190 & ~a36188;
assign a36194 = ~l1434 & l1054;
assign a36196 = ~a36194 & ~a36192;
assign a36198 = l1454 & ~l1058;
assign a36200 = ~a36198 & ~a36196;
assign a36202 = ~l1454 & l1058;
assign a36204 = ~a36202 & ~a36200;
assign a36206 = ~a36204 & a36154;
assign a36208 = ~a6254 & ~l1334;
assign a36210 = ~a36208 & ~a36162;
assign a36212 = ~a36210 & ~a36158;
assign a36214 = ~a36212 & ~a36170;
assign a36216 = ~a36214 & ~a36166;
assign a36218 = ~a36216 & ~a36178;
assign a36220 = ~a36218 & ~a36174;
assign a36222 = ~a36220 & ~a36186;
assign a36224 = ~a36222 & ~a36182;
assign a36226 = ~a36224 & ~a36194;
assign a36228 = ~a36226 & ~a36190;
assign a36230 = ~a36228 & ~a36202;
assign a36232 = ~a36230 & ~a36198;
assign a36234 = ~a36232 & ~a36154;
assign a36236 = ~a36234 & ~a36206;
assign a36238 = ~a36236 & ~a36148;
assign a36240 = a36238 & l968;
assign a36242 = ~a36240 & ~l886;
assign a36244 = ~l2078 & l2076;
assign a36246 = ~l2082 & l2080;
assign a36248 = a36246 & a36244;
assign a36250 = a36248 & ~a36242;
assign a36252 = a36250 & l886;
assign a36254 = ~l1322 & l978;
assign a36256 = l1322 & ~l978;
assign a36258 = ~a36256 & ~a36254;
assign a36260 = a6254 & l1342;
assign a36262 = a6262 & l1362;
assign a36264 = ~a36262 & ~a36260;
assign a36266 = ~a6262 & ~l1362;
assign a36268 = ~a36266 & ~a36264;
assign a36270 = a6270 & l1382;
assign a36272 = ~a36270 & ~a36268;
assign a36274 = ~a6270 & ~l1382;
assign a36276 = ~a36274 & ~a36272;
assign a36278 = a6278 & l1402;
assign a36280 = ~a36278 & ~a36276;
assign a36282 = ~a6278 & ~l1402;
assign a36284 = ~a36282 & ~a36280;
assign a36286 = a6286 & l1422;
assign a36288 = ~a36286 & ~a36284;
assign a36290 = ~a6286 & ~l1422;
assign a36292 = ~a36290 & ~a36288;
assign a36294 = l1442 & ~l1054;
assign a36296 = ~a36294 & ~a36292;
assign a36298 = ~l1442 & l1054;
assign a36300 = ~a36298 & ~a36296;
assign a36302 = l1462 & ~l1058;
assign a36304 = ~a36302 & ~a36300;
assign a36306 = ~l1462 & l1058;
assign a36308 = ~a36306 & ~a36304;
assign a36310 = ~a36308 & a36258;
assign a36312 = ~a6254 & ~l1342;
assign a36314 = ~a36312 & ~a36266;
assign a36316 = ~a36314 & ~a36262;
assign a36318 = ~a36316 & ~a36274;
assign a36320 = ~a36318 & ~a36270;
assign a36322 = ~a36320 & ~a36282;
assign a36324 = ~a36322 & ~a36278;
assign a36326 = ~a36324 & ~a36290;
assign a36328 = ~a36326 & ~a36286;
assign a36330 = ~a36328 & ~a36298;
assign a36332 = ~a36330 & ~a36294;
assign a36334 = ~a36332 & ~a36306;
assign a36336 = ~a36334 & ~a36302;
assign a36338 = ~a36336 & ~a36258;
assign a36340 = ~a36338 & ~a36310;
assign a36342 = ~l1320 & l978;
assign a36344 = l1320 & ~l978;
assign a36346 = ~a36344 & ~a36342;
assign a36348 = a6254 & l1340;
assign a36350 = a6262 & l1360;
assign a36352 = ~a36350 & ~a36348;
assign a36354 = ~a6262 & ~l1360;
assign a36356 = ~a36354 & ~a36352;
assign a36358 = a6270 & l1380;
assign a36360 = ~a36358 & ~a36356;
assign a36362 = ~a6270 & ~l1380;
assign a36364 = ~a36362 & ~a36360;
assign a36366 = a6278 & l1400;
assign a36368 = ~a36366 & ~a36364;
assign a36370 = ~a6278 & ~l1400;
assign a36372 = ~a36370 & ~a36368;
assign a36374 = a6286 & l1420;
assign a36376 = ~a36374 & ~a36372;
assign a36378 = ~a6286 & ~l1420;
assign a36380 = ~a36378 & ~a36376;
assign a36382 = l1440 & ~l1054;
assign a36384 = ~a36382 & ~a36380;
assign a36386 = ~l1440 & l1054;
assign a36388 = ~a36386 & ~a36384;
assign a36390 = l1460 & ~l1058;
assign a36392 = ~a36390 & ~a36388;
assign a36394 = ~l1460 & l1058;
assign a36396 = ~a36394 & ~a36392;
assign a36398 = ~a36396 & a36346;
assign a36400 = ~a6254 & ~l1340;
assign a36402 = ~a36400 & ~a36354;
assign a36404 = ~a36402 & ~a36350;
assign a36406 = ~a36404 & ~a36362;
assign a36408 = ~a36406 & ~a36358;
assign a36410 = ~a36408 & ~a36370;
assign a36412 = ~a36410 & ~a36366;
assign a36414 = ~a36412 & ~a36378;
assign a36416 = ~a36414 & ~a36374;
assign a36418 = ~a36416 & ~a36386;
assign a36420 = ~a36418 & ~a36382;
assign a36422 = ~a36420 & ~a36394;
assign a36424 = ~a36422 & ~a36390;
assign a36426 = ~a36424 & ~a36346;
assign a36428 = ~a36426 & ~a36398;
assign a36430 = a36428 & l964;
assign a36432 = ~a36430 & ~a15232;
assign a36434 = ~a36432 & ~a36340;
assign a36436 = a36434 & l962;
assign a36438 = ~a36436 & ~l886;
assign a36440 = ~a36438 & ~a36252;
assign a36442 = ~l1318 & l978;
assign a36444 = l1318 & ~l978;
assign a36446 = ~a36444 & ~a36442;
assign a36448 = a6254 & l1338;
assign a36450 = a6262 & l1358;
assign a36452 = ~a36450 & ~a36448;
assign a36454 = ~a6262 & ~l1358;
assign a36456 = ~a36454 & ~a36452;
assign a36458 = a6270 & l1378;
assign a36460 = ~a36458 & ~a36456;
assign a36462 = ~a6270 & ~l1378;
assign a36464 = ~a36462 & ~a36460;
assign a36466 = a6278 & l1398;
assign a36468 = ~a36466 & ~a36464;
assign a36470 = ~a6278 & ~l1398;
assign a36472 = ~a36470 & ~a36468;
assign a36474 = a6286 & l1418;
assign a36476 = ~a36474 & ~a36472;
assign a36478 = ~a6286 & ~l1418;
assign a36480 = ~a36478 & ~a36476;
assign a36482 = l1438 & ~l1054;
assign a36484 = ~a36482 & ~a36480;
assign a36486 = ~l1438 & l1054;
assign a36488 = ~a36486 & ~a36484;
assign a36490 = l1458 & ~l1058;
assign a36492 = ~a36490 & ~a36488;
assign a36494 = ~l1458 & l1058;
assign a36496 = ~a36494 & ~a36492;
assign a36498 = ~a36496 & a36446;
assign a36500 = ~a6254 & ~l1338;
assign a36502 = ~a36500 & ~a36454;
assign a36504 = ~a36502 & ~a36450;
assign a36506 = ~a36504 & ~a36462;
assign a36508 = ~a36506 & ~a36458;
assign a36510 = ~a36508 & ~a36470;
assign a36512 = ~a36510 & ~a36466;
assign a36514 = ~a36512 & ~a36478;
assign a36516 = ~a36514 & ~a36474;
assign a36518 = ~a36516 & ~a36486;
assign a36520 = ~a36518 & ~a36482;
assign a36522 = ~a36520 & ~a36494;
assign a36524 = ~a36522 & ~a36490;
assign a36526 = ~a36524 & ~a36446;
assign a36528 = ~a36526 & ~a36498;
assign a36530 = ~l1316 & l978;
assign a36532 = l1316 & ~l978;
assign a36534 = ~a36532 & ~a36530;
assign a36536 = a6254 & l1336;
assign a36538 = a6262 & l1356;
assign a36540 = ~a36538 & ~a36536;
assign a36542 = ~a6262 & ~l1356;
assign a36544 = ~a36542 & ~a36540;
assign a36546 = a6270 & l1376;
assign a36548 = ~a36546 & ~a36544;
assign a36550 = ~a6270 & ~l1376;
assign a36552 = ~a36550 & ~a36548;
assign a36554 = a6278 & l1396;
assign a36556 = ~a36554 & ~a36552;
assign a36558 = ~a6278 & ~l1396;
assign a36560 = ~a36558 & ~a36556;
assign a36562 = a6286 & l1416;
assign a36564 = ~a36562 & ~a36560;
assign a36566 = ~a6286 & ~l1416;
assign a36568 = ~a36566 & ~a36564;
assign a36570 = l1436 & ~l1054;
assign a36572 = ~a36570 & ~a36568;
assign a36574 = ~l1436 & l1054;
assign a36576 = ~a36574 & ~a36572;
assign a36578 = l1456 & ~l1058;
assign a36580 = ~a36578 & ~a36576;
assign a36582 = ~l1456 & l1058;
assign a36584 = ~a36582 & ~a36580;
assign a36586 = ~a36584 & a36534;
assign a36588 = ~a6254 & ~l1336;
assign a36590 = ~a36588 & ~a36542;
assign a36592 = ~a36590 & ~a36538;
assign a36594 = ~a36592 & ~a36550;
assign a36596 = ~a36594 & ~a36546;
assign a36598 = ~a36596 & ~a36558;
assign a36600 = ~a36598 & ~a36554;
assign a36602 = ~a36600 & ~a36566;
assign a36604 = ~a36602 & ~a36562;
assign a36606 = ~a36604 & ~a36574;
assign a36608 = ~a36606 & ~a36570;
assign a36610 = ~a36608 & ~a36582;
assign a36612 = ~a36610 & ~a36578;
assign a36614 = ~a36612 & ~a36534;
assign a36616 = ~a36614 & ~a36586;
assign a36618 = a36616 & l970;
assign a36620 = ~a36618 & ~a15564;
assign a36622 = ~a36620 & ~a36528;
assign a36624 = a36622 & l966;
assign a36626 = ~a36624 & ~l886;
assign a36628 = ~a36626 & ~a36252;
assign a36630 = ~l1326 & l978;
assign a36632 = l1326 & ~l978;
assign a36634 = ~a36632 & ~a36630;
assign a36636 = ~a12954 & a6254;
assign a36638 = ~a13138 & a6262;
assign a36640 = ~a36638 & ~a36636;
assign a36642 = a13138 & ~a6262;
assign a36644 = ~a36642 & ~a36640;
assign a36646 = ~a13328 & a6270;
assign a36648 = ~a36646 & ~a36644;
assign a36650 = a13328 & ~a6270;
assign a36652 = ~a36650 & ~a36648;
assign a36654 = ~a13518 & a6278;
assign a36656 = ~a36654 & ~a36652;
assign a36658 = a13518 & ~a6278;
assign a36660 = ~a36658 & ~a36656;
assign a36662 = ~a13708 & a6286;
assign a36664 = ~a36662 & ~a36660;
assign a36666 = a13708 & ~a6286;
assign a36668 = ~a36666 & ~a36664;
assign a36670 = ~a13886 & ~l1054;
assign a36672 = ~a36670 & ~a36668;
assign a36674 = a13886 & l1054;
assign a36676 = ~a36674 & ~a36672;
assign a36678 = ~a14050 & ~l1058;
assign a36680 = ~a36678 & ~a36676;
assign a36682 = a14050 & l1058;
assign a36684 = ~a36682 & ~a36680;
assign a36686 = ~a36684 & a36634;
assign a36688 = a12954 & ~a6254;
assign a36690 = ~a36688 & ~a36642;
assign a36692 = ~a36690 & ~a36638;
assign a36694 = ~a36692 & ~a36650;
assign a36696 = ~a36694 & ~a36646;
assign a36698 = ~a36696 & ~a36658;
assign a36700 = ~a36698 & ~a36654;
assign a36702 = ~a36700 & ~a36666;
assign a36704 = ~a36702 & ~a36662;
assign a36706 = ~a36704 & ~a36674;
assign a36708 = ~a36706 & ~a36670;
assign a36710 = ~a36708 & ~a36682;
assign a36712 = ~a36710 & ~a36678;
assign a36714 = ~a36712 & ~a36634;
assign a36716 = ~a36714 & ~a36686;
assign a36718 = ~l1324 & l978;
assign a36720 = l1324 & ~l978;
assign a36722 = ~a36720 & ~a36718;
assign a36724 = a6254 & l1344;
assign a36726 = a6262 & l1364;
assign a36728 = ~a36726 & ~a36724;
assign a36730 = ~a6262 & ~l1364;
assign a36732 = ~a36730 & ~a36728;
assign a36734 = a6270 & l1384;
assign a36736 = ~a36734 & ~a36732;
assign a36738 = ~a6270 & ~l1384;
assign a36740 = ~a36738 & ~a36736;
assign a36742 = a6278 & l1404;
assign a36744 = ~a36742 & ~a36740;
assign a36746 = ~a6278 & ~l1404;
assign a36748 = ~a36746 & ~a36744;
assign a36750 = a6286 & l1424;
assign a36752 = ~a36750 & ~a36748;
assign a36754 = ~a6286 & ~l1424;
assign a36756 = ~a36754 & ~a36752;
assign a36758 = l1444 & ~l1054;
assign a36760 = ~a36758 & ~a36756;
assign a36762 = ~l1444 & l1054;
assign a36764 = ~a36762 & ~a36760;
assign a36766 = l1464 & ~l1058;
assign a36768 = ~a36766 & ~a36764;
assign a36770 = ~l1464 & l1058;
assign a36772 = ~a36770 & ~a36768;
assign a36774 = ~a36772 & a36722;
assign a36776 = ~a6254 & ~l1344;
assign a36778 = ~a36776 & ~a36730;
assign a36780 = ~a36778 & ~a36726;
assign a36782 = ~a36780 & ~a36738;
assign a36784 = ~a36782 & ~a36734;
assign a36786 = ~a36784 & ~a36746;
assign a36788 = ~a36786 & ~a36742;
assign a36790 = ~a36788 & ~a36754;
assign a36792 = ~a36790 & ~a36750;
assign a36794 = ~a36792 & ~a36762;
assign a36796 = ~a36794 & ~a36758;
assign a36798 = ~a36796 & ~a36770;
assign a36800 = ~a36798 & ~a36766;
assign a36802 = ~a36800 & ~a36722;
assign a36804 = ~a36802 & ~a36774;
assign a36806 = a36804 & l960;
assign a36808 = ~a36806 & ~a14896;
assign a36810 = ~a36808 & ~a36716;
assign a36812 = a36810 & a5606;
assign a36814 = ~a36812 & ~l886;
assign a36816 = ~a36814 & ~a36252;
assign a36818 = ~l1330 & l978;
assign a36820 = l1330 & ~l978;
assign a36822 = ~a36820 & ~a36818;
assign a36824 = ~a12974 & a6254;
assign a36826 = ~a13158 & a6262;
assign a36828 = ~a36826 & ~a36824;
assign a36830 = a13158 & ~a6262;
assign a36832 = ~a36830 & ~a36828;
assign a36834 = ~a13348 & a6270;
assign a36836 = ~a36834 & ~a36832;
assign a36838 = a13348 & ~a6270;
assign a36840 = ~a36838 & ~a36836;
assign a36842 = ~a13538 & a6278;
assign a36844 = ~a36842 & ~a36840;
assign a36846 = a13538 & ~a6278;
assign a36848 = ~a36846 & ~a36844;
assign a36850 = ~a13728 & a6286;
assign a36852 = ~a36850 & ~a36848;
assign a36854 = a13728 & ~a6286;
assign a36856 = ~a36854 & ~a36852;
assign a36858 = ~a13906 & ~l1054;
assign a36860 = ~a36858 & ~a36856;
assign a36862 = a13906 & l1054;
assign a36864 = ~a36862 & ~a36860;
assign a36866 = l1470 & ~l1058;
assign a36868 = ~a36866 & ~a36864;
assign a36870 = ~l1470 & l1058;
assign a36872 = ~a36870 & ~a36868;
assign a36874 = a36872 & a36822;
assign a36876 = a12974 & ~a6254;
assign a36878 = ~a36876 & ~a36830;
assign a36880 = ~a36878 & ~a36826;
assign a36882 = ~a36880 & ~a36838;
assign a36884 = ~a36882 & ~a36834;
assign a36886 = ~a36884 & ~a36846;
assign a36888 = ~a36886 & ~a36842;
assign a36890 = ~a36888 & ~a36854;
assign a36892 = ~a36890 & ~a36850;
assign a36894 = ~a36892 & ~a36862;
assign a36896 = ~a36894 & ~a36858;
assign a36898 = ~a36896 & ~a36870;
assign a36900 = ~a36866 & ~a36822;
assign a36902 = a36900 & ~a36898;
assign a36904 = ~a36902 & ~a36874;
assign a36906 = ~l1328 & l978;
assign a36908 = l1328 & ~l978;
assign a36910 = ~a36908 & ~a36906;
assign a36912 = ~a12962 & a6254;
assign a36914 = ~a13146 & a6262;
assign a36916 = ~a36914 & ~a36912;
assign a36918 = a13146 & ~a6262;
assign a36920 = ~a36918 & ~a36916;
assign a36922 = ~a13336 & a6270;
assign a36924 = ~a36922 & ~a36920;
assign a36926 = a13336 & ~a6270;
assign a36928 = ~a36926 & ~a36924;
assign a36930 = ~a13526 & a6278;
assign a36932 = ~a36930 & ~a36928;
assign a36934 = a13526 & ~a6278;
assign a36936 = ~a36934 & ~a36932;
assign a36938 = ~a13716 & a6286;
assign a36940 = ~a36938 & ~a36936;
assign a36942 = a13716 & ~a6286;
assign a36944 = ~a36942 & ~a36940;
assign a36946 = ~a13894 & ~l1054;
assign a36948 = ~a36946 & ~a36944;
assign a36950 = a13894 & l1054;
assign a36952 = ~a36950 & ~a36948;
assign a36954 = ~a14058 & ~l1058;
assign a36956 = ~a36954 & ~a36952;
assign a36958 = a14058 & l1058;
assign a36960 = ~a36958 & ~a36956;
assign a36962 = ~a36960 & a36910;
assign a36964 = a12962 & ~a6254;
assign a36966 = ~a36964 & ~a36918;
assign a36968 = ~a36966 & ~a36914;
assign a36970 = ~a36968 & ~a36926;
assign a36972 = ~a36970 & ~a36922;
assign a36974 = ~a36972 & ~a36934;
assign a36976 = ~a36974 & ~a36930;
assign a36978 = ~a36976 & ~a36942;
assign a36980 = ~a36978 & ~a36938;
assign a36982 = ~a36980 & ~a36950;
assign a36984 = ~a36982 & ~a36946;
assign a36986 = ~a36984 & ~a36958;
assign a36988 = ~a36986 & ~a36954;
assign a36990 = ~a36988 & ~a36910;
assign a36992 = ~a36990 & ~a36962;
assign a36994 = a36992 & a5600;
assign a36996 = ~a36994 & ~a14558;
assign a36998 = ~a36996 & a36904;
assign a37000 = a36998 & a5594;
assign a37002 = ~a37000 & ~l886;
assign a37004 = ~a37002 & ~a36252;
assign a37006 = a36236 & l968;
assign a37008 = ~a37006 & ~a15734;
assign a37010 = ~a37008 & ~a36616;
assign a37012 = a37010 & l970;
assign a37014 = ~a37012 & ~l886;
assign a37016 = a36528 & l966;
assign a37018 = ~a37016 & ~a15398;
assign a37020 = ~a37018 & ~a36428;
assign a37022 = a37020 & l964;
assign a37024 = ~a37022 & ~l886;
assign a37026 = a36340 & l962;
assign a37028 = ~a37026 & ~a15066;
assign a37030 = ~a37028 & ~a36804;
assign a37032 = a37030 & l960;
assign a37034 = ~a37032 & ~l886;
assign a37036 = a36716 & a5606;
assign a37038 = ~a37036 & ~a14728;
assign a37040 = ~a37038 & ~a36992;
assign a37042 = a37040 & a5600;
assign a37044 = ~a37042 & ~l886;
assign a37046 = ~a36904 & a5594;
assign a37048 = ~a37046 & ~a16068;
assign a37050 = ~a37048 & ~a36144;
assign a37052 = a37050 & a5568;
assign a37054 = ~a37052 & ~l886;
assign a37056 = ~a36252 & ~a36242;
assign a37058 = ~a37056 & a37054;
assign a37060 = a37058 & a37044;
assign a37062 = a37060 & a37034;
assign a37064 = a37062 & a37024;
assign a37066 = a37064 & a37014;
assign a37068 = a37066 & ~a37004;
assign a37070 = a37068 & ~a36816;
assign a37072 = a37070 & ~a36628;
assign a37074 = a37072 & a36440;
assign a37076 = a37070 & ~a36440;
assign a37078 = a37076 & a36628;
assign a37080 = ~a37078 & ~a37074;
assign a37082 = ~a36628 & ~a36440;
assign a37084 = a37082 & ~a36816;
assign a37086 = a37084 & a37066;
assign a37088 = a37086 & a37004;
assign a37090 = ~a37044 & a36816;
assign a37092 = a37090 & a37004;
assign a37094 = a37092 & ~l2076;
assign a37096 = a37076 & ~a36628;
assign a37098 = a37096 & l2076;
assign a37100 = a37054 & ~a37004;
assign a37102 = a37024 & a37014;
assign a37104 = a37102 & a37084;
assign a37106 = a37104 & a37034;
assign a37108 = a37106 & a37044;
assign a37110 = a37108 & a37056;
assign a37112 = a37110 & a37100;
assign a37114 = a37082 & a37068;
assign a37116 = a37114 & a36816;
assign a37118 = ~a37116 & ~a37112;
assign a37120 = a37118 & ~a37098;
assign a37122 = a37120 & ~a37094;
assign a37124 = a37122 & ~a37088;
assign a37126 = a37124 & a37080;
assign a37128 = a37084 & ~a37004;
assign a37130 = a37128 & a37014;
assign a37132 = a37130 & a37024;
assign a37134 = a37132 & ~a37044;
assign a37136 = a37134 & a37058;
assign a37138 = a37136 & a37034;
assign a37140 = a37096 & l2078;
assign a37142 = l2078 & ~l2076;
assign a37144 = ~a37142 & ~a36244;
assign a37146 = ~a37144 & a37092;
assign a37148 = a37130 & ~a37024;
assign a37150 = a37148 & a37062;
assign a37152 = ~a37116 & ~a37078;
assign a37154 = a37152 & ~a37150;
assign a37156 = a37154 & ~a37146;
assign a37158 = a37156 & ~a37140;
assign a37160 = a37158 & ~a37138;
assign a37162 = a37128 & ~a37014;
assign a37164 = a37162 & a37064;
assign a37166 = l2078 & l2076;
assign a37168 = a37166 & l2082;
assign a37170 = ~a37168 & l2080;
assign a37172 = a37168 & ~l2080;
assign a37174 = ~a37172 & ~a37170;
assign a37176 = ~a37174 & a37092;
assign a37178 = a37096 & l2080;
assign a37180 = ~a37178 & ~a37112;
assign a37182 = a37180 & ~a37176;
assign a37184 = a37182 & ~a37164;
assign a37186 = a37132 & ~a37034;
assign a37188 = a37186 & a37060;
assign a37190 = a37096 & l2082;
assign a37192 = ~a37166 & l2082;
assign a37194 = a37166 & ~l2082;
assign a37196 = ~a37194 & ~a37192;
assign a37198 = ~a37196 & a37092;
assign a37200 = ~a37198 & ~a37150;
assign a37202 = a37200 & ~a37190;
assign a37204 = a37202 & ~a37188;
assign a37206 = a37204 & a37080;
assign a37208 = l2084 & ~l2074;
assign a37210 = ~a37208 & ~a36022;
assign a37212 = ~a37210 & a36026;
assign a37214 = a37210 & a36042;
assign a37216 = ~a36042 & l2084;
assign a37218 = ~a37216 & ~a37214;
assign a37220 = ~a37218 & ~a36026;
assign a37222 = ~a37220 & ~a37212;
assign a37224 = l2084 & l2074;
assign a37226 = ~a37224 & l2086;
assign a37228 = a37224 & ~l2086;
assign a37230 = ~a37228 & ~a37226;
assign a37232 = ~a37230 & a36026;
assign a37234 = ~a36036 & l2086;
assign a37236 = ~a37234 & ~a36038;
assign a37238 = ~a37236 & a36042;
assign a37240 = ~a36042 & l2086;
assign a37242 = ~a37240 & ~a37238;
assign a37244 = ~a37242 & ~a36026;
assign a37246 = ~a37244 & ~a37232;
assign a37248 = a37224 & l2086;
assign a37250 = ~a37248 & ~l2088;
assign a37252 = ~a37250 & a36026;
assign a37254 = ~a36040 & ~a36024;
assign a37256 = ~a37254 & a36042;
assign a37258 = ~a36046 & ~l2088;
assign a37260 = ~a37258 & ~a36042;
assign a37262 = ~a37260 & ~a37256;
assign a37264 = ~a37262 & a36020;
assign a37266 = ~a37264 & ~a37252;
assign a37268 = ~a37126 & l1560;
assign a37270 = a37126 & l1564;
assign a37272 = ~a37270 & ~a37268;
assign a37274 = ~a37272 & ~a37184;
assign a37276 = ~a37126 & l1548;
assign a37278 = a37126 & l1570;
assign a37280 = ~a37278 & ~a37276;
assign a37282 = ~a37280 & ~a37160;
assign a37284 = ~a37126 & l1572;
assign a37286 = a37126 & l1574;
assign a37288 = ~a37286 & ~a37284;
assign a37290 = ~a37288 & a37160;
assign a37292 = ~a37290 & ~a37282;
assign a37294 = ~a37292 & ~a37206;
assign a37296 = ~a37126 & l1576;
assign a37298 = a37126 & l1578;
assign a37300 = ~a37298 & ~a37296;
assign a37302 = ~a37300 & ~a37160;
assign a37304 = ~a37126 & l1580;
assign a37306 = a37126 & l1582;
assign a37308 = ~a37306 & ~a37304;
assign a37310 = ~a37308 & a37160;
assign a37312 = ~a37310 & ~a37302;
assign a37314 = ~a37312 & a37206;
assign a37316 = ~a37314 & ~a37294;
assign a37318 = ~a37316 & a37184;
assign a37320 = ~a37318 & ~a37274;
assign a37322 = ~a37320 & ~l886;
assign a37324 = l2076 & l1560;
assign a37326 = ~l2076 & l1564;
assign a37328 = ~a37326 & ~a37324;
assign a37330 = ~a37328 & l2080;
assign a37332 = l2076 & l1548;
assign a37334 = ~l2076 & l1570;
assign a37336 = ~a37334 & ~a37332;
assign a37338 = ~a37336 & l2078;
assign a37340 = l2076 & l1572;
assign a37342 = ~l2076 & l1574;
assign a37344 = ~a37342 & ~a37340;
assign a37346 = ~a37344 & ~l2078;
assign a37348 = ~a37346 & ~a37338;
assign a37350 = ~a37348 & l2082;
assign a37352 = l2076 & l1576;
assign a37354 = ~l2076 & l1578;
assign a37356 = ~a37354 & ~a37352;
assign a37358 = ~a37356 & l2078;
assign a37360 = l2076 & l1580;
assign a37362 = ~l2076 & l1582;
assign a37364 = ~a37362 & ~a37360;
assign a37366 = ~a37364 & ~l2078;
assign a37368 = ~a37366 & ~a37358;
assign a37370 = ~a37368 & ~l2082;
assign a37372 = ~a37370 & ~a37350;
assign a37374 = ~a37372 & ~l2080;
assign a37376 = ~a37374 & ~a37330;
assign a37378 = ~a37376 & ~a36248;
assign a37380 = a37376 & a36248;
assign a37382 = ~a37380 & ~a37378;
assign a37384 = ~a37382 & l886;
assign a37386 = ~a37384 & ~a37322;
assign a37388 = a36024 & ~a36020;
assign a37390 = a37388 & ~l2092;
assign a37392 = a36046 & ~l2092;
assign a37394 = ~a36046 & l2092;
assign a37396 = ~a37394 & ~a37392;
assign a37398 = ~a37396 & ~a37388;
assign a37400 = ~a37398 & ~a37390;
assign a37402 = ~a33538 & l884;
assign a37404 = a30140 & l2004;
assign a37406 = a30132 & l1524;
assign a37408 = a30182 & l1988;
assign a37410 = a30120 & l1990;
assign a37412 = a30170 & l1992;
assign a37414 = a30104 & l1994;
assign a37416 = a30096 & l1996;
assign a37418 = a30156 & l1998;
assign a37420 = a30930 & l2000;
assign a37422 = a30934 & l2002;
assign a37424 = ~a37422 & ~a37420;
assign a37426 = a37424 & ~a37418;
assign a37428 = a37426 & ~a37416;
assign a37430 = a37428 & ~a37414;
assign a37432 = a37430 & ~a37412;
assign a37434 = a37432 & ~a37410;
assign a37436 = a37434 & ~a37408;
assign a37438 = a37436 & ~a37406;
assign a37440 = a37438 & ~a37404;
assign a37442 = ~a37440 & a30066;
assign a37444 = a30062 & l2094;
assign a37446 = ~a37444 & ~a37442;
assign a37448 = a37446 & ~a37402;
assign a37450 = l2098 & l884;
assign a37452 = a34274 & l1554;
assign a37454 = ~a37452 & l2096;
assign a37456 = a37452 & ~l2096;
assign a37458 = ~a37456 & ~a37454;
assign a37460 = ~a37458 & a34242;
assign a37462 = a34240 & a34184;
assign a37464 = a37462 & ~l2096;
assign a37466 = ~a37462 & l2096;
assign a37468 = ~a37466 & ~a37464;
assign a37470 = ~a37468 & ~a34242;
assign a37472 = ~a37470 & ~a37460;
assign a37474 = ~a37472 & ~l884;
assign a37476 = ~a37474 & ~a37450;
assign a37478 = ~a33538 & a5360;
assign a37480 = ~a5360 & l2098;
assign a37482 = ~a37480 & ~a37478;
assign a37484 = ~l2102 & l890;
assign a37486 = i576 & ~i574;
assign a37488 = ~a37486 & ~i574;
assign a37490 = a37488 & i578;
assign a37492 = ~a37490 & a37488;
assign a37494 = ~a37492 & i554;
assign a37496 = a37492 & i554;
assign a37498 = a37496 & i580;
assign a37500 = ~a37498 & ~a37494;
assign a37502 = ~a37500 & i572;
assign a37504 = a37502 & ~i570;
assign a37506 = a37504 & ~i568;
assign a37508 = a37506 & ~i566;
assign a37510 = a37508 & i564;
assign a37512 = a37496 & ~i580;
assign a37514 = a37512 & i572;
assign a37516 = a37514 & ~i570;
assign a37518 = a37516 & ~i568;
assign a37520 = a37518 & ~i566;
assign a37522 = a37520 & i564;
assign a37524 = ~a37522 & ~a37510;
assign a37526 = ~a37524 & ~i562;
assign a37528 = a37508 & ~i564;
assign a37530 = a37528 & ~i562;
assign a37532 = a37530 & ~i584;
assign a37534 = a37520 & ~i564;
assign a37536 = a37534 & ~i562;
assign a37538 = ~a37536 & ~a37532;
assign a37540 = a37492 & ~i554;
assign a37542 = a37540 & i580;
assign a37544 = a37542 & i572;
assign a37546 = a37544 & ~i570;
assign a37548 = a37546 & ~i568;
assign a37550 = a37548 & ~i566;
assign a37552 = a37550 & ~i564;
assign a37554 = a37552 & ~i562;
assign a37556 = a37554 & i584;
assign a37558 = a37556 & ~i586;
assign a37560 = ~a37558 & a37538;
assign a37562 = ~a37560 & i582;
assign a37564 = ~a37562 & ~a37526;
assign a37566 = ~a37560 & ~i582;
assign a37568 = a37566 & ~i588;
assign a37570 = ~a37568 & a37564;
assign a37572 = ~a37492 & ~i554;
assign a37574 = a37540 & ~i580;
assign a37576 = ~a37574 & ~a37572;
assign a37578 = ~a37576 & i572;
assign a37580 = a37578 & ~i570;
assign a37582 = a37580 & ~i568;
assign a37584 = a37582 & ~i566;
assign a37586 = a37584 & i564;
assign a37588 = a37550 & i564;
assign a37590 = ~a37588 & ~a37586;
assign a37592 = ~a37590 & i562;
assign a37594 = a37592 & i586;
assign a37596 = a37584 & ~i564;
assign a37598 = a37596 & i562;
assign a37600 = a37598 & ~i584;
assign a37602 = a37552 & i562;
assign a37604 = ~a37602 & ~a37600;
assign a37606 = ~a37604 & i586;
assign a37608 = a37606 & i582;
assign a37610 = ~a37608 & ~a37594;
assign a37612 = a37606 & ~i582;
assign a37614 = a37612 & ~i588;
assign a37616 = ~a37614 & a37610;
assign a37618 = ~a37616 & ~i590;
assign a37620 = ~a37618 & a37570;
assign a37622 = ~a37620 & i560;
assign a37624 = a37622 & i592;
assign a37626 = a37624 & i594;
assign a37628 = a37626 & i596;
assign a37630 = a37622 & ~i592;
assign a37632 = a37630 & ~i594;
assign a37634 = a37632 & i596;
assign a37636 = ~a37634 & ~a37628;
assign a37638 = ~a37636 & i598;
assign a37640 = a37626 & ~i596;
assign a37642 = a37640 & ~i598;
assign a37644 = ~a37642 & ~a37638;
assign a37646 = ~a37644 & i600;
assign a37648 = a37632 & ~i596;
assign a37650 = a37648 & ~i598;
assign a37652 = a37650 & i600;
assign a37654 = ~a37652 & ~a37646;
assign a37656 = ~a37654 & i602;
assign a37658 = ~a37644 & ~i600;
assign a37660 = a37658 & ~i602;
assign a37662 = ~a37660 & ~a37656;
assign a37664 = ~a37616 & i590;
assign a37666 = a37664 & i560;
assign a37668 = a37666 & i592;
assign a37670 = a37668 & i594;
assign a37672 = a37670 & i596;
assign a37674 = a37666 & ~i592;
assign a37676 = a37674 & ~i594;
assign a37678 = a37676 & i596;
assign a37680 = ~a37678 & ~a37672;
assign a37682 = ~a37680 & i598;
assign a37684 = a37670 & ~i596;
assign a37686 = a37684 & ~i598;
assign a37688 = ~a37686 & ~a37682;
assign a37690 = ~a37688 & ~i600;
assign a37692 = a37690 & ~i602;
assign a37694 = ~a37692 & a37662;
assign a37696 = ~a37694 & i604;
assign a37698 = a37696 & i606;
assign a37700 = ~a37694 & ~i604;
assign a37702 = ~a37688 & i600;
assign a37704 = a37676 & ~i596;
assign a37706 = a37704 & ~i598;
assign a37708 = a37706 & i600;
assign a37710 = ~a37708 & ~a37702;
assign a37712 = ~a37710 & i602;
assign a37714 = a37712 & ~i604;
assign a37716 = ~a37714 & ~a37700;
assign a37718 = ~a37716 & ~i606;
assign a37720 = ~a37718 & ~a37698;
assign a37722 = a37650 & ~i600;
assign a37724 = a37722 & ~i602;
assign a37726 = a37706 & ~i600;
assign a37728 = a37726 & ~i602;
assign a37730 = ~a37728 & ~a37724;
assign a37732 = ~a37730 & i604;
assign a37734 = a37732 & i606;
assign a37736 = ~a37734 & a37720;
assign a37738 = a37598 & i584;
assign a37740 = a37738 & i586;
assign a37742 = a37612 & i588;
assign a37744 = ~a37742 & ~a37740;
assign a37746 = ~a37744 & i590;
assign a37748 = a37746 & ~i560;
assign a37750 = a37748 & i592;
assign a37752 = a37748 & ~i592;
assign a37754 = a37752 & i598;
assign a37756 = ~a37754 & ~a37750;
assign a37758 = ~a37756 & i602;
assign a37760 = a37752 & ~i598;
assign a37762 = a37760 & i602;
assign a37764 = ~a37762 & ~a37758;
assign a37766 = ~a37764 & i604;
assign a37768 = a37746 & i560;
assign a37770 = a37768 & i592;
assign a37772 = a37770 & ~i594;
assign a37774 = a37772 & ~i596;
assign a37776 = a37768 & ~i592;
assign a37778 = a37776 & ~i594;
assign a37780 = a37778 & ~i596;
assign a37782 = a37780 & i598;
assign a37784 = ~a37782 & ~a37774;
assign a37786 = ~a37784 & ~i600;
assign a37788 = a37786 & i602;
assign a37790 = a37780 & ~i598;
assign a37792 = a37790 & ~i600;
assign a37794 = a37792 & i602;
assign a37796 = ~a37794 & ~a37788;
assign a37798 = ~a37796 & i604;
assign a37800 = a37798 & ~i606;
assign a37802 = a37770 & i594;
assign a37804 = a37802 & i596;
assign a37806 = a37778 & i596;
assign a37808 = ~a37806 & ~a37804;
assign a37810 = ~a37808 & i598;
assign a37812 = a37802 & ~i596;
assign a37814 = a37812 & ~i598;
assign a37816 = ~a37814 & ~a37810;
assign a37818 = ~a37816 & i600;
assign a37820 = a37790 & i600;
assign a37822 = ~a37820 & ~a37818;
assign a37824 = ~a37822 & i602;
assign a37826 = a37824 & i604;
assign a37828 = a37826 & ~i606;
assign a37830 = ~a37816 & ~i600;
assign a37832 = a37830 & i602;
assign a37834 = a37812 & i598;
assign a37836 = a37772 & i596;
assign a37838 = ~a37836 & ~a37834;
assign a37840 = ~a37784 & i600;
assign a37842 = ~a37840 & a37838;
assign a37844 = ~a37842 & i602;
assign a37846 = ~a37844 & ~a37832;
assign a37848 = ~a37846 & i604;
assign a37850 = ~a37848 & ~a37828;
assign a37852 = a37798 & i606;
assign a37854 = ~a37852 & a37850;
assign a37856 = a37826 & i606;
assign a37858 = a37592 & ~i586;
assign a37860 = ~a37604 & ~i586;
assign a37862 = a37534 & i562;
assign a37864 = a37862 & i584;
assign a37866 = ~a37864 & ~a37860;
assign a37868 = ~a37866 & i582;
assign a37870 = ~a37868 & ~a37858;
assign a37872 = ~a37866 & ~i582;
assign a37874 = a37872 & ~i588;
assign a37876 = ~a37874 & a37870;
assign a37878 = ~a37876 & i590;
assign a37880 = a37878 & ~i560;
assign a37882 = a37880 & i592;
assign a37884 = a37880 & ~i592;
assign a37886 = a37884 & i598;
assign a37888 = ~a37886 & ~a37882;
assign a37890 = ~a37888 & i602;
assign a37892 = a37884 & ~i598;
assign a37894 = a37892 & i602;
assign a37896 = ~a37894 & ~a37890;
assign a37898 = ~a37896 & i604;
assign a37900 = a37878 & i560;
assign a37902 = a37900 & i592;
assign a37904 = a37902 & ~i594;
assign a37906 = a37904 & ~i596;
assign a37908 = a37900 & ~i592;
assign a37910 = a37908 & ~i594;
assign a37912 = a37910 & ~i596;
assign a37914 = a37912 & i598;
assign a37916 = ~a37914 & ~a37906;
assign a37918 = ~a37916 & ~i600;
assign a37920 = a37918 & i602;
assign a37922 = a37912 & ~i598;
assign a37924 = a37922 & ~i600;
assign a37926 = a37924 & i602;
assign a37928 = ~a37926 & ~a37920;
assign a37930 = ~a37928 & i604;
assign a37932 = a37930 & ~i606;
assign a37934 = a37902 & i594;
assign a37936 = a37934 & i596;
assign a37938 = a37910 & i596;
assign a37940 = ~a37938 & ~a37936;
assign a37942 = ~a37940 & i598;
assign a37944 = a37934 & ~i596;
assign a37946 = a37944 & ~i598;
assign a37948 = ~a37946 & ~a37942;
assign a37950 = ~a37948 & i600;
assign a37952 = a37922 & i600;
assign a37954 = ~a37952 & ~a37950;
assign a37956 = ~a37954 & i602;
assign a37958 = a37956 & i604;
assign a37960 = a37958 & ~i606;
assign a37962 = ~a37948 & ~i600;
assign a37964 = a37962 & i602;
assign a37966 = a37944 & i598;
assign a37968 = a37904 & i596;
assign a37970 = ~a37968 & ~a37966;
assign a37972 = ~a37916 & i600;
assign a37974 = ~a37972 & a37970;
assign a37976 = ~a37974 & i602;
assign a37978 = ~a37976 & ~a37964;
assign a37980 = ~a37978 & i604;
assign a37982 = ~a37980 & ~a37960;
assign a37984 = a37930 & i606;
assign a37986 = ~a37984 & a37982;
assign a37988 = a37958 & i606;
assign a37990 = a37664 & ~i560;
assign a37992 = a37990 & i592;
assign a37994 = a37990 & ~i592;
assign a37996 = a37994 & i598;
assign a37998 = ~a37996 & ~a37992;
assign a38000 = ~a37998 & i602;
assign a38002 = a37994 & ~i598;
assign a38004 = a38002 & i602;
assign a38006 = ~a38004 & ~a38000;
assign a38008 = ~a38006 & i604;
assign a38010 = a37668 & ~i594;
assign a38012 = a38010 & ~i596;
assign a38014 = a37704 & i598;
assign a38016 = ~a38014 & ~a38012;
assign a38018 = ~a38016 & ~i600;
assign a38020 = a38018 & i602;
assign a38022 = a37726 & i602;
assign a38024 = ~a38022 & ~a38020;
assign a38026 = ~a38024 & i604;
assign a38028 = a38026 & ~i606;
assign a38030 = ~a37680 & ~i598;
assign a38032 = a37674 & i594;
assign a38034 = ~a38032 & ~a38030;
assign a38036 = ~a37940 & ~i598;
assign a38038 = ~a38036 & a38034;
assign a38040 = a37908 & i594;
assign a38042 = ~a38040 & a38038;
assign a38044 = ~a38042 & i602;
assign a38046 = a38044 & i604;
assign a38048 = a37712 & i604;
assign a38050 = a38048 & ~i606;
assign a38052 = a37690 & i602;
assign a38054 = a37684 & i598;
assign a38056 = a38010 & i596;
assign a38058 = ~a38056 & ~a38054;
assign a38060 = ~a38016 & i600;
assign a38062 = ~a38060 & a38058;
assign a38064 = ~a38062 & i602;
assign a38066 = ~a38064 & ~a38052;
assign a38068 = ~a38066 & i604;
assign a38070 = ~a38068 & ~a38050;
assign a38072 = a38026 & i606;
assign a38074 = ~a38072 & a38070;
assign a38076 = a38048 & i606;
assign a38078 = ~a37524 & i562;
assign a38080 = a37528 & i562;
assign a38082 = ~a38080 & ~a38078;
assign a38084 = a37738 & ~i586;
assign a38086 = ~a38084 & a38082;
assign a38088 = a37872 & i588;
assign a38090 = ~a38088 & a38086;
assign a38092 = a37862 & ~i584;
assign a38094 = ~a38092 & a38090;
assign a38096 = ~a38094 & i590;
assign a38098 = a38096 & ~i560;
assign a38100 = a38098 & i592;
assign a38102 = a38098 & ~i592;
assign a38104 = a38102 & i598;
assign a38106 = ~a38104 & ~a38100;
assign a38108 = ~a38106 & i602;
assign a38110 = a38102 & ~i598;
assign a38112 = a38110 & i602;
assign a38114 = ~a38112 & ~a38108;
assign a38116 = ~a38114 & i604;
assign a38118 = a38096 & i560;
assign a38120 = a38118 & i592;
assign a38122 = a38120 & ~i594;
assign a38124 = a38122 & ~i596;
assign a38126 = a38118 & ~i592;
assign a38128 = a38126 & ~i594;
assign a38130 = a38128 & ~i596;
assign a38132 = a38130 & i598;
assign a38134 = ~a38132 & ~a38124;
assign a38136 = ~a38134 & ~i600;
assign a38138 = a38136 & i602;
assign a38140 = a38130 & ~i598;
assign a38142 = a38140 & ~i600;
assign a38144 = a38142 & i602;
assign a38146 = ~a38144 & ~a38138;
assign a38148 = ~a38146 & i604;
assign a38150 = a38148 & ~i606;
assign a38152 = a38120 & i594;
assign a38154 = a38152 & i596;
assign a38156 = a38128 & i596;
assign a38158 = ~a38156 & ~a38154;
assign a38160 = ~a38158 & ~i598;
assign a38162 = a38126 & i594;
assign a38164 = ~a38162 & ~a38160;
assign a38166 = ~a37808 & ~i598;
assign a38168 = ~a38166 & a38164;
assign a38170 = a37776 & i594;
assign a38172 = ~a38170 & a38168;
assign a38174 = ~a38172 & i602;
assign a38176 = a38174 & i604;
assign a38178 = ~a38158 & i598;
assign a38180 = a38152 & ~i596;
assign a38182 = a38180 & ~i598;
assign a38184 = ~a38182 & ~a38178;
assign a38186 = ~a38184 & i600;
assign a38188 = a38140 & i600;
assign a38190 = ~a38188 & ~a38186;
assign a38192 = ~a38190 & i602;
assign a38194 = a38192 & i604;
assign a38196 = a38194 & i606;
assign a38198 = a38194 & ~i606;
assign a38200 = ~a38184 & ~i600;
assign a38202 = a38200 & i602;
assign a38204 = a38180 & i598;
assign a38206 = a38122 & i596;
assign a38208 = ~a38206 & ~a38204;
assign a38210 = ~a38134 & i600;
assign a38212 = ~a38210 & a38208;
assign a38214 = ~a38212 & i602;
assign a38216 = ~a38214 & ~a38202;
assign a38218 = ~a38216 & i604;
assign a38220 = ~a38218 & ~a38198;
assign a38222 = a38148 & i606;
assign a38224 = ~a38222 & a38220;
assign a38226 = a38224 & ~a38196;
assign a38228 = a38226 & ~a38176;
assign a38230 = a38228 & ~a38150;
assign a38232 = a38230 & ~a38116;
assign a38234 = a38232 & ~a38076;
assign a38236 = a38234 & a38074;
assign a38238 = a38236 & ~a38046;
assign a38240 = a38238 & ~a38028;
assign a38242 = a38240 & ~a38008;
assign a38244 = a38242 & ~a37988;
assign a38246 = a38244 & a37986;
assign a38248 = a38246 & ~a37932;
assign a38250 = a38248 & ~a37898;
assign a38252 = a38250 & ~a37856;
assign a38254 = a38252 & a37854;
assign a38256 = a38254 & ~a37800;
assign a38258 = a38256 & ~a37766;
assign a38260 = a38258 & i608;
assign a38262 = a38260 & ~a37736;
assign a38264 = a38262 & i610;
assign a38266 = ~a38260 & ~a37736;
assign a38268 = ~a38266 & ~a38076;
assign a38270 = ~a38268 & ~i610;
assign a38272 = ~a38270 & ~a38264;
assign a38274 = ~a37730 & ~i604;
assign a38276 = a38274 & ~i606;
assign a38278 = a38276 & a38260;
assign a38280 = a38278 & i610;
assign a38282 = ~a38280 & a38272;
assign a38284 = a37956 & ~i604;
assign a38286 = a37962 & ~i602;
assign a38288 = ~a37876 & ~i590;
assign a38290 = a37548 & i566;
assign a38292 = a38290 & ~i564;
assign a38294 = a38292 & ~i562;
assign a38296 = a38294 & i584;
assign a38298 = a38296 & i586;
assign a38300 = a38298 & i582;
assign a38302 = ~a38300 & ~a38288;
assign a38304 = a38298 & ~i582;
assign a38306 = a38304 & ~i588;
assign a38308 = ~a38306 & a38302;
assign a38310 = ~a38308 & i560;
assign a38312 = a38310 & i592;
assign a38314 = a38312 & i594;
assign a38316 = a38314 & i596;
assign a38318 = a38310 & ~i592;
assign a38320 = a38318 & ~i594;
assign a38322 = a38320 & i596;
assign a38324 = ~a38322 & ~a38316;
assign a38326 = ~a38324 & i598;
assign a38328 = a38314 & ~i596;
assign a38330 = a38328 & ~i598;
assign a38332 = ~a38330 & ~a38326;
assign a38334 = ~a38332 & i600;
assign a38336 = a38320 & ~i596;
assign a38338 = a38336 & ~i598;
assign a38340 = a38338 & i600;
assign a38342 = ~a38340 & ~a38334;
assign a38344 = ~a38342 & i602;
assign a38346 = ~a38344 & ~a38286;
assign a38348 = ~a38332 & ~i600;
assign a38350 = a38348 & ~i602;
assign a38352 = ~a38350 & a38346;
assign a38354 = ~a38352 & ~i604;
assign a38356 = ~a38354 & ~a38284;
assign a38358 = ~a38356 & ~i606;
assign a38360 = ~a38352 & i604;
assign a38362 = a38360 & i606;
assign a38364 = ~a38362 & ~a38358;
assign a38366 = a37924 & ~i602;
assign a38368 = a38338 & ~i600;
assign a38370 = a38368 & ~i602;
assign a38372 = ~a38370 & ~a38366;
assign a38374 = ~a38372 & i604;
assign a38376 = a38374 & i606;
assign a38378 = ~a38376 & a38364;
assign a38380 = ~a38378 & a38260;
assign a38382 = a38380 & ~i610;
assign a38384 = ~a38382 & a37986;
assign a38386 = ~a37978 & ~i604;
assign a38388 = ~a38386 & a38384;
assign a38390 = a38360 & ~i606;
assign a38392 = ~a38390 & a38388;
assign a38394 = ~a37974 & ~i602;
assign a38396 = ~a38394 & a38392;
assign a38398 = ~a37928 & ~i604;
assign a38400 = a37918 & ~i602;
assign a38402 = ~a38400 & ~a38398;
assign a38404 = a38312 & ~i594;
assign a38406 = a38404 & ~i596;
assign a38408 = a38336 & i598;
assign a38410 = ~a38408 & ~a38406;
assign a38412 = ~a38410 & ~i600;
assign a38414 = ~a38412 & a38402;
assign a38416 = a38368 & i602;
assign a38418 = ~a38416 & a38414;
assign a38420 = ~a38418 & ~i606;
assign a38422 = ~a38420 & ~a37932;
assign a38424 = a38374 & ~i606;
assign a38426 = ~a38424 & a38422;
assign a38428 = ~a38426 & i610;
assign a38430 = ~a38428 & a38396;
assign a38432 = ~a38418 & i606;
assign a38434 = ~a38432 & a38430;
assign a38436 = a38348 & i602;
assign a38438 = ~a38436 & a38434;
assign a38440 = a38328 & i598;
assign a38442 = ~a38440 & a38438;
assign a38444 = a38404 & i596;
assign a38446 = ~a38444 & a38442;
assign a38448 = ~a38410 & i600;
assign a38450 = ~a38448 & a38446;
assign a38452 = ~a38378 & ~a38260;
assign a38454 = ~a38452 & ~a37988;
assign a38456 = ~a38454 & ~i610;
assign a38458 = a38380 & i610;
assign a38460 = ~a38458 & ~a38456;
assign a38462 = ~a38372 & ~i604;
assign a38464 = a38462 & ~i606;
assign a38466 = a38464 & a38260;
assign a38468 = a38466 & i610;
assign a38470 = ~a38468 & a38460;
assign a38472 = ~a38268 & i610;
assign a38474 = ~a37716 & i606;
assign a38476 = ~a38474 & ~a38472;
assign a38478 = ~a37654 & ~i602;
assign a38480 = ~a38478 & a38476;
assign a38482 = ~a37636 & ~i598;
assign a38484 = ~a38482 & a38480;
assign a38486 = a37630 & i594;
assign a38488 = ~a38486 & a38484;
assign a38490 = a38274 & i606;
assign a38492 = ~a38490 & a38488;
assign a38494 = a38276 & ~a38260;
assign a38496 = ~a37500 & ~i572;
assign a38498 = a38496 & i564;
assign a38500 = a38496 & ~i564;
assign a38502 = a38500 & ~i584;
assign a38504 = a37514 & i570;
assign a38506 = a37516 & i568;
assign a38508 = ~a38506 & ~a38504;
assign a38510 = a37518 & i566;
assign a38512 = ~a38510 & a38508;
assign a38514 = a37544 & i570;
assign a38516 = ~a38514 & a38512;
assign a38518 = a37546 & i568;
assign a38520 = ~a38518 & a38516;
assign a38522 = a37542 & ~i572;
assign a38524 = ~a38522 & a38520;
assign a38526 = ~a38524 & ~i564;
assign a38528 = a38292 & i562;
assign a38530 = ~a38528 & ~a38526;
assign a38532 = ~a38530 & i584;
assign a38534 = ~a38532 & ~a38502;
assign a38536 = a37512 & ~i572;
assign a38538 = a38536 & ~i564;
assign a38540 = ~a38538 & a38534;
assign a38542 = a38296 & ~i586;
assign a38544 = ~a38542 & a38540;
assign a38546 = a37556 & i586;
assign a38548 = ~a38546 & a38544;
assign a38550 = ~a38548 & i582;
assign a38552 = ~a38550 & ~a38498;
assign a38554 = ~a38548 & ~i582;
assign a38556 = a38554 & ~i588;
assign a38558 = ~a38556 & a38552;
assign a38560 = a38536 & i564;
assign a38562 = ~a38560 & a38558;
assign a38564 = ~a38562 & i560;
assign a38566 = a38564 & ~i594;
assign a38568 = a38566 & ~i596;
assign a38570 = a38568 & ~i600;
assign a38572 = a38570 & ~i606;
assign a38574 = ~a38572 & ~a38494;
assign a38576 = a38464 & ~a38260;
assign a38578 = ~a38576 & a38574;
assign a38580 = ~a38578 & i610;
assign a38582 = ~a38580 & a38492;
assign a38584 = a38564 & i594;
assign a38586 = ~a38584 & a38582;
assign a38588 = a38566 & i596;
assign a38590 = ~a38588 & a38586;
assign a38592 = a38568 & i600;
assign a38594 = ~a38592 & a38590;
assign a38596 = a38570 & i606;
assign a38598 = ~a38596 & a38594;
assign a38600 = ~a37710 & ~i602;
assign a38602 = ~a38600 & a38598;
assign a38604 = a38602 & ~a38046;
assign a38606 = a38044 & ~i604;
assign a38608 = ~a38606 & a38604;
assign a38610 = ~a38042 & ~i602;
assign a38612 = ~a38610 & a38608;
assign a38614 = ~a38454 & i610;
assign a38616 = ~a38614 & a38612;
assign a38618 = ~a38356 & i606;
assign a38620 = ~a38618 & a38616;
assign a38622 = ~a37954 & ~i602;
assign a38624 = ~a38622 & a38620;
assign a38626 = a38462 & i606;
assign a38628 = ~a38626 & a38624;
assign a38630 = ~a38342 & ~i602;
assign a38632 = ~a38630 & a38628;
assign a38634 = ~a38324 & ~i598;
assign a38636 = ~a38634 & a38632;
assign a38638 = a38318 & i594;
assign a38640 = ~a38638 & a38636;
assign a38642 = a38192 & ~i604;
assign a38644 = a38200 & ~i602;
assign a38646 = ~a38094 & ~i590;
assign a38648 = a37582 & i566;
assign a38650 = a38290 & i564;
assign a38652 = ~a38650 & ~a38648;
assign a38654 = ~a38652 & ~i562;
assign a38656 = a38294 & ~i584;
assign a38658 = ~a38656 & ~a38654;
assign a38660 = ~a38658 & i586;
assign a38662 = ~a38660 & ~a38646;
assign a38664 = a38304 & i588;
assign a38666 = ~a38664 & a38662;
assign a38668 = ~a38666 & i560;
assign a38670 = a38668 & i592;
assign a38672 = a38670 & i594;
assign a38674 = a38672 & i596;
assign a38676 = a38668 & ~i592;
assign a38678 = a38676 & ~i594;
assign a38680 = a38678 & i596;
assign a38682 = ~a38680 & ~a38674;
assign a38684 = ~a38682 & i598;
assign a38686 = a38672 & ~i596;
assign a38688 = a38686 & ~i598;
assign a38690 = ~a38688 & ~a38684;
assign a38692 = ~a38690 & i600;
assign a38694 = a38678 & ~i596;
assign a38696 = a38694 & ~i598;
assign a38698 = a38696 & i600;
assign a38700 = ~a38698 & ~a38692;
assign a38702 = ~a38700 & i602;
assign a38704 = ~a38702 & ~a38644;
assign a38706 = ~a38690 & ~i600;
assign a38708 = a38706 & ~i602;
assign a38710 = ~a38708 & a38704;
assign a38712 = ~a38710 & ~i604;
assign a38714 = ~a38712 & ~a38642;
assign a38716 = ~a38714 & ~i606;
assign a38718 = ~a38710 & i604;
assign a38720 = a38718 & i606;
assign a38722 = ~a38720 & ~a38716;
assign a38724 = a38142 & ~i602;
assign a38726 = a38696 & ~i600;
assign a38728 = a38726 & ~i602;
assign a38730 = ~a38728 & ~a38724;
assign a38732 = ~a38730 & i604;
assign a38734 = a38732 & i606;
assign a38736 = ~a38734 & a38722;
assign a38738 = ~a38736 & a38260;
assign a38740 = a38738 & ~i610;
assign a38742 = ~a38740 & a38224;
assign a38744 = ~a38216 & ~i604;
assign a38746 = ~a38744 & a38742;
assign a38748 = a38718 & ~i606;
assign a38750 = ~a38748 & a38746;
assign a38752 = ~a38212 & ~i602;
assign a38754 = ~a38752 & a38750;
assign a38756 = ~a38146 & ~i604;
assign a38758 = a38136 & ~i602;
assign a38760 = ~a38758 & ~a38756;
assign a38762 = a38670 & ~i594;
assign a38764 = a38762 & ~i596;
assign a38766 = a38694 & i598;
assign a38768 = ~a38766 & ~a38764;
assign a38770 = ~a38768 & ~i600;
assign a38772 = ~a38770 & a38760;
assign a38774 = a38726 & i602;
assign a38776 = ~a38774 & a38772;
assign a38778 = ~a38776 & ~i606;
assign a38780 = ~a38778 & ~a38150;
assign a38782 = a38732 & ~i606;
assign a38784 = ~a38782 & a38780;
assign a38786 = ~a38784 & i610;
assign a38788 = ~a38786 & a38754;
assign a38790 = ~a38776 & i606;
assign a38792 = ~a38790 & a38788;
assign a38794 = a38706 & i602;
assign a38796 = ~a38794 & a38792;
assign a38798 = a38686 & i598;
assign a38800 = ~a38798 & a38796;
assign a38802 = a38762 & i596;
assign a38804 = ~a38802 & a38800;
assign a38806 = ~a38768 & i600;
assign a38808 = ~a38806 & a38804;
assign a38810 = a37502 & i570;
assign a38812 = a37504 & i568;
assign a38814 = ~a38812 & ~a38810;
assign a38816 = a37506 & i566;
assign a38818 = ~a38816 & a38814;
assign a38820 = a38500 & i584;
assign a38822 = ~a38820 & a38818;
assign a38824 = a38554 & i588;
assign a38826 = ~a38824 & a38822;
assign a38828 = a37578 & i570;
assign a38830 = ~a38828 & a38826;
assign a38832 = a37580 & i568;
assign a38834 = ~a38832 & a38830;
assign a38836 = ~a38652 & i562;
assign a38838 = ~a38836 & a38834;
assign a38840 = ~a38658 & ~i586;
assign a38842 = ~a38840 & a38838;
assign a38844 = ~a37590 & ~i562;
assign a38846 = a37596 & ~i562;
assign a38848 = ~a38846 & ~a38844;
assign a38850 = a37554 & ~i584;
assign a38852 = ~a38850 & a38848;
assign a38854 = ~a38852 & i586;
assign a38856 = ~a38854 & a38842;
assign a38858 = ~a37576 & ~i572;
assign a38860 = ~a38858 & a38856;
assign a38862 = ~a38524 & i564;
assign a38864 = ~a38862 & a38860;
assign a38866 = ~a38530 & ~i584;
assign a38868 = ~a38866 & a38864;
assign a38870 = ~a38868 & i560;
assign a38872 = a38870 & i594;
assign a38874 = a38870 & ~i594;
assign a38876 = a38874 & i596;
assign a38878 = ~a38876 & ~a38872;
assign a38880 = a38874 & ~i596;
assign a38882 = a38880 & i600;
assign a38884 = ~a38882 & a38878;
assign a38886 = a38880 & ~i600;
assign a38888 = a38886 & i606;
assign a38890 = ~a38888 & a38884;
assign a38892 = a38886 & ~i606;
assign a38894 = ~a38730 & ~i604;
assign a38896 = a38894 & ~i606;
assign a38898 = a38896 & ~a38260;
assign a38900 = ~a38898 & ~a38892;
assign a38902 = a37530 & i584;
assign a38904 = a37566 & i588;
assign a38906 = ~a38904 & ~a38902;
assign a38908 = ~a38852 & ~i586;
assign a38910 = ~a38908 & a38906;
assign a38912 = ~a37744 & ~i590;
assign a38914 = ~a38912 & a38910;
assign a38916 = ~a38914 & i560;
assign a38918 = a38916 & ~i592;
assign a38920 = a38918 & ~i594;
assign a38922 = a38920 & ~i596;
assign a38924 = a38922 & ~i598;
assign a38926 = a38924 & ~i600;
assign a38928 = a38926 & ~i602;
assign a38930 = a37792 & ~i602;
assign a38932 = ~a38930 & ~a38928;
assign a38934 = ~a38932 & ~i604;
assign a38936 = a38934 & ~i606;
assign a38938 = a38936 & ~a38260;
assign a38940 = ~a38938 & a38900;
assign a38942 = ~a38940 & i610;
assign a38944 = ~a38942 & a38890;
assign a38946 = ~a38736 & ~a38260;
assign a38948 = ~a38946 & ~a38196;
assign a38950 = ~a38948 & i610;
assign a38952 = ~a38950 & a38944;
assign a38954 = ~a38714 & i606;
assign a38956 = ~a38954 & a38952;
assign a38958 = ~a38190 & ~i602;
assign a38960 = ~a38958 & a38956;
assign a38962 = a38960 & ~a38176;
assign a38964 = a38174 & ~i604;
assign a38966 = ~a38964 & a38962;
assign a38968 = ~a38172 & ~i602;
assign a38970 = ~a38968 & a38966;
assign a38972 = a38894 & i606;
assign a38974 = ~a38972 & a38970;
assign a38976 = ~a38700 & ~i602;
assign a38978 = ~a38976 & a38974;
assign a38980 = ~a38682 & ~i598;
assign a38982 = ~a38980 & a38978;
assign a38984 = a38676 & i594;
assign a38986 = ~a38984 & a38982;
assign a38988 = a38916 & i592;
assign a38990 = a38988 & i594;
assign a38992 = a38990 & i596;
assign a38994 = a38920 & i596;
assign a38996 = ~a38994 & ~a38992;
assign a38998 = ~a38996 & i598;
assign a39000 = a38990 & ~i596;
assign a39002 = a39000 & ~i598;
assign a39004 = ~a39002 & ~a38998;
assign a39006 = ~a39004 & i600;
assign a39008 = a38924 & i600;
assign a39010 = ~a39008 & ~a39006;
assign a39012 = ~a39010 & i602;
assign a39014 = ~a39004 & ~i600;
assign a39016 = a39014 & ~i602;
assign a39018 = ~a39016 & ~a39012;
assign a39020 = a37830 & ~i602;
assign a39022 = ~a39020 & a39018;
assign a39024 = ~a39022 & i604;
assign a39026 = a39024 & i606;
assign a39028 = ~a39022 & ~i604;
assign a39030 = a37824 & ~i604;
assign a39032 = ~a39030 & ~a39028;
assign a39034 = ~a39032 & ~i606;
assign a39036 = ~a39034 & ~a39026;
assign a39038 = ~a38932 & i604;
assign a39040 = a39038 & i606;
assign a39042 = ~a39040 & a39036;
assign a39044 = ~a39042 & ~a38260;
assign a39046 = ~a39044 & ~a37856;
assign a39048 = ~a39046 & i610;
assign a39050 = ~a39048 & a38986;
assign a39052 = ~a39032 & i606;
assign a39054 = ~a39052 & a39050;
assign a39056 = ~a39010 & ~i602;
assign a39058 = ~a39056 & a39054;
assign a39060 = ~a38996 & ~i598;
assign a39062 = ~a39060 & a39058;
assign a39064 = a38918 & i594;
assign a39066 = ~a39064 & a39062;
assign a39068 = a38934 & i606;
assign a39070 = ~a39068 & a39066;
assign a39072 = ~a37822 & ~i602;
assign a39074 = ~a39072 & a39070;
assign a39076 = ~a38948 & ~i610;
assign a39078 = a38738 & i610;
assign a39080 = ~a39078 & ~a39076;
assign a39082 = a38896 & a38260;
assign a39084 = a39082 & i610;
assign a39086 = ~a39084 & a39080;
assign a39088 = a39086 & a39074;
assign a39090 = a39088 & a38808;
assign a39092 = a39090 & a38640;
assign a39094 = a39092 & a38470;
assign a39096 = a39094 & a38450;
assign a39098 = ~a38426 & ~i610;
assign a39100 = a38466 & ~i610;
assign a39102 = ~a39100 & ~a39098;
assign a39104 = ~a38914 & ~i560;
assign a39106 = a39104 & i592;
assign a39108 = a39106 & i598;
assign a39110 = a39108 & i602;
assign a39112 = a39110 & i604;
assign a39114 = a39112 & a38260;
assign a39116 = a38988 & ~i594;
assign a39118 = a39116 & ~i596;
assign a39120 = a38922 & i598;
assign a39122 = ~a39120 & ~a39118;
assign a39124 = ~a39122 & ~i600;
assign a39126 = a38926 & i602;
assign a39128 = ~a39126 & ~a39124;
assign a39130 = ~a37796 & ~i604;
assign a39132 = ~a39130 & a39128;
assign a39134 = a37786 & ~i602;
assign a39136 = ~a39134 & a39132;
assign a39138 = ~a39136 & ~i606;
assign a39140 = a39038 & ~i606;
assign a39142 = ~a39140 & ~a39138;
assign a39144 = a39142 & ~a37800;
assign a39146 = ~a39144 & ~i610;
assign a39148 = a38936 & a38260;
assign a39150 = a39148 & ~i610;
assign a39152 = ~a39150 & ~a39146;
assign a39154 = ~a39042 & a38260;
assign a39156 = a39154 & ~i610;
assign a39158 = a39024 & ~i606;
assign a39160 = ~a39158 & ~a39156;
assign a39162 = a39014 & i602;
assign a39164 = ~a39162 & a39160;
assign a39166 = a39000 & i598;
assign a39168 = ~a39166 & a39164;
assign a39170 = a39116 & i596;
assign a39172 = ~a39170 & a39168;
assign a39174 = ~a39122 & i600;
assign a39176 = ~a39174 & a39172;
assign a39178 = ~a39136 & i606;
assign a39180 = ~a39178 & a39176;
assign a39182 = ~a39144 & i610;
assign a39184 = ~a39182 & a39180;
assign a39186 = a39184 & a37854;
assign a39188 = ~a37846 & ~i604;
assign a39190 = ~a39188 & a39186;
assign a39192 = ~a37842 & ~i602;
assign a39194 = ~a39192 & a39190;
assign a39196 = a39154 & i610;
assign a39198 = ~a39046 & ~i610;
assign a39200 = ~a39198 & ~a39196;
assign a39202 = a39148 & i610;
assign a39204 = ~a39202 & a39200;
assign a39206 = ~a37620 & ~i560;
assign a39208 = a39206 & i592;
assign a39210 = a39208 & i598;
assign a39212 = a39210 & i602;
assign a39214 = a39212 & i604;
assign a39216 = a39214 & a38260;
assign a39218 = ~a38578 & ~i610;
assign a39220 = a37624 & ~i594;
assign a39222 = a39220 & ~i596;
assign a39224 = a37648 & i598;
assign a39226 = ~a39224 & ~a39222;
assign a39228 = ~a39226 & ~i600;
assign a39230 = a37722 & i602;
assign a39232 = ~a39230 & ~a39228;
assign a39234 = ~a38024 & ~i604;
assign a39236 = ~a39234 & a39232;
assign a39238 = a38018 & ~i602;
assign a39240 = ~a39238 & a39236;
assign a39242 = ~a39240 & ~i606;
assign a39244 = a37732 & ~i606;
assign a39246 = ~a39244 & ~a39242;
assign a39248 = a39246 & ~a38028;
assign a39250 = ~a39248 & ~i610;
assign a39252 = a38278 & ~i610;
assign a39254 = ~a39252 & ~a39250;
assign a39256 = a38262 & ~i610;
assign a39258 = a37696 & ~i606;
assign a39260 = ~a39258 & ~a39256;
assign a39262 = a37658 & i602;
assign a39264 = ~a39262 & a39260;
assign a39266 = a37640 & i598;
assign a39268 = ~a39266 & a39264;
assign a39270 = a39220 & i596;
assign a39272 = ~a39270 & a39268;
assign a39274 = ~a39226 & i600;
assign a39276 = ~a39274 & a39272;
assign a39278 = ~a39240 & i606;
assign a39280 = ~a39278 & a39276;
assign a39282 = ~a39248 & i610;
assign a39284 = ~a39282 & a39280;
assign a39286 = a39284 & a38074;
assign a39288 = ~a38066 & ~i604;
assign a39290 = ~a39288 & a39286;
assign a39292 = ~a38062 & ~i602;
assign a39294 = ~a39292 & a39290;
assign a39296 = ~a38940 & ~i610;
assign a39298 = ~a38784 & ~i610;
assign a39300 = a39082 & ~i610;
assign a39302 = ~a39300 & ~a39298;
assign a39304 = a39302 & ~a39296;
assign a39306 = a39304 & a38282;
assign a39308 = a39306 & a39294;
assign a39310 = a39308 & a39254;
assign a39312 = a39310 & ~a39218;
assign a39314 = a39312 & ~a39216;
assign a39316 = a39314 & a39204;
assign a39318 = a39316 & a39194;
assign a39320 = a39318 & a39152;
assign a39322 = a39320 & ~a39114;
assign a39324 = a39322 & a39102;
assign a39326 = a39324 & a39096;
assign a39328 = a39326 & i612;
assign a39330 = ~a39328 & a39096;
assign a39332 = a39330 & ~a38282;
assign a39334 = ~a39330 & ~a38640;
assign a39336 = ~a39334 & ~a39332;
assign a39338 = a39214 & ~a38260;
assign a39340 = a39212 & ~i604;
assign a39342 = ~a39340 & ~a39338;
assign a39344 = a39210 & ~i602;
assign a39346 = ~a39344 & a39342;
assign a39348 = a39208 & ~i598;
assign a39350 = ~a39348 & a39346;
assign a39352 = a39206 & ~i592;
assign a39354 = a39352 & i598;
assign a39356 = ~a39354 & a39350;
assign a39358 = a39352 & ~i598;
assign a39360 = a39358 & i602;
assign a39362 = ~a39360 & a39356;
assign a39364 = a39358 & ~i602;
assign a39366 = a38002 & ~i602;
assign a39368 = ~a39366 & ~a39364;
assign a39370 = ~a39368 & i604;
assign a39372 = ~a39370 & a39362;
assign a39374 = a39372 & ~a38008;
assign a39376 = ~a38006 & ~i604;
assign a39378 = ~a39376 & a39374;
assign a39380 = ~a37998 & ~i602;
assign a39382 = ~a39380 & a39378;
assign a39384 = ~a39382 & ~a39330;
assign a39386 = ~a39384 & a39336;
assign a39388 = ~a39368 & ~i604;
assign a39390 = a39388 & a38260;
assign a39392 = a39390 & ~a39330;
assign a39394 = ~a39392 & a39386;
assign a39396 = a39388 & ~a38260;
assign a39398 = ~a38562 & ~i560;
assign a39400 = ~a39398 & ~a39396;
assign a39402 = a37892 & ~i602;
assign a39404 = ~a38308 & ~i560;
assign a39406 = a39404 & ~i592;
assign a39408 = a39406 & ~i598;
assign a39410 = a39408 & ~i602;
assign a39412 = ~a39410 & ~a39402;
assign a39414 = ~a39412 & ~i604;
assign a39416 = a39414 & ~a38260;
assign a39418 = ~a39416 & a39400;
assign a39420 = ~a39418 & ~a39330;
assign a39422 = ~a39420 & a39394;
assign a39424 = a39330 & ~a39194;
assign a39426 = a39330 & ~a39294;
assign a39428 = ~a39330 & ~a39074;
assign a39430 = ~a38868 & ~i560;
assign a39432 = a38110 & ~i602;
assign a39434 = ~a38666 & ~i560;
assign a39436 = a39434 & ~i592;
assign a39438 = a39436 & ~i598;
assign a39440 = a39438 & ~i602;
assign a39442 = ~a39440 & ~a39432;
assign a39444 = ~a39442 & ~i604;
assign a39446 = a39444 & ~a38260;
assign a39448 = ~a39446 & ~a39430;
assign a39450 = a39104 & ~i592;
assign a39452 = a39450 & ~i598;
assign a39454 = a39452 & ~i602;
assign a39456 = a37760 & ~i602;
assign a39458 = ~a39456 & ~a39454;
assign a39460 = ~a39458 & ~i604;
assign a39462 = a39460 & ~a38260;
assign a39464 = ~a39462 & a39448;
assign a39466 = ~a39464 & ~a39330;
assign a39468 = ~a39466 & ~a39428;
assign a39470 = a39330 & ~a39204;
assign a39472 = ~a39470 & a39468;
assign a39474 = a39112 & ~a38260;
assign a39476 = a39110 & ~i604;
assign a39478 = ~a39476 & ~a39474;
assign a39480 = a39108 & ~i602;
assign a39482 = ~a39480 & a39478;
assign a39484 = a39106 & ~i598;
assign a39486 = ~a39484 & a39482;
assign a39488 = a39450 & i598;
assign a39490 = ~a39488 & a39486;
assign a39492 = a39452 & i602;
assign a39494 = ~a39492 & a39490;
assign a39496 = ~a39458 & i604;
assign a39498 = ~a39496 & a39494;
assign a39500 = a39498 & ~a37766;
assign a39502 = ~a37764 & ~i604;
assign a39504 = ~a39502 & a39500;
assign a39506 = ~a37756 & ~i602;
assign a39508 = ~a39506 & a39504;
assign a39510 = ~a39508 & ~a39330;
assign a39512 = ~a39510 & a39472;
assign a39514 = a39460 & a38260;
assign a39516 = a39514 & ~a39330;
assign a39518 = ~a39516 & a39512;
assign a39520 = a39518 & a39422;
assign a39522 = a39520 & ~a39426;
assign a39524 = a39522 & ~a39424;
assign a39526 = a39404 & i592;
assign a39528 = a39526 & i598;
assign a39530 = a39528 & i602;
assign a39532 = a39530 & i604;
assign a39534 = a39532 & a38260;
assign a39536 = a39534 & ~a39330;
assign a39538 = ~a39330 & ~a38450;
assign a39540 = a39330 & ~a39102;
assign a39542 = ~a39540 & ~a39538;
assign a39544 = ~a37888 & ~i602;
assign a39546 = ~a39544 & a37896;
assign a39548 = ~a39412 & i604;
assign a39550 = ~a39548 & a39546;
assign a39552 = a39532 & ~a38260;
assign a39554 = ~a39552 & a39550;
assign a39556 = a39530 & ~i604;
assign a39558 = ~a39556 & a39554;
assign a39560 = a39528 & ~i602;
assign a39562 = ~a39560 & a39558;
assign a39564 = a39526 & ~i598;
assign a39566 = ~a39564 & a39562;
assign a39568 = a39406 & i598;
assign a39570 = ~a39568 & a39566;
assign a39572 = a39408 & i602;
assign a39574 = ~a39572 & a39570;
assign a39576 = ~a39574 & a39330;
assign a39578 = ~a39576 & a39542;
assign a39580 = a39414 & a38260;
assign a39582 = a39580 & a39330;
assign a39584 = ~a39582 & a39578;
assign a39586 = a39534 & a39330;
assign a39588 = ~a39586 & a39584;
assign a39590 = a39330 & ~a39152;
assign a39592 = a39330 & a39218;
assign a39594 = ~a39418 & a39330;
assign a39596 = ~a39594 & ~a39592;
assign a39598 = ~a39330 & ~a38470;
assign a39600 = ~a39598 & a39596;
assign a39602 = a39330 & ~a39254;
assign a39604 = a39434 & i592;
assign a39606 = a39604 & i598;
assign a39608 = a39606 & i602;
assign a39610 = a39608 & i604;
assign a39612 = a39610 & a38260;
assign a39614 = a39612 & ~a39330;
assign a39616 = a39330 & a39296;
assign a39618 = ~a39464 & a39330;
assign a39620 = ~a39618 & ~a39616;
assign a39622 = ~a39330 & ~a39086;
assign a39624 = ~a39622 & a39620;
assign a39626 = ~a39330 & ~a38808;
assign a39628 = a39330 & ~a39302;
assign a39630 = ~a39628 & ~a39626;
assign a39632 = ~a38106 & ~i602;
assign a39634 = ~a39632 & a38114;
assign a39636 = ~a39442 & i604;
assign a39638 = ~a39636 & a39634;
assign a39640 = a39610 & ~a38260;
assign a39642 = ~a39640 & a39638;
assign a39644 = a39608 & ~i604;
assign a39646 = ~a39644 & a39642;
assign a39648 = a39606 & ~i602;
assign a39650 = ~a39648 & a39646;
assign a39652 = a39604 & ~i598;
assign a39654 = ~a39652 & a39650;
assign a39656 = a39436 & i598;
assign a39658 = ~a39656 & a39654;
assign a39660 = a39438 & i602;
assign a39662 = ~a39660 & a39658;
assign a39664 = ~a39662 & a39330;
assign a39666 = ~a39664 & a39630;
assign a39668 = a39444 & a38260;
assign a39670 = a39668 & a39330;
assign a39672 = ~a39670 & a39666;
assign a39674 = a39612 & a39330;
assign a39676 = ~a39674 & a39672;
assign a39678 = a39676 & a39624;
assign a39680 = a39678 & ~a39614;
assign a39682 = a39680 & ~a39602;
assign a39684 = a39682 & a39600;
assign a39686 = a39684 & ~a39590;
assign a39688 = a39686 & a39588;
assign a39690 = a39688 & ~a39536;
assign a39692 = a39690 & a39524;
assign a39694 = a39692 & i614;
assign a39696 = ~a39694 & a39524;
assign a39698 = ~a39696 & ~a39422;
assign a39700 = a39696 & ~a39600;
assign a39702 = ~a39700 & ~a39698;
assign a39704 = a39390 & a39330;
assign a39706 = a39704 & ~a39696;
assign a39708 = ~a39706 & a39702;
assign a39710 = ~a39574 & ~a39330;
assign a39712 = a39710 & ~a39696;
assign a39714 = ~a39712 & a39708;
assign a39716 = a39580 & ~a39330;
assign a39718 = ~a39716 & a39714;
assign a39720 = a39696 & ~a39676;
assign a39722 = a39696 & ~a39588;
assign a39724 = ~a39722 & ~a39720;
assign a39726 = a39330 & a39114;
assign a39728 = ~a39508 & a39330;
assign a39730 = ~a39728 & ~a39726;
assign a39732 = ~a39730 & ~a39696;
assign a39734 = ~a39696 & a39424;
assign a39736 = a39696 & a39590;
assign a39738 = ~a39736 & ~a39734;
assign a39740 = ~a39730 & a39696;
assign a39742 = ~a39740 & a39738;
assign a39744 = a39514 & a39330;
assign a39746 = a39744 & a39696;
assign a39748 = ~a39746 & a39742;
assign a39750 = a39330 & a39216;
assign a39752 = ~a39382 & a39330;
assign a39754 = ~a39752 & ~a39750;
assign a39756 = ~a39754 & ~a39696;
assign a39758 = ~a39696 & a39426;
assign a39760 = a39696 & a39602;
assign a39762 = ~a39760 & ~a39758;
assign a39764 = ~a39754 & a39696;
assign a39766 = ~a39764 & a39762;
assign a39768 = a39704 & a39696;
assign a39770 = ~a39768 & a39766;
assign a39772 = ~a39696 & ~a39518;
assign a39774 = a39696 & ~a39624;
assign a39776 = ~a39774 & ~a39772;
assign a39778 = ~a39662 & ~a39330;
assign a39780 = a39778 & ~a39696;
assign a39782 = ~a39780 & a39776;
assign a39784 = a39668 & ~a39330;
assign a39786 = ~a39784 & a39782;
assign a39788 = a39744 & ~a39696;
assign a39790 = ~a39788 & a39786;
assign a39792 = a39790 & a39718;
assign a39794 = a39792 & a39770;
assign a39796 = a39794 & ~a39756;
assign a39798 = a39796 & a39748;
assign a39800 = a39798 & ~a39732;
assign a39802 = a39800 & a39724;
assign a39804 = a39802 & i616;
assign a39806 = ~a39804 & a39724;
assign a39808 = a39806 & ~a39718;
assign a39810 = ~a39806 & a39722;
assign a39812 = ~a39810 & ~a39808;
assign a39814 = a39710 & a39696;
assign a39816 = ~a39814 & a39812;
assign a39818 = a39696 & a39536;
assign a39820 = ~a39818 & a39816;
assign a39822 = a39806 & ~a39770;
assign a39824 = a39806 & ~a39748;
assign a39826 = ~a39824 & ~a39822;
assign a39828 = a39806 & ~a39790;
assign a39830 = ~a39806 & a39720;
assign a39832 = ~a39830 & ~a39828;
assign a39834 = a39778 & a39696;
assign a39836 = ~a39834 & a39832;
assign a39838 = a39696 & a39614;
assign a39840 = ~a39838 & a39836;
assign a39842 = a39840 & a39820;
assign a39844 = a39842 & a39826;
assign a39846 = a39844 & i618;
assign a39848 = ~a39846 & a39826;
assign a39850 = a39848 & ~a39820;
assign a39852 = ~a39848 & a39822;
assign a39854 = ~a39852 & ~a39850;
assign a39856 = a39806 & a39756;
assign a39858 = ~a39856 & a39854;
assign a39860 = a39858 & i558;
assign a39862 = ~i564 & ~i554;
assign a39864 = a39862 & i580;
assign a39866 = a39864 & i578;
assign a39868 = a39864 & ~i578;
assign a39870 = a39868 & i576;
assign a39872 = ~a39870 & ~a39866;
assign a39874 = a39868 & ~i576;
assign a39876 = a39874 & i574;
assign a39878 = ~a39876 & a39872;
assign a39880 = a39862 & ~i580;
assign a39882 = ~a39880 & a39878;
assign a39884 = ~a39882 & i572;
assign a39886 = a39884 & i568;
assign a39888 = a39884 & ~i568;
assign a39890 = a39888 & i570;
assign a39892 = ~a39890 & ~a39886;
assign a39894 = a39888 & ~i570;
assign a39896 = a39894 & i566;
assign a39898 = a39896 & i562;
assign a39900 = ~a39898 & a39892;
assign a39902 = a39900 & ~a38846;
assign a39904 = ~a39882 & ~i572;
assign a39906 = ~a39904 & a39902;
assign a39908 = a39874 & ~i574;
assign a39910 = a39908 & i572;
assign a39912 = a39910 & i568;
assign a39914 = a39910 & ~i568;
assign a39916 = a39914 & i570;
assign a39918 = ~a39916 & ~a39912;
assign a39920 = a39918 & ~a38528;
assign a39922 = a39920 & ~a37554;
assign a39924 = a39908 & ~i572;
assign a39926 = ~a39924 & a39922;
assign a39928 = ~a39926 & ~i584;
assign a39930 = ~a39928 & a39906;
assign a39932 = ~a39930 & ~i582;
assign a39934 = a39932 & i588;
assign a39936 = a39896 & ~i562;
assign a39938 = ~a39936 & ~a38656;
assign a39940 = ~a39938 & ~i582;
assign a39942 = a39940 & i588;
assign a39944 = a38296 & ~i582;
assign a39946 = a39944 & i588;
assign a39948 = ~a39946 & ~a39942;
assign a39950 = ~a39948 & a38260;
assign a39952 = a39950 & ~i622;
assign a39954 = ~a39952 & ~a39934;
assign a39956 = ~a39948 & ~a38260;
assign a39958 = ~a39956 & a39954;
assign a39960 = a37738 & ~i582;
assign a39962 = a39960 & i588;
assign a39964 = ~a37604 & ~i582;
assign a39966 = a39964 & i588;
assign a39968 = ~a39966 & ~a39962;
assign a39970 = ~a39968 & a38260;
assign a39972 = a39970 & i590;
assign a39974 = a39972 & i622;
assign a39976 = ~a39974 & a39958;
assign a39978 = ~a39968 & ~a38260;
assign a39980 = a39978 & i590;
assign a39982 = ~a39980 & a39976;
assign a39984 = a39978 & ~i590;
assign a39986 = a39984 & ~i604;
assign a39988 = a39986 & ~i602;
assign a39990 = ~a39988 & a39982;
assign a39992 = ~a39926 & i584;
assign a39994 = a39992 & ~i582;
assign a39996 = a39994 & i588;
assign a39998 = ~a39996 & a39990;
assign a40000 = a39970 & ~i590;
assign a40002 = a40000 & i622;
assign a40004 = ~a40002 & a39998;
assign a40006 = a39984 & i604;
assign a40008 = ~a40006 & a40004;
assign a40010 = a39986 & i602;
assign a40012 = ~a40010 & a40008;
assign a40014 = ~i564 & i554;
assign a40016 = a40014 & i580;
assign a40018 = a40014 & ~i580;
assign a40020 = a40018 & i578;
assign a40022 = ~a40020 & ~a40016;
assign a40024 = a40018 & ~i578;
assign a40026 = a40024 & i576;
assign a40028 = ~a40026 & a40022;
assign a40030 = a40024 & ~i576;
assign a40032 = a40030 & i574;
assign a40034 = ~a40032 & a40028;
assign a40036 = ~a40034 & i572;
assign a40038 = a40036 & i568;
assign a40040 = a40036 & ~i568;
assign a40042 = a40040 & i570;
assign a40044 = ~a40042 & ~a40038;
assign a40046 = a40040 & ~i570;
assign a40048 = a40046 & i566;
assign a40050 = a40048 & i562;
assign a40052 = ~a40050 & a40044;
assign a40054 = ~a38500 & ~a37530;
assign a40056 = ~a40054 & i584;
assign a40058 = ~a40056 & a40052;
assign a40060 = a40030 & ~i574;
assign a40062 = a40060 & i572;
assign a40064 = a40062 & i568;
assign a40066 = a40062 & ~i568;
assign a40068 = a40066 & i570;
assign a40070 = ~a40068 & ~a40064;
assign a40072 = a40066 & ~i570;
assign a40074 = a40072 & i566;
assign a40076 = a40074 & i562;
assign a40078 = ~a40076 & a40070;
assign a40080 = ~a40078 & ~i584;
assign a40082 = ~a40080 & a40058;
assign a40084 = ~a40082 & ~i582;
assign a40086 = a40084 & i588;
assign a40088 = a40048 & ~i562;
assign a40090 = a40074 & ~i562;
assign a40092 = a40090 & ~i584;
assign a40094 = ~a40092 & ~a40088;
assign a40096 = ~a40094 & ~i582;
assign a40098 = a40096 & i588;
assign a40100 = a40090 & i584;
assign a40102 = a40100 & ~i582;
assign a40104 = a40102 & i588;
assign a40106 = ~a40104 & ~a40098;
assign a40108 = ~a40106 & a38260;
assign a40110 = a40108 & ~i622;
assign a40112 = ~a40110 & ~a40086;
assign a40114 = ~a40106 & ~a38260;
assign a40116 = ~a40114 & a40112;
assign a40118 = ~a38092 & ~a38080;
assign a40120 = ~a40118 & ~i582;
assign a40122 = a40120 & i588;
assign a40124 = a37864 & ~i582;
assign a40126 = a40124 & i588;
assign a40128 = ~a40126 & ~a40122;
assign a40130 = ~a40128 & a38260;
assign a40132 = a40130 & i590;
assign a40134 = a40132 & i622;
assign a40136 = ~a40134 & a40116;
assign a40138 = ~a40128 & ~a38260;
assign a40140 = a40138 & i590;
assign a40142 = ~a40140 & a40136;
assign a40144 = a40138 & ~i590;
assign a40146 = a40144 & ~i604;
assign a40148 = a40146 & ~i602;
assign a40150 = ~a40148 & a40142;
assign a40152 = ~a40054 & ~i584;
assign a40154 = ~a40078 & i584;
assign a40156 = ~a40154 & ~a40152;
assign a40158 = a40156 & ~a37536;
assign a40160 = a40158 & ~a38538;
assign a40162 = ~a40160 & ~i582;
assign a40164 = a40162 & i588;
assign a40166 = ~a40164 & a40150;
assign a40168 = a40130 & ~i590;
assign a40170 = a40168 & i622;
assign a40172 = ~a40170 & a40166;
assign a40174 = a40144 & i604;
assign a40176 = ~a40174 & a40172;
assign a40178 = a40146 & i602;
assign a40180 = ~a40178 & a40176;
assign a40182 = i564 & i554;
assign a40184 = a40182 & ~i572;
assign a40186 = ~a40184 & ~a37526;
assign a40188 = ~a40160 & i582;
assign a40190 = ~a40188 & a40186;
assign a40192 = a40162 & ~i588;
assign a40194 = ~a40192 & a40190;
assign a40196 = a40100 & i582;
assign a40198 = a40102 & ~i588;
assign a40200 = ~a40198 & ~a40196;
assign a40202 = a38296 & i582;
assign a40204 = ~a40202 & a40200;
assign a40206 = a39944 & ~i588;
assign a40208 = ~a40206 & a40204;
assign a40210 = ~a40208 & a38260;
assign a40212 = a40210 & ~i622;
assign a40214 = ~a40212 & a40194;
assign a40216 = ~a40208 & ~a38260;
assign a40218 = ~a40216 & a40214;
assign a40220 = a37864 & i582;
assign a40222 = a40124 & ~i588;
assign a40224 = ~a40222 & ~a40220;
assign a40226 = a40224 & ~a37592;
assign a40228 = ~a37604 & i582;
assign a40230 = ~a40228 & a40226;
assign a40232 = a39964 & ~i588;
assign a40234 = ~a40232 & a40230;
assign a40236 = ~a40234 & a38260;
assign a40238 = a40236 & i590;
assign a40240 = a40238 & i622;
assign a40242 = ~a40240 & a40218;
assign a40244 = ~a40234 & ~a38260;
assign a40246 = a40244 & i590;
assign a40248 = ~a40246 & a40242;
assign a40250 = a40244 & ~i590;
assign a40252 = a40250 & ~i604;
assign a40254 = a40252 & ~i602;
assign a40256 = ~a40254 & a40248;
assign a40258 = a39992 & i582;
assign a40260 = ~a40258 & a40256;
assign a40262 = a39994 & ~i588;
assign a40264 = ~a40262 & a40260;
assign a40266 = a40236 & ~i590;
assign a40268 = a40266 & i622;
assign a40270 = ~a40268 & a40264;
assign a40272 = a40250 & i604;
assign a40274 = ~a40272 & a40270;
assign a40276 = a40252 & i602;
assign a40278 = ~a40276 & a40274;
assign a40280 = a40182 & i572;
assign a40282 = a40280 & i568;
assign a40284 = a40280 & ~i568;
assign a40286 = a40284 & i570;
assign a40288 = ~a40286 & ~a40282;
assign a40290 = a40284 & ~i570;
assign a40292 = a40290 & i566;
assign a40294 = i564 & ~i554;
assign a40296 = a40294 & i572;
assign a40298 = a40296 & ~i568;
assign a40300 = a40298 & ~i570;
assign a40302 = a40300 & i566;
assign a40304 = ~a40302 & ~a40292;
assign a40306 = ~a40304 & i562;
assign a40308 = ~a40306 & a40288;
assign a40310 = ~a40304 & ~i562;
assign a40312 = ~a40094 & i582;
assign a40314 = ~a40312 & ~a40310;
assign a40316 = a40096 & ~i588;
assign a40318 = ~a40316 & a40314;
assign a40320 = ~a39938 & i582;
assign a40322 = ~a40320 & a40318;
assign a40324 = a39940 & ~i588;
assign a40326 = ~a40324 & a40322;
assign a40328 = ~a40326 & a38260;
assign a40330 = a40328 & ~i622;
assign a40332 = ~a40330 & a40308;
assign a40334 = ~a40326 & ~a38260;
assign a40336 = ~a40334 & a40332;
assign a40338 = ~a40118 & i582;
assign a40340 = ~a40338 & ~a38078;
assign a40342 = a40120 & ~i588;
assign a40344 = ~a40342 & a40340;
assign a40346 = a37738 & i582;
assign a40348 = ~a40346 & a40344;
assign a40350 = a39960 & ~i588;
assign a40352 = ~a40350 & a40348;
assign a40354 = ~a40352 & a38260;
assign a40356 = a40354 & i590;
assign a40358 = a40356 & i622;
assign a40360 = ~a40358 & a40336;
assign a40362 = ~a40352 & ~a38260;
assign a40364 = a40362 & i590;
assign a40366 = ~a40364 & a40360;
assign a40368 = a40362 & ~i590;
assign a40370 = a40368 & ~i604;
assign a40372 = a40370 & ~i602;
assign a40374 = ~a40372 & a40366;
assign a40376 = ~a40082 & i582;
assign a40378 = ~a40376 & a40374;
assign a40380 = a40084 & ~i588;
assign a40382 = ~a40380 & a40378;
assign a40384 = a40296 & i568;
assign a40386 = ~a40384 & a40382;
assign a40388 = a40298 & i570;
assign a40390 = ~a40388 & a40386;
assign a40392 = a40390 & ~a38844;
assign a40394 = a40294 & ~i572;
assign a40396 = ~a40394 & a40392;
assign a40398 = ~a39930 & i582;
assign a40400 = ~a40398 & a40396;
assign a40402 = a39932 & ~i588;
assign a40404 = ~a40402 & a40400;
assign a40406 = a40354 & ~i590;
assign a40408 = a40406 & i622;
assign a40410 = ~a40408 & a40404;
assign a40412 = a40368 & i604;
assign a40414 = ~a40412 & a40410;
assign a40416 = a40370 & i602;
assign a40418 = ~a40416 & a40414;
assign a40420 = a40418 & a40278;
assign a40422 = a40420 & a40180;
assign a40424 = a40422 & a40012;
assign a40426 = a40424 & i620;
assign a40428 = ~a40426 & a39860;
assign a40430 = i572 & i570;
assign a40432 = i572 & i566;
assign a40434 = i572 & i562;
assign a40436 = i572 & i568;
assign a40438 = ~a40436 & i572;
assign a40440 = a40438 & ~a40434;
assign a40442 = a40440 & a40432;
assign a40444 = a40442 & ~a40430;
assign a40446 = a40444 & i604;
assign a40448 = a40446 & i622;
assign a40450 = a40438 & a40434;
assign a40452 = a40450 & ~a40432;
assign a40454 = a40452 & ~a40430;
assign a40456 = a40454 & i604;
assign a40458 = a40456 & ~i622;
assign a40460 = ~a40458 & ~a40448;
assign a40462 = a40460 & i624;
assign a40464 = ~a40462 & a40428;
assign a40466 = ~a40460 & ~i624;
assign a40468 = ~a40466 & a40464;
assign a40470 = a40444 & i602;
assign a40472 = a40470 & i622;
assign a40474 = a40454 & i602;
assign a40476 = a40474 & ~i622;
assign a40478 = ~a40476 & ~a40472;
assign a40480 = a40478 & i626;
assign a40482 = ~a40480 & a40468;
assign a40484 = ~a40478 & ~i626;
assign a40486 = ~a40484 & a40482;
assign a40488 = a40444 & i598;
assign a40490 = a40488 & i622;
assign a40492 = a40454 & i598;
assign a40494 = a40492 & ~i622;
assign a40496 = ~a40494 & ~a40490;
assign a40498 = a40496 & i628;
assign a40500 = ~a40498 & a40486;
assign a40502 = ~a40496 & ~i628;
assign a40504 = ~a40502 & a40500;
assign a40506 = a40444 & i592;
assign a40508 = a40506 & i622;
assign a40510 = a40454 & i592;
assign a40512 = a40510 & ~i622;
assign a40514 = ~a40512 & ~a40508;
assign a40516 = a40514 & i630;
assign a40518 = ~a40516 & a40504;
assign a40520 = ~a40514 & ~i630;
assign a40522 = ~a40520 & a40518;
assign a40524 = a40444 & i634;
assign a40526 = a40524 & i622;
assign a40528 = a40454 & i634;
assign a40530 = a40528 & ~i622;
assign a40532 = ~a40530 & ~a40526;
assign a40534 = a40532 & i632;
assign a40536 = ~a40534 & a40522;
assign a40538 = ~a40532 & ~i632;
assign a40540 = ~a40538 & a40536;
assign a40542 = a40444 & i638;
assign a40544 = a40542 & i622;
assign a40546 = a40454 & i638;
assign a40548 = a40546 & ~i622;
assign a40550 = ~a40548 & ~a40544;
assign a40552 = a40550 & i636;
assign a40554 = ~a40552 & a40540;
assign a40556 = ~a40550 & ~i636;
assign a40558 = ~a40556 & a40554;
assign a40560 = a40444 & i642;
assign a40562 = a40560 & i622;
assign a40564 = a40454 & i642;
assign a40566 = a40564 & ~i622;
assign a40568 = ~a40566 & ~a40562;
assign a40570 = a40568 & i640;
assign a40572 = ~a40570 & a40558;
assign a40574 = ~a40568 & ~i640;
assign a40576 = ~a40574 & a40572;
assign a40578 = i586 & ~i554;
assign a40580 = ~a40578 & a40444;
assign a40582 = ~a40436 & ~a40430;
assign a40584 = a40432 & ~a40430;
assign a40586 = ~a40584 & a40582;
assign a40588 = ~a40586 & i564;
assign a40590 = ~a40588 & a40580;
assign a40592 = a40590 & i622;
assign a40594 = ~a40578 & a40454;
assign a40596 = a40434 & ~a40430;
assign a40598 = a40596 & ~a40436;
assign a40600 = ~a40598 & a40586;
assign a40602 = ~a40600 & i564;
assign a40604 = ~a40602 & a40594;
assign a40606 = a40604 & ~i622;
assign a40608 = ~a40606 & ~a40592;
assign a40610 = ~a40608 & a40576;
assign a40612 = ~a40610 & i556;
assign a40614 = a40612 & ~i554;
assign a40616 = ~i556 & i552;
assign a40618 = ~a40616 & ~i556;
assign a40620 = a40618 & i644;
assign a40622 = ~a40620 & ~a40616;
assign a40624 = a40618 & i646;
assign a40626 = ~a40624 & a40610;
assign a40628 = a40626 & a40622;
assign a40630 = a40628 & i554;
assign a40632 = ~a40630 & ~a40614;
assign a40634 = a40632 & ~i552;
assign a40636 = a40624 & ~a40578;
assign a40638 = ~a40636 & a40634;
assign a40640 = ~a40638 & ~l890;
assign a40644 = ~l2104 & l890;
assign a40646 = ~l890 & ~i560;
assign a40648 = ~a40646 & ~a40644;
assign a40650 = ~a40648 & ~i652;
assign a40652 = ~l2108 & l890;
assign a40654 = i588 & ~i564;
assign a40656 = a40654 & ~i582;
assign a40658 = i584 & ~i564;
assign a40660 = ~a40658 & a40434;
assign a40662 = a40658 & i580;
assign a40664 = ~a40662 & ~a40660;
assign a40666 = ~a40664 & ~a40656;
assign a40668 = a40108 & i622;
assign a40670 = a40132 & ~i622;
assign a40672 = ~a40670 & ~a40668;
assign a40674 = a40672 & a40180;
assign a40676 = a40168 & ~i622;
assign a40678 = ~a40676 & a40674;
assign a40680 = ~a40678 & ~i660;
assign a40682 = a40680 & ~i658;
assign a40684 = a40682 & ~i656;
assign a40686 = a40684 & a39860;
assign a40688 = a39950 & i622;
assign a40690 = a39972 & ~i622;
assign a40692 = ~a40690 & ~a40688;
assign a40694 = a40692 & a40012;
assign a40696 = a40000 & ~i622;
assign a40698 = ~a40696 & a40694;
assign a40700 = ~a40698 & ~i660;
assign a40702 = a40700 & ~i658;
assign a40704 = a40702 & ~i656;
assign a40706 = a40704 & a39860;
assign a40708 = ~a40706 & ~a40686;
assign a40710 = a40708 & i662;
assign a40712 = ~a40710 & ~a40686;
assign a40714 = ~a40712 & a40656;
assign a40716 = ~a40714 & ~a40666;
assign a40718 = i666 & ~i582;
assign a40720 = a40718 & ~i664;
assign a40722 = ~a40720 & ~a40716;
assign a40724 = a40720 & i668;
assign a40726 = ~a40724 & ~a40722;
assign a40728 = a40726 & ~l890;
assign a40730 = ~a40728 & ~a40652;
assign a40732 = ~a40730 & ~a40642;
assign a40734 = a40730 & a40642;
assign a40736 = ~l2114 & l890;
assign a40738 = ~a40658 & a40432;
assign a40740 = a40658 & i576;
assign a40742 = ~a40740 & ~a40738;
assign a40744 = ~a40742 & ~a40656;
assign a40746 = a40656 & i658;
assign a40748 = ~a40746 & ~a40744;
assign a40750 = ~a40748 & ~a40720;
assign a40752 = a40720 & i682;
assign a40754 = ~a40752 & ~a40750;
assign a40756 = a40754 & ~l890;
assign a40758 = ~a40756 & ~a40736;
assign a40760 = ~l2116 & l890;
assign a40762 = ~a40658 & a40436;
assign a40764 = a40658 & i574;
assign a40766 = ~a40764 & ~a40762;
assign a40768 = ~a40766 & ~a40656;
assign a40770 = a40656 & i660;
assign a40772 = ~a40770 & ~a40768;
assign a40774 = ~a40658 & a40430;
assign a40776 = a40658 & i578;
assign a40778 = ~a40776 & ~a40774;
assign a40780 = ~a40778 & ~a40656;
assign a40782 = a40656 & i656;
assign a40784 = ~a40782 & ~a40780;
assign a40786 = a40784 & a40748;
assign a40788 = a40786 & a40772;
assign a40790 = a40716 & a40578;
assign a40792 = ~a40790 & a40788;
assign a40794 = ~a40716 & ~a40578;
assign a40796 = ~a40794 & a40792;
assign a40798 = a37768 & ~i686;
assign a40800 = a38310 & ~i686;
assign a40802 = a37900 & ~i686;
assign a40804 = a37666 & ~i686;
assign a40806 = a38564 & ~i686;
assign a40808 = a38916 & ~i686;
assign a40810 = a37622 & ~i686;
assign a40812 = a38668 & ~i686;
assign a40814 = a38870 & ~i686;
assign a40816 = a38118 & ~i686;
assign a40818 = ~a40816 & ~a40814;
assign a40820 = a40818 & ~a40812;
assign a40822 = a40820 & ~a40810;
assign a40824 = a40822 & ~a40808;
assign a40826 = a40824 & ~a40806;
assign a40828 = a40826 & ~a40804;
assign a40830 = a40828 & ~a40802;
assign a40832 = a40830 & ~a40800;
assign a40834 = a40832 & ~a40798;
assign a40836 = i688 & ~i560;
assign a40838 = ~a40836 & a40834;
assign a40840 = ~a40578 & a40528;
assign a40842 = a40578 & a40524;
assign a40844 = ~a40842 & ~a40840;
assign a40846 = a40844 & a40838;
assign a40848 = ~a40846 & a39696;
assign a40850 = ~a40844 & ~a40838;
assign a40852 = ~a40850 & ~a40848;
assign a40854 = a37768 & ~i690;
assign a40856 = a38310 & ~i690;
assign a40858 = a37900 & ~i690;
assign a40860 = a37666 & ~i690;
assign a40862 = a38564 & ~i690;
assign a40864 = a38916 & ~i690;
assign a40866 = a37622 & ~i690;
assign a40868 = a38668 & ~i690;
assign a40870 = a38870 & ~i690;
assign a40872 = a38118 & ~i690;
assign a40874 = ~a40872 & ~a40870;
assign a40876 = a40874 & ~a40868;
assign a40878 = a40876 & ~a40866;
assign a40880 = a40878 & ~a40864;
assign a40882 = a40880 & ~a40862;
assign a40884 = a40882 & ~a40860;
assign a40886 = a40884 & ~a40858;
assign a40888 = a40886 & ~a40856;
assign a40890 = a40888 & ~a40854;
assign a40892 = i692 & ~i560;
assign a40894 = ~a40892 & a40890;
assign a40896 = ~a40578 & a40546;
assign a40898 = a40578 & a40542;
assign a40900 = ~a40898 & ~a40896;
assign a40902 = a40900 & a40894;
assign a40904 = ~a40902 & ~a40852;
assign a40906 = ~a40900 & ~a40894;
assign a40908 = ~a40906 & ~a40904;
assign a40910 = a37768 & ~i694;
assign a40912 = a38310 & ~i694;
assign a40914 = a37900 & ~i694;
assign a40916 = a37666 & ~i694;
assign a40918 = a38564 & ~i694;
assign a40920 = a38916 & ~i694;
assign a40922 = a37622 & ~i694;
assign a40924 = a38668 & ~i694;
assign a40926 = a38870 & ~i694;
assign a40928 = a38118 & ~i694;
assign a40930 = ~a40928 & ~a40926;
assign a40932 = a40930 & ~a40924;
assign a40934 = a40932 & ~a40922;
assign a40936 = a40934 & ~a40920;
assign a40938 = a40936 & ~a40918;
assign a40940 = a40938 & ~a40916;
assign a40942 = a40940 & ~a40914;
assign a40944 = a40942 & ~a40912;
assign a40946 = a40944 & ~a40910;
assign a40948 = i696 & ~i560;
assign a40950 = ~a40948 & a40946;
assign a40952 = ~a40578 & a40564;
assign a40954 = a40578 & a40560;
assign a40956 = ~a40954 & ~a40952;
assign a40958 = a40956 & a40950;
assign a40960 = ~a40956 & ~a40950;
assign a40962 = ~a40960 & ~a40958;
assign a40964 = ~a40962 & a40908;
assign a40966 = ~a40964 & ~a40796;
assign a40968 = a40962 & ~a40902;
assign a40970 = ~a40850 & a39806;
assign a40972 = ~a40970 & ~a40846;
assign a40974 = ~a40972 & ~a40906;
assign a40976 = ~a40974 & a40968;
assign a40978 = ~a40976 & a40966;
assign a40980 = a40978 & a40604;
assign a40982 = ~a40980 & ~a40624;
assign a40984 = ~a40982 & a40578;
assign a40986 = a40628 & ~i554;
assign a40988 = ~a40986 & ~a40984;
assign a40990 = ~a40988 & ~l890;
assign a40992 = ~a40990 & ~a40760;
assign a40994 = ~a40992 & ~a40758;
assign a40996 = a40992 & a40758;
assign a40998 = ~l2118 & l890;
assign a41000 = ~a40784 & ~a40720;
assign a41002 = a40720 & i698;
assign a41004 = ~a41002 & ~a41000;
assign a41006 = a41004 & ~l890;
assign a41008 = ~a41006 & ~a40998;
assign a41010 = ~a41008 & l2120;
assign a41012 = a41008 & ~l2120;
assign a41014 = ~l2122 & l890;
assign a41016 = ~a40772 & ~a40720;
assign a41018 = a40720 & i702;
assign a41020 = ~a41018 & ~a41016;
assign a41022 = a41020 & ~l890;
assign a41024 = ~a41022 & ~a41014;
assign a41026 = ~a41024 & l2124;
assign a41028 = a41024 & ~l2124;
assign a41030 = ~a41028 & ~a41026;
assign a41032 = a41030 & ~a41012;
assign a41034 = a41032 & ~a41010;
assign a41036 = a41034 & ~a40996;
assign a41038 = a41036 & ~a40994;
assign a41040 = a41038 & ~a40734;
assign a41042 = a41040 & ~a40732;
assign a41044 = ~l2126 & l890;
assign a41046 = a40622 & i706;
assign a41048 = a40778 & a40766;
assign a41050 = a40778 & ~a40742;
assign a41052 = ~a41050 & a41048;
assign a41054 = ~a41052 & i582;
assign a41056 = ~a41054 & ~a40624;
assign a41058 = a40766 & a40658;
assign a41060 = a41058 & a40664;
assign a41062 = a41060 & ~a40742;
assign a41064 = a41062 & a40778;
assign a41066 = ~a41064 & ~a40590;
assign a41068 = ~a41066 & a41056;
assign a41070 = a41068 & ~i554;
assign a41072 = a40778 & ~a40664;
assign a41074 = a41072 & a40766;
assign a41076 = ~a41074 & a41052;
assign a41078 = ~a41076 & i582;
assign a41080 = ~a41078 & ~a40624;
assign a41082 = a41058 & ~a40664;
assign a41084 = a41082 & a40742;
assign a41086 = a41084 & a40778;
assign a41088 = ~a41086 & ~a40604;
assign a41090 = ~a41088 & a41080;
assign a41092 = a41090 & i554;
assign a41094 = ~a41092 & ~a41070;
assign a41096 = ~a41094 & ~a40610;
assign a41098 = a41050 & ~a40664;
assign a41100 = ~a41098 & a41048;
assign a41102 = ~a41100 & i582;
assign a41104 = ~a41102 & ~a40624;
assign a41106 = a41082 & ~a40742;
assign a41108 = a41106 & a40778;
assign a41110 = a40450 & a40432;
assign a41112 = a41110 & ~a40430;
assign a41114 = a41112 & ~a40578;
assign a41116 = a40584 & a40434;
assign a41118 = ~a41116 & a40582;
assign a41120 = ~a41118 & i564;
assign a41122 = ~a41120 & a41114;
assign a41124 = ~a41122 & ~a41108;
assign a41126 = ~a41124 & a41104;
assign a41128 = a41126 & ~i554;
assign a41130 = a41068 & i554;
assign a41132 = ~a41130 & ~a41128;
assign a41134 = ~a41132 & a40610;
assign a41136 = ~a41134 & ~a41096;
assign a41138 = ~a41136 & a41046;
assign a41140 = ~a41064 & a40560;
assign a41142 = a41064 & i710;
assign a41144 = ~a41142 & ~a41140;
assign a41146 = ~a41144 & ~i554;
assign a41148 = ~a41086 & a40564;
assign a41150 = a41086 & i710;
assign a41152 = ~a41150 & ~a41148;
assign a41154 = ~a41152 & i554;
assign a41156 = ~a41154 & ~a41146;
assign a41158 = ~a41156 & ~a40610;
assign a41160 = a41112 & i642;
assign a41162 = a41160 & ~a41108;
assign a41164 = a41108 & i710;
assign a41166 = ~a41164 & ~a41162;
assign a41168 = ~a41166 & ~i554;
assign a41170 = ~a41144 & i554;
assign a41172 = ~a41170 & ~a41168;
assign a41174 = ~a41172 & a40610;
assign a41176 = ~a41174 & ~a41158;
assign a41178 = ~a41176 & ~i708;
assign a41180 = ~a41178 & a41138;
assign a41182 = a41176 & i708;
assign a41184 = ~a41182 & a41180;
assign a41186 = ~a41064 & a40542;
assign a41188 = a41064 & i714;
assign a41190 = ~a41188 & ~a41186;
assign a41192 = ~a41190 & ~i554;
assign a41194 = ~a41086 & a40546;
assign a41196 = a41086 & i714;
assign a41198 = ~a41196 & ~a41194;
assign a41200 = ~a41198 & i554;
assign a41202 = ~a41200 & ~a41192;
assign a41204 = ~a41202 & ~a40610;
assign a41206 = a41112 & i638;
assign a41208 = a41206 & ~a41108;
assign a41210 = a41108 & i714;
assign a41212 = ~a41210 & ~a41208;
assign a41214 = ~a41212 & ~i554;
assign a41216 = ~a41190 & i554;
assign a41218 = ~a41216 & ~a41214;
assign a41220 = ~a41218 & a40610;
assign a41222 = ~a41220 & ~a41204;
assign a41224 = ~a41222 & ~i712;
assign a41226 = ~a41224 & a41184;
assign a41228 = a41222 & i712;
assign a41230 = ~a41228 & a41226;
assign a41232 = ~a41064 & a40524;
assign a41234 = a41064 & i718;
assign a41236 = ~a41234 & ~a41232;
assign a41238 = ~a41236 & ~i554;
assign a41240 = ~a41086 & a40528;
assign a41242 = a41086 & i718;
assign a41244 = ~a41242 & ~a41240;
assign a41246 = ~a41244 & i554;
assign a41248 = ~a41246 & ~a41238;
assign a41250 = ~a41248 & ~a40610;
assign a41252 = a41112 & i634;
assign a41254 = a41252 & ~a41108;
assign a41256 = a41108 & i718;
assign a41258 = ~a41256 & ~a41254;
assign a41260 = ~a41258 & ~i554;
assign a41262 = ~a41236 & i554;
assign a41264 = ~a41262 & ~a41260;
assign a41266 = ~a41264 & a40610;
assign a41268 = ~a41266 & ~a41250;
assign a41270 = ~a41268 & ~i716;
assign a41272 = ~a41270 & a41230;
assign a41274 = a41268 & i716;
assign a41276 = ~a41274 & a41272;
assign a41278 = ~a41064 & a40506;
assign a41280 = a41064 & i722;
assign a41282 = ~a41280 & ~a41278;
assign a41284 = ~a41282 & ~i554;
assign a41286 = ~a41086 & a40510;
assign a41288 = a41086 & i722;
assign a41290 = ~a41288 & ~a41286;
assign a41292 = ~a41290 & i554;
assign a41294 = ~a41292 & ~a41284;
assign a41296 = ~a41294 & ~a40610;
assign a41298 = a41112 & i592;
assign a41300 = a41298 & ~a41108;
assign a41302 = a41108 & i722;
assign a41304 = ~a41302 & ~a41300;
assign a41306 = ~a41304 & ~i554;
assign a41308 = ~a41282 & i554;
assign a41310 = ~a41308 & ~a41306;
assign a41312 = ~a41310 & a40610;
assign a41314 = ~a41312 & ~a41296;
assign a41316 = ~a41314 & ~i720;
assign a41318 = ~a41316 & a41276;
assign a41320 = a41314 & i720;
assign a41322 = ~a41320 & a41318;
assign a41324 = ~a41064 & a40488;
assign a41326 = a41064 & i726;
assign a41328 = ~a41326 & ~a41324;
assign a41330 = ~a41328 & ~i554;
assign a41332 = ~a41086 & a40492;
assign a41334 = a41086 & i726;
assign a41336 = ~a41334 & ~a41332;
assign a41338 = ~a41336 & i554;
assign a41340 = ~a41338 & ~a41330;
assign a41342 = ~a41340 & ~a40610;
assign a41344 = a41112 & i598;
assign a41346 = a41344 & ~a41108;
assign a41348 = a41108 & i726;
assign a41350 = ~a41348 & ~a41346;
assign a41352 = ~a41350 & ~i554;
assign a41354 = ~a41328 & i554;
assign a41356 = ~a41354 & ~a41352;
assign a41358 = ~a41356 & a40610;
assign a41360 = ~a41358 & ~a41342;
assign a41362 = ~a41360 & ~i724;
assign a41364 = ~a41362 & a41322;
assign a41366 = a41360 & i724;
assign a41368 = ~a41366 & a41364;
assign a41370 = ~a41064 & a40470;
assign a41372 = a41064 & i730;
assign a41374 = ~a41372 & ~a41370;
assign a41376 = ~a41374 & ~i554;
assign a41378 = ~a41086 & a40474;
assign a41380 = a41086 & i730;
assign a41382 = ~a41380 & ~a41378;
assign a41384 = ~a41382 & i554;
assign a41386 = ~a41384 & ~a41376;
assign a41388 = ~a41386 & ~a40610;
assign a41390 = a41112 & i602;
assign a41392 = a41390 & ~a41108;
assign a41394 = a41108 & i730;
assign a41396 = ~a41394 & ~a41392;
assign a41398 = ~a41396 & ~i554;
assign a41400 = ~a41374 & i554;
assign a41402 = ~a41400 & ~a41398;
assign a41404 = ~a41402 & a40610;
assign a41406 = ~a41404 & ~a41388;
assign a41408 = ~a41406 & ~i728;
assign a41410 = ~a41408 & a41368;
assign a41412 = a41406 & i728;
assign a41414 = ~a41412 & a41410;
assign a41416 = ~a41064 & a40446;
assign a41418 = a41064 & i734;
assign a41420 = ~a41418 & ~a41416;
assign a41422 = ~a41420 & ~i554;
assign a41424 = ~a41086 & a40456;
assign a41426 = a41086 & i734;
assign a41428 = ~a41426 & ~a41424;
assign a41430 = ~a41428 & i554;
assign a41432 = ~a41430 & ~a41422;
assign a41434 = ~a41432 & ~a40610;
assign a41436 = a41112 & i604;
assign a41438 = a41436 & ~a41108;
assign a41440 = a41108 & i734;
assign a41442 = ~a41440 & ~a41438;
assign a41444 = ~a41442 & ~i554;
assign a41446 = ~a41420 & i554;
assign a41448 = ~a41446 & ~a41444;
assign a41450 = ~a41448 & a40610;
assign a41452 = ~a41450 & ~a41434;
assign a41454 = ~a41452 & ~i732;
assign a41456 = ~a41454 & a41414;
assign a41458 = a41452 & i732;
assign a41460 = ~a41458 & a41456;
assign a41462 = a40444 & a38260;
assign a41464 = a41462 & ~a41064;
assign a41466 = a41064 & i738;
assign a41468 = ~a41466 & ~a41464;
assign a41470 = ~a41468 & ~i554;
assign a41472 = a40454 & a38260;
assign a41474 = a41472 & ~a41086;
assign a41476 = a41086 & i738;
assign a41478 = ~a41476 & ~a41474;
assign a41480 = ~a41478 & i554;
assign a41482 = ~a41480 & ~a41470;
assign a41484 = ~a41482 & ~a40610;
assign a41486 = a41112 & a38260;
assign a41488 = a41486 & ~a41108;
assign a41490 = a41108 & i738;
assign a41492 = ~a41490 & ~a41488;
assign a41494 = ~a41492 & ~i554;
assign a41496 = ~a41468 & i554;
assign a41498 = ~a41496 & ~a41494;
assign a41500 = ~a41498 & a40610;
assign a41502 = ~a41500 & ~a41484;
assign a41504 = ~a41502 & ~i736;
assign a41506 = ~a41504 & a41460;
assign a41508 = a41502 & i736;
assign a41510 = ~a41508 & a41506;
assign a41512 = ~a41510 & ~l890;
assign a41514 = ~a41512 & ~a41044;
assign a41516 = a41514 & ~a41042;
assign a41518 = ~a41516 & ~i654;
assign a41520 = a41518 & a40650;
assign a41522 = a41520 & ~a40642;
assign a41524 = ~a40648 & ~i654;
assign a41526 = a41524 & a41516;
assign a41528 = a41526 & a40642;
assign a41530 = a40650 & i862;
assign a41532 = a41530 & ~l2410;
assign a41534 = l2428 & i652;
assign a41536 = a40650 & ~i862;
assign a41538 = a41536 & i654;
assign a41540 = a41538 & l2410;
assign a41542 = ~l2310 & l890;
assign a41544 = a40440 & ~a40432;
assign a41546 = a41544 & ~a40430;
assign a41548 = a41546 & ~a40578;
assign a41550 = a41546 & i642;
assign a41552 = a41550 & ~a40578;
assign a41554 = a40578 & a40564;
assign a41556 = ~a41554 & ~a41552;
assign a41558 = a41556 & a40950;
assign a41560 = ~a41556 & ~a40950;
assign a41562 = ~a41560 & ~a41558;
assign a41564 = a41546 & i634;
assign a41566 = a41564 & ~a40578;
assign a41568 = a40578 & a40528;
assign a41570 = ~a41568 & ~a41566;
assign a41572 = ~a41570 & ~a40838;
assign a41574 = ~a41572 & a39848;
assign a41576 = a41570 & a40838;
assign a41578 = ~a41576 & ~a41574;
assign a41580 = a41546 & i638;
assign a41582 = a41580 & ~a40578;
assign a41584 = a40578 & a40546;
assign a41586 = ~a41584 & ~a41582;
assign a41588 = ~a41586 & ~a40894;
assign a41590 = ~a41588 & ~a41578;
assign a41592 = ~a41590 & a41562;
assign a41594 = a41586 & a40894;
assign a41596 = ~a41594 & a41592;
assign a41598 = ~a41588 & ~a41562;
assign a41600 = ~a41576 & a39330;
assign a41602 = ~a41600 & ~a41572;
assign a41604 = ~a41602 & ~a41594;
assign a41606 = ~a41604 & a41598;
assign a41608 = ~a41606 & ~a41596;
assign a41610 = ~a41608 & ~a40624;
assign a41612 = a41610 & a41548;
assign a41614 = ~a41612 & a40982;
assign a41616 = a41614 & a40578;
assign a41618 = ~a41616 & ~a41612;
assign a41620 = ~a40982 & ~a40578;
assign a41622 = ~a41620 & a41618;
assign a41624 = ~a41622 & ~l890;
assign a41626 = ~a41624 & ~a41542;
assign a41628 = a41626 & a40648;
assign a41630 = ~a41628 & ~a41540;
assign a41632 = a41630 & ~a41534;
assign a41634 = a41632 & ~a41532;
assign a41636 = a41634 & ~a41528;
assign a41640 = ~l2106 & l890;
assign a41642 = ~l890 & ~i648;
assign a41646 = ~l2110 & l890;
assign a41648 = i672 & ~i664;
assign a41650 = a41648 & ~i670;
assign a41652 = ~a41650 & ~l890;
assign a41656 = ~a41654 & a40730;
assign a41658 = a41654 & i680;
assign a41660 = ~a41658 & ~a41656;
assign a41662 = ~l2112 & l890;
assign a41664 = i676 & ~i670;
assign a41666 = ~a41664 & ~l890;
assign a41668 = ~a41666 & ~a41662;
assign a41674 = ~a41654 & a40758;
assign a41676 = a41654 & i684;
assign a41678 = ~a41676 & ~a41674;
assign a41680 = a41520 & ~a40992;
assign a41682 = ~a40992 & a40642;
assign a41684 = a40992 & ~a40642;
assign a41686 = a41684 & ~l2124;
assign a41688 = ~a41686 & ~a41682;
assign a41690 = ~a41688 & a41526;
assign a41692 = ~l2414 & l2410;
assign a41694 = a41692 & ~l2418;
assign a41696 = l2414 & ~l2410;
assign a41698 = ~a41696 & ~a41694;
assign a41700 = ~a41698 & a41530;
assign a41702 = l2426 & i652;
assign a41704 = a41538 & l2414;
assign a41706 = ~l2316 & l890;
assign a41708 = a40984 & ~l890;
assign a41710 = ~a41708 & ~a41706;
assign a41712 = ~a41710 & a41626;
assign a41714 = ~l2314 & l890;
assign a41716 = a41612 & ~l890;
assign a41718 = ~a41716 & ~a41714;
assign a41720 = a41710 & ~a41626;
assign a41722 = a41720 & a41718;
assign a41724 = ~a41722 & ~a41712;
assign a41726 = ~a41724 & a40648;
assign a41728 = ~a41726 & ~a41704;
assign a41730 = a41728 & ~a41702;
assign a41732 = a41730 & ~a41700;
assign a41734 = a41732 & ~a41690;
assign a41738 = ~a41654 & a41008;
assign a41740 = a41654 & i700;
assign a41742 = ~a41740 & ~a41738;
assign a41744 = a41520 & l2120;
assign a41746 = a40992 & l2120;
assign a41748 = ~a40992 & ~a40642;
assign a41750 = a41748 & ~l2120;
assign a41752 = a40642 & l2120;
assign a41754 = ~a41752 & ~a41750;
assign a41756 = a41754 & ~a41746;
assign a41758 = ~a41756 & a41526;
assign a41760 = ~l2414 & l2406;
assign a41762 = ~l2410 & l2406;
assign a41764 = l2414 & l2410;
assign a41766 = a41764 & ~l2406;
assign a41768 = ~a41766 & ~a41762;
assign a41770 = a41768 & ~a41760;
assign a41772 = ~a41770 & a41530;
assign a41774 = l2424 & i652;
assign a41776 = a41538 & l2406;
assign a41778 = ~a41710 & ~a41626;
assign a41780 = a41778 & ~l2318;
assign a41782 = a41626 & l2318;
assign a41784 = ~a41782 & ~a41780;
assign a41786 = a41710 & l2318;
assign a41788 = ~a41786 & a41784;
assign a41790 = ~a41788 & a40648;
assign a41792 = ~a41790 & ~a41776;
assign a41794 = a41792 & ~a41774;
assign a41796 = a41794 & ~a41772;
assign a41798 = a41796 & ~a41758;
assign a41800 = a41798 & ~a41744;
assign a41802 = ~a41654 & a41024;
assign a41804 = a41654 & i704;
assign a41806 = ~a41804 & ~a41802;
assign a41808 = a41520 & l2124;
assign a41810 = a41748 & l2120;
assign a41812 = a40642 & l2124;
assign a41814 = ~a41812 & ~a41810;
assign a41816 = ~a41814 & a41526;
assign a41818 = a41764 & l2406;
assign a41820 = l2418 & ~l2410;
assign a41822 = ~a41820 & ~a41818;
assign a41824 = ~a41822 & a41530;
assign a41826 = l2422 & i652;
assign a41828 = a41538 & l2418;
assign a41830 = ~a41718 & a41626;
assign a41832 = a41778 & l2318;
assign a41834 = ~a41832 & ~a41830;
assign a41836 = ~a41834 & a40648;
assign a41838 = ~a41836 & ~a41828;
assign a41840 = a41838 & ~a41826;
assign a41842 = a41840 & ~a41824;
assign a41844 = a41842 & ~a41816;
assign a41846 = a41844 & ~a41808;
assign a41848 = ~l2128 & l890;
assign a41850 = a41060 & a40742;
assign a41852 = a41850 & a40778;
assign a41854 = a41546 & a38260;
assign a41856 = a41854 & ~a41852;
assign a41858 = a41852 & i738;
assign a41860 = ~a41858 & ~a41856;
assign a41862 = a40772 & a40656;
assign a41864 = a41862 & a40716;
assign a41866 = a41864 & a40748;
assign a41868 = a41866 & a40784;
assign a41870 = ~a41868 & ~a41860;
assign a41872 = a41868 & i742;
assign a41874 = ~a41872 & ~a41870;
assign a41876 = ~a41874 & ~l890;
assign a41878 = ~a41876 & ~a41848;
assign a41880 = a40992 & ~l2120;
assign a41882 = a41880 & ~a41878;
assign a41884 = a41882 & l2124;
assign a41886 = a41884 & ~a40642;
assign a41888 = ~l2132 & l890;
assign a41890 = a40778 & a40742;
assign a41892 = a41890 & ~a40766;
assign a41894 = a41892 & a40658;
assign a41896 = a41894 & ~a40664;
assign a41898 = ~a40432 & ~a40430;
assign a41900 = a41898 & a40436;
assign a41902 = a41900 & a40434;
assign a41904 = a41902 & a38260;
assign a41906 = a41904 & ~a41896;
assign a41908 = a41896 & i738;
assign a41910 = ~a41908 & ~a41906;
assign a41912 = a40786 & ~a40772;
assign a41914 = a41912 & a40656;
assign a41916 = a41914 & ~a40716;
assign a41918 = ~a41916 & ~a41910;
assign a41920 = a41916 & i742;
assign a41922 = ~a41920 & ~a41918;
assign a41924 = ~a41922 & ~l890;
assign a41926 = ~a41924 & ~a41888;
assign a41928 = a41880 & l2124;
assign a41930 = a41928 & ~a41926;
assign a41932 = a41930 & a40642;
assign a41934 = ~l2134 & l890;
assign a41936 = a41900 & ~a40434;
assign a41938 = a41936 & a38260;
assign a41940 = a41894 & a40664;
assign a41942 = ~a41940 & a41938;
assign a41944 = a41940 & i738;
assign a41946 = ~a41944 & ~a41942;
assign a41948 = a41914 & a40716;
assign a41950 = ~a41948 & ~a41946;
assign a41952 = a41948 & i742;
assign a41954 = ~a41952 & ~a41950;
assign a41956 = ~a41954 & ~l890;
assign a41958 = ~a41956 & ~a41934;
assign a41960 = ~l2124 & l2120;
assign a41962 = a41960 & ~a40992;
assign a41964 = a41962 & ~a41958;
assign a41966 = a41964 & ~a40642;
assign a41968 = ~l2136 & l890;
assign a41970 = a41110 & a40430;
assign a41972 = a41970 & a38260;
assign a41974 = a41106 & ~a40778;
assign a41976 = ~a41974 & a41972;
assign a41978 = a41974 & i738;
assign a41980 = ~a41978 & ~a41976;
assign a41982 = a41862 & ~a40716;
assign a41984 = a41982 & ~a40748;
assign a41986 = a41984 & ~a40784;
assign a41988 = ~a41986 & ~a41980;
assign a41990 = a41986 & i742;
assign a41992 = ~a41990 & ~a41988;
assign a41994 = ~a41992 & ~l890;
assign a41996 = ~a41994 & ~a41968;
assign a41998 = ~a41996 & a41960;
assign a42000 = a41998 & ~a40992;
assign a42002 = a42000 & a40642;
assign a42004 = ~l2138 & l890;
assign a42006 = a40442 & a40430;
assign a42008 = a42006 & a38260;
assign a42010 = a41062 & ~a40778;
assign a42012 = ~a42010 & a42008;
assign a42014 = a42010 & i738;
assign a42016 = ~a42014 & ~a42012;
assign a42018 = a41864 & ~a40748;
assign a42020 = a42018 & ~a40784;
assign a42022 = ~a42020 & ~a42016;
assign a42024 = a42020 & i742;
assign a42026 = ~a42024 & ~a42022;
assign a42028 = ~a42026 & ~l890;
assign a42030 = ~a42028 & ~a42004;
assign a42032 = ~a42030 & a41960;
assign a42034 = a42032 & a41684;
assign a42036 = ~l2140 & l890;
assign a42038 = a40452 & a40430;
assign a42040 = a42038 & a38260;
assign a42042 = a41084 & ~a40778;
assign a42044 = ~a42042 & a42040;
assign a42046 = a42042 & i738;
assign a42048 = ~a42046 & ~a42044;
assign a42050 = a41982 & a40748;
assign a42052 = a42050 & ~a40784;
assign a42054 = ~a42052 & ~a42048;
assign a42056 = a42052 & i742;
assign a42058 = ~a42056 & ~a42054;
assign a42060 = ~a42058 & ~l890;
assign a42062 = ~a42060 & ~a42036;
assign a42064 = ~a42062 & ~l2124;
assign a42066 = a42064 & a41746;
assign a42068 = a42066 & a40642;
assign a42070 = ~a40992 & ~l2120;
assign a42072 = ~l2142 & l890;
assign a42074 = a41544 & a40430;
assign a42076 = a42074 & a38260;
assign a42078 = a41850 & ~a40778;
assign a42080 = ~a42078 & a42076;
assign a42082 = a42078 & i738;
assign a42084 = ~a42082 & ~a42080;
assign a42086 = a41866 & ~a40784;
assign a42088 = ~a42086 & ~a42084;
assign a42090 = a42086 & i742;
assign a42092 = ~a42090 & ~a42088;
assign a42094 = ~a42092 & ~l890;
assign a42096 = ~a42094 & ~a42072;
assign a42098 = ~a42096 & ~l2124;
assign a42100 = a42098 & a42070;
assign a42102 = a42100 & ~a40642;
assign a42104 = ~l2144 & l890;
assign a42106 = a41984 & a40784;
assign a42108 = ~a42106 & ~a41492;
assign a42110 = a42106 & i742;
assign a42112 = ~a42110 & ~a42108;
assign a42114 = ~a42112 & ~l890;
assign a42116 = ~a42114 & ~a42104;
assign a42118 = ~l2124 & ~l2120;
assign a42120 = a42118 & ~a42116;
assign a42122 = a42120 & ~a40992;
assign a42124 = a42122 & a40642;
assign a42126 = ~l2146 & l890;
assign a42128 = a42018 & a40784;
assign a42130 = ~a42128 & ~a41468;
assign a42132 = a42128 & i742;
assign a42134 = ~a42132 & ~a42130;
assign a42136 = ~a42134 & ~l890;
assign a42138 = ~a42136 & ~a42126;
assign a42140 = ~a42138 & a42118;
assign a42142 = a42140 & a40992;
assign a42144 = a42142 & ~a40642;
assign a42146 = ~l2148 & l890;
assign a42148 = a42050 & a40784;
assign a42150 = ~a42148 & ~a41478;
assign a42152 = a42148 & i742;
assign a42154 = ~a42152 & ~a42150;
assign a42156 = ~a42154 & ~l890;
assign a42158 = ~a42156 & ~a42146;
assign a42160 = ~a42158 & a41880;
assign a42162 = a40642 & ~l2124;
assign a42164 = a42162 & a42160;
assign a42166 = ~a42164 & ~a42144;
assign a42168 = a42166 & ~a42124;
assign a42170 = a42168 & ~a42102;
assign a42172 = a42170 & ~a42068;
assign a42174 = a42172 & ~a42034;
assign a42176 = a42174 & ~a42002;
assign a42178 = a42176 & ~a41966;
assign a42180 = a42178 & ~a41932;
assign a42182 = a42180 & ~a41886;
assign a42184 = ~a42182 & ~a41516;
assign a42186 = a42120 & a41684;
assign a42188 = a42142 & a40642;
assign a42190 = ~a42188 & ~a42186;
assign a42192 = a42100 & a40642;
assign a42194 = ~a42192 & a42190;
assign a42196 = a42064 & a41750;
assign a42198 = ~a42196 & a42194;
assign a42200 = a42032 & a40642;
assign a42202 = a42200 & a40992;
assign a42204 = ~a42202 & a42198;
assign a42206 = a41998 & a41684;
assign a42208 = ~a42206 & a42204;
assign a42210 = a41964 & a40642;
assign a42212 = ~a42210 & a42208;
assign a42214 = a41960 & a41748;
assign a42216 = a42214 & ~a41926;
assign a42218 = ~a42216 & a42212;
assign a42220 = a41884 & a40642;
assign a42222 = ~a42220 & a42218;
assign a42224 = a42160 & ~a40642;
assign a42226 = a42224 & l2124;
assign a42228 = ~a42226 & a42222;
assign a42230 = ~a42228 & a41516;
assign a42232 = ~a42230 & ~a42184;
assign a42234 = a42232 & i740;
assign a42236 = ~a42232 & ~i740;
assign a42238 = ~l2150 & l890;
assign a42240 = a41546 & i604;
assign a42242 = a42240 & ~a41852;
assign a42244 = a41852 & i734;
assign a42246 = ~a42244 & ~a42242;
assign a42248 = ~a42246 & ~a41868;
assign a42250 = a41868 & i748;
assign a42252 = ~a42250 & ~a42248;
assign a42254 = ~a42252 & ~l890;
assign a42256 = ~a42254 & ~a42238;
assign a42258 = ~a42256 & a41880;
assign a42260 = a42258 & l2124;
assign a42262 = a42260 & ~a40642;
assign a42264 = ~l2152 & l890;
assign a42266 = a41902 & i604;
assign a42268 = a42266 & ~a41896;
assign a42270 = a41896 & i734;
assign a42272 = ~a42270 & ~a42268;
assign a42274 = ~a42272 & ~a41916;
assign a42276 = a41916 & i748;
assign a42278 = ~a42276 & ~a42274;
assign a42280 = ~a42278 & ~l890;
assign a42282 = ~a42280 & ~a42264;
assign a42284 = ~a42282 & a41928;
assign a42286 = a42284 & a40642;
assign a42288 = ~l2154 & l890;
assign a42290 = a41936 & i604;
assign a42292 = a42290 & ~a41940;
assign a42294 = a41940 & i734;
assign a42296 = ~a42294 & ~a42292;
assign a42298 = ~a42296 & ~a41948;
assign a42300 = a41948 & i748;
assign a42302 = ~a42300 & ~a42298;
assign a42304 = ~a42302 & ~l890;
assign a42306 = ~a42304 & ~a42288;
assign a42308 = ~a42306 & a41962;
assign a42310 = a42308 & ~a40642;
assign a42312 = ~l2156 & l890;
assign a42314 = a41970 & i604;
assign a42316 = a42314 & ~a41974;
assign a42318 = a41974 & i734;
assign a42320 = ~a42318 & ~a42316;
assign a42322 = ~a42320 & ~a41986;
assign a42324 = a41986 & i748;
assign a42326 = ~a42324 & ~a42322;
assign a42328 = ~a42326 & ~l890;
assign a42330 = ~a42328 & ~a42312;
assign a42332 = ~a42330 & a41960;
assign a42334 = a42332 & ~a40992;
assign a42336 = a42334 & a40642;
assign a42338 = ~l2158 & l890;
assign a42340 = a42006 & i604;
assign a42342 = a42340 & ~a42010;
assign a42344 = a42010 & i734;
assign a42346 = ~a42344 & ~a42342;
assign a42348 = ~a42346 & ~a42020;
assign a42350 = a42020 & i748;
assign a42352 = ~a42350 & ~a42348;
assign a42354 = ~a42352 & ~l890;
assign a42356 = ~a42354 & ~a42338;
assign a42358 = ~a42356 & a41960;
assign a42360 = a42358 & a41684;
assign a42362 = ~l2160 & l890;
assign a42364 = a42038 & i604;
assign a42366 = a42364 & ~a42042;
assign a42368 = a42042 & i734;
assign a42370 = ~a42368 & ~a42366;
assign a42372 = ~a42370 & ~a42052;
assign a42374 = a42052 & i748;
assign a42376 = ~a42374 & ~a42372;
assign a42378 = ~a42376 & ~l890;
assign a42380 = ~a42378 & ~a42362;
assign a42382 = ~a42380 & ~l2124;
assign a42384 = a42382 & a41746;
assign a42386 = a42384 & a40642;
assign a42388 = ~l2162 & l890;
assign a42390 = a42074 & i604;
assign a42392 = a42390 & ~a42078;
assign a42394 = a42078 & i734;
assign a42396 = ~a42394 & ~a42392;
assign a42398 = ~a42396 & ~a42086;
assign a42400 = a42086 & i748;
assign a42402 = ~a42400 & ~a42398;
assign a42404 = ~a42402 & ~l890;
assign a42406 = ~a42404 & ~a42388;
assign a42408 = ~a42406 & ~l2124;
assign a42410 = a42408 & a42070;
assign a42412 = a42410 & ~a40642;
assign a42414 = ~l2164 & l890;
assign a42416 = ~a42106 & ~a41442;
assign a42418 = a42106 & i748;
assign a42420 = ~a42418 & ~a42416;
assign a42422 = ~a42420 & ~l890;
assign a42424 = ~a42422 & ~a42414;
assign a42426 = ~a42424 & a42118;
assign a42428 = a42426 & ~a40992;
assign a42430 = a42428 & a40642;
assign a42432 = ~l2166 & l890;
assign a42434 = ~a42128 & ~a41420;
assign a42436 = a42128 & i748;
assign a42438 = ~a42436 & ~a42434;
assign a42440 = ~a42438 & ~l890;
assign a42442 = ~a42440 & ~a42432;
assign a42444 = ~a42442 & a42118;
assign a42446 = a42444 & a40992;
assign a42448 = a42446 & ~a40642;
assign a42450 = ~l2168 & l890;
assign a42452 = ~a42148 & ~a41428;
assign a42454 = a42148 & i748;
assign a42456 = ~a42454 & ~a42452;
assign a42458 = ~a42456 & ~l890;
assign a42460 = ~a42458 & ~a42450;
assign a42462 = ~a42460 & a41880;
assign a42464 = a42462 & a42162;
assign a42466 = ~a42464 & ~a42448;
assign a42468 = a42466 & ~a42430;
assign a42470 = a42468 & ~a42412;
assign a42472 = a42470 & ~a42386;
assign a42474 = a42472 & ~a42360;
assign a42476 = a42474 & ~a42336;
assign a42478 = a42476 & ~a42310;
assign a42480 = a42478 & ~a42286;
assign a42482 = a42480 & ~a42262;
assign a42484 = ~a42482 & ~a41516;
assign a42486 = a42426 & a41684;
assign a42488 = a42446 & a40642;
assign a42490 = ~a42488 & ~a42486;
assign a42492 = a42410 & a40642;
assign a42494 = ~a42492 & a42490;
assign a42496 = a42382 & a41750;
assign a42498 = ~a42496 & a42494;
assign a42500 = a42358 & a40642;
assign a42502 = a42500 & a40992;
assign a42504 = ~a42502 & a42498;
assign a42506 = a42332 & a41684;
assign a42508 = ~a42506 & a42504;
assign a42510 = a42308 & a40642;
assign a42512 = ~a42510 & a42508;
assign a42514 = ~a42282 & a42214;
assign a42516 = ~a42514 & a42512;
assign a42518 = a42260 & a40642;
assign a42520 = ~a42518 & a42516;
assign a42522 = a42462 & ~a40642;
assign a42524 = a42522 & l2124;
assign a42526 = ~a42524 & a42520;
assign a42528 = ~a42526 & a41516;
assign a42530 = ~a42528 & ~a42484;
assign a42532 = a42530 & i746;
assign a42534 = ~a42530 & ~i746;
assign a42536 = ~l2170 & l890;
assign a42538 = a41546 & i602;
assign a42540 = a42538 & ~a41852;
assign a42542 = a41852 & i730;
assign a42544 = ~a42542 & ~a42540;
assign a42546 = ~a42544 & ~a41868;
assign a42548 = a41868 & i754;
assign a42550 = ~a42548 & ~a42546;
assign a42552 = ~a42550 & ~l890;
assign a42554 = ~a42552 & ~a42536;
assign a42556 = ~a42554 & a41880;
assign a42558 = a42556 & l2124;
assign a42560 = a42558 & ~a40642;
assign a42562 = ~l2172 & l890;
assign a42564 = a41902 & i602;
assign a42566 = a42564 & ~a41896;
assign a42568 = a41896 & i730;
assign a42570 = ~a42568 & ~a42566;
assign a42572 = ~a42570 & ~a41916;
assign a42574 = a41916 & i754;
assign a42576 = ~a42574 & ~a42572;
assign a42578 = ~a42576 & ~l890;
assign a42580 = ~a42578 & ~a42562;
assign a42582 = ~a42580 & a41928;
assign a42584 = a42582 & a40642;
assign a42586 = ~l2174 & l890;
assign a42588 = a41936 & i602;
assign a42590 = a42588 & ~a41940;
assign a42592 = a41940 & i730;
assign a42594 = ~a42592 & ~a42590;
assign a42596 = ~a42594 & ~a41948;
assign a42598 = a41948 & i754;
assign a42600 = ~a42598 & ~a42596;
assign a42602 = ~a42600 & ~l890;
assign a42604 = ~a42602 & ~a42586;
assign a42606 = ~a42604 & a41962;
assign a42608 = a42606 & ~a40642;
assign a42610 = ~l2176 & l890;
assign a42612 = a41970 & i602;
assign a42614 = a42612 & ~a41974;
assign a42616 = a41974 & i730;
assign a42618 = ~a42616 & ~a42614;
assign a42620 = ~a42618 & ~a41986;
assign a42622 = a41986 & i754;
assign a42624 = ~a42622 & ~a42620;
assign a42626 = ~a42624 & ~l890;
assign a42628 = ~a42626 & ~a42610;
assign a42630 = ~a42628 & a41960;
assign a42632 = a42630 & ~a40992;
assign a42634 = a42632 & a40642;
assign a42636 = ~l2178 & l890;
assign a42638 = a42006 & i602;
assign a42640 = a42638 & ~a42010;
assign a42642 = a42010 & i730;
assign a42644 = ~a42642 & ~a42640;
assign a42646 = ~a42644 & ~a42020;
assign a42648 = a42020 & i754;
assign a42650 = ~a42648 & ~a42646;
assign a42652 = ~a42650 & ~l890;
assign a42654 = ~a42652 & ~a42636;
assign a42656 = ~a42654 & a41960;
assign a42658 = a42656 & a41684;
assign a42660 = ~l2180 & l890;
assign a42662 = a42038 & i602;
assign a42664 = a42662 & ~a42042;
assign a42666 = a42042 & i730;
assign a42668 = ~a42666 & ~a42664;
assign a42670 = ~a42668 & ~a42052;
assign a42672 = a42052 & i754;
assign a42674 = ~a42672 & ~a42670;
assign a42676 = ~a42674 & ~l890;
assign a42678 = ~a42676 & ~a42660;
assign a42680 = ~a42678 & ~l2124;
assign a42682 = a42680 & a41746;
assign a42684 = a42682 & a40642;
assign a42686 = ~l2182 & l890;
assign a42688 = a42074 & i602;
assign a42690 = a42688 & ~a42078;
assign a42692 = a42078 & i730;
assign a42694 = ~a42692 & ~a42690;
assign a42696 = ~a42694 & ~a42086;
assign a42698 = a42086 & i754;
assign a42700 = ~a42698 & ~a42696;
assign a42702 = ~a42700 & ~l890;
assign a42704 = ~a42702 & ~a42686;
assign a42706 = ~a42704 & ~l2124;
assign a42708 = a42706 & a42070;
assign a42710 = a42708 & ~a40642;
assign a42712 = ~l2184 & l890;
assign a42714 = ~a42106 & ~a41396;
assign a42716 = a42106 & i754;
assign a42718 = ~a42716 & ~a42714;
assign a42720 = ~a42718 & ~l890;
assign a42722 = ~a42720 & ~a42712;
assign a42724 = ~a42722 & a42118;
assign a42726 = a42724 & ~a40992;
assign a42728 = a42726 & a40642;
assign a42730 = ~l2186 & l890;
assign a42732 = ~a42128 & ~a41374;
assign a42734 = a42128 & i754;
assign a42736 = ~a42734 & ~a42732;
assign a42738 = ~a42736 & ~l890;
assign a42740 = ~a42738 & ~a42730;
assign a42742 = ~a42740 & a42118;
assign a42744 = a42742 & a40992;
assign a42746 = a42744 & ~a40642;
assign a42748 = ~l2188 & l890;
assign a42750 = ~a42148 & ~a41382;
assign a42752 = a42148 & i754;
assign a42754 = ~a42752 & ~a42750;
assign a42756 = ~a42754 & ~l890;
assign a42758 = ~a42756 & ~a42748;
assign a42760 = ~a42758 & a41880;
assign a42762 = a42760 & a42162;
assign a42764 = ~a42762 & ~a42746;
assign a42766 = a42764 & ~a42728;
assign a42768 = a42766 & ~a42710;
assign a42770 = a42768 & ~a42684;
assign a42772 = a42770 & ~a42658;
assign a42774 = a42772 & ~a42634;
assign a42776 = a42774 & ~a42608;
assign a42778 = a42776 & ~a42584;
assign a42780 = a42778 & ~a42560;
assign a42782 = ~a42780 & ~a41516;
assign a42784 = a42724 & a41684;
assign a42786 = a42744 & a40642;
assign a42788 = ~a42786 & ~a42784;
assign a42790 = a42708 & a40642;
assign a42792 = ~a42790 & a42788;
assign a42794 = a42680 & a41750;
assign a42796 = ~a42794 & a42792;
assign a42798 = a42656 & a40642;
assign a42800 = a42798 & a40992;
assign a42802 = ~a42800 & a42796;
assign a42804 = a42630 & a41684;
assign a42806 = ~a42804 & a42802;
assign a42808 = a42606 & a40642;
assign a42810 = ~a42808 & a42806;
assign a42812 = ~a42580 & a42214;
assign a42814 = ~a42812 & a42810;
assign a42816 = a42558 & a40642;
assign a42818 = ~a42816 & a42814;
assign a42820 = a42760 & ~a40642;
assign a42822 = a42820 & l2124;
assign a42824 = ~a42822 & a42818;
assign a42826 = ~a42824 & a41516;
assign a42828 = ~a42826 & ~a42782;
assign a42830 = a42828 & i752;
assign a42832 = ~a42828 & ~i752;
assign a42834 = ~l2190 & l890;
assign a42836 = a41546 & i598;
assign a42838 = a42836 & ~a41852;
assign a42840 = a41852 & i726;
assign a42842 = ~a42840 & ~a42838;
assign a42844 = ~a42842 & ~a41868;
assign a42846 = a41868 & i760;
assign a42848 = ~a42846 & ~a42844;
assign a42850 = ~a42848 & ~l890;
assign a42852 = ~a42850 & ~a42834;
assign a42854 = ~a42852 & a41880;
assign a42856 = a42854 & l2124;
assign a42858 = a42856 & ~a40642;
assign a42860 = ~l2192 & l890;
assign a42862 = a41902 & i598;
assign a42864 = a42862 & ~a41896;
assign a42866 = a41896 & i726;
assign a42868 = ~a42866 & ~a42864;
assign a42870 = ~a42868 & ~a41916;
assign a42872 = a41916 & i760;
assign a42874 = ~a42872 & ~a42870;
assign a42876 = ~a42874 & ~l890;
assign a42878 = ~a42876 & ~a42860;
assign a42880 = ~a42878 & a41928;
assign a42882 = a42880 & a40642;
assign a42884 = ~l2194 & l890;
assign a42886 = a41936 & i598;
assign a42888 = a42886 & ~a41940;
assign a42890 = a41940 & i726;
assign a42892 = ~a42890 & ~a42888;
assign a42894 = ~a42892 & ~a41948;
assign a42896 = a41948 & i760;
assign a42898 = ~a42896 & ~a42894;
assign a42900 = ~a42898 & ~l890;
assign a42902 = ~a42900 & ~a42884;
assign a42904 = ~a42902 & a41962;
assign a42906 = a42904 & ~a40642;
assign a42908 = ~l2196 & l890;
assign a42910 = a41970 & i598;
assign a42912 = a42910 & ~a41974;
assign a42914 = a41974 & i726;
assign a42916 = ~a42914 & ~a42912;
assign a42918 = ~a42916 & ~a41986;
assign a42920 = a41986 & i760;
assign a42922 = ~a42920 & ~a42918;
assign a42924 = ~a42922 & ~l890;
assign a42926 = ~a42924 & ~a42908;
assign a42928 = ~a42926 & a41960;
assign a42930 = a42928 & ~a40992;
assign a42932 = a42930 & a40642;
assign a42934 = ~l2198 & l890;
assign a42936 = a42006 & i598;
assign a42938 = a42936 & ~a42010;
assign a42940 = a42010 & i726;
assign a42942 = ~a42940 & ~a42938;
assign a42944 = ~a42942 & ~a42020;
assign a42946 = a42020 & i760;
assign a42948 = ~a42946 & ~a42944;
assign a42950 = ~a42948 & ~l890;
assign a42952 = ~a42950 & ~a42934;
assign a42954 = ~a42952 & a41960;
assign a42956 = a42954 & a41684;
assign a42958 = ~l2200 & l890;
assign a42960 = a42038 & i598;
assign a42962 = a42960 & ~a42042;
assign a42964 = a42042 & i726;
assign a42966 = ~a42964 & ~a42962;
assign a42968 = ~a42966 & ~a42052;
assign a42970 = a42052 & i760;
assign a42972 = ~a42970 & ~a42968;
assign a42974 = ~a42972 & ~l890;
assign a42976 = ~a42974 & ~a42958;
assign a42978 = ~a42976 & ~l2124;
assign a42980 = a42978 & a41746;
assign a42982 = a42980 & a40642;
assign a42984 = ~l2202 & l890;
assign a42986 = a42074 & i598;
assign a42988 = a42986 & ~a42078;
assign a42990 = a42078 & i726;
assign a42992 = ~a42990 & ~a42988;
assign a42994 = ~a42992 & ~a42086;
assign a42996 = a42086 & i760;
assign a42998 = ~a42996 & ~a42994;
assign a43000 = ~a42998 & ~l890;
assign a43002 = ~a43000 & ~a42984;
assign a43004 = ~a43002 & ~l2124;
assign a43006 = a43004 & a42070;
assign a43008 = a43006 & ~a40642;
assign a43010 = ~l2204 & l890;
assign a43012 = ~a42106 & ~a41350;
assign a43014 = a42106 & i760;
assign a43016 = ~a43014 & ~a43012;
assign a43018 = ~a43016 & ~l890;
assign a43020 = ~a43018 & ~a43010;
assign a43022 = ~a43020 & a42118;
assign a43024 = a43022 & ~a40992;
assign a43026 = a43024 & a40642;
assign a43028 = ~l2206 & l890;
assign a43030 = ~a42128 & ~a41328;
assign a43032 = a42128 & i760;
assign a43034 = ~a43032 & ~a43030;
assign a43036 = ~a43034 & ~l890;
assign a43038 = ~a43036 & ~a43028;
assign a43040 = ~a43038 & a42118;
assign a43042 = a43040 & a40992;
assign a43044 = a43042 & ~a40642;
assign a43046 = ~l2208 & l890;
assign a43048 = ~a42148 & ~a41336;
assign a43050 = a42148 & i760;
assign a43052 = ~a43050 & ~a43048;
assign a43054 = ~a43052 & ~l890;
assign a43056 = ~a43054 & ~a43046;
assign a43058 = ~a43056 & a41880;
assign a43060 = a43058 & a42162;
assign a43062 = ~a43060 & ~a43044;
assign a43064 = a43062 & ~a43026;
assign a43066 = a43064 & ~a43008;
assign a43068 = a43066 & ~a42982;
assign a43070 = a43068 & ~a42956;
assign a43072 = a43070 & ~a42932;
assign a43074 = a43072 & ~a42906;
assign a43076 = a43074 & ~a42882;
assign a43078 = a43076 & ~a42858;
assign a43080 = ~a43078 & ~a41516;
assign a43082 = a43022 & a41684;
assign a43084 = a43042 & a40642;
assign a43086 = ~a43084 & ~a43082;
assign a43088 = a43006 & a40642;
assign a43090 = ~a43088 & a43086;
assign a43092 = a42978 & a41750;
assign a43094 = ~a43092 & a43090;
assign a43096 = a42954 & a40642;
assign a43098 = a43096 & a40992;
assign a43100 = ~a43098 & a43094;
assign a43102 = a42928 & a41684;
assign a43104 = ~a43102 & a43100;
assign a43106 = a42904 & a40642;
assign a43108 = ~a43106 & a43104;
assign a43110 = ~a42878 & a42214;
assign a43112 = ~a43110 & a43108;
assign a43114 = a42856 & a40642;
assign a43116 = ~a43114 & a43112;
assign a43118 = a43058 & ~a40642;
assign a43120 = a43118 & l2124;
assign a43122 = ~a43120 & a43116;
assign a43124 = ~a43122 & a41516;
assign a43126 = ~a43124 & ~a43080;
assign a43128 = a43126 & i758;
assign a43130 = ~a43126 & ~i758;
assign a43132 = ~l2210 & l890;
assign a43134 = a41546 & i592;
assign a43136 = a43134 & ~a41852;
assign a43138 = a41852 & i722;
assign a43140 = ~a43138 & ~a43136;
assign a43142 = ~a43140 & ~a41868;
assign a43144 = a41868 & i766;
assign a43146 = ~a43144 & ~a43142;
assign a43148 = ~a43146 & ~l890;
assign a43150 = ~a43148 & ~a43132;
assign a43152 = ~a43150 & a41880;
assign a43154 = a43152 & l2124;
assign a43156 = a43154 & ~a40642;
assign a43158 = ~l2212 & l890;
assign a43160 = a41902 & i592;
assign a43162 = a43160 & ~a41896;
assign a43164 = a41896 & i722;
assign a43166 = ~a43164 & ~a43162;
assign a43168 = ~a43166 & ~a41916;
assign a43170 = a41916 & i766;
assign a43172 = ~a43170 & ~a43168;
assign a43174 = ~a43172 & ~l890;
assign a43176 = ~a43174 & ~a43158;
assign a43178 = ~a43176 & a41928;
assign a43180 = a43178 & a40642;
assign a43182 = ~l2214 & l890;
assign a43184 = a41936 & i592;
assign a43186 = a43184 & ~a41940;
assign a43188 = a41940 & i722;
assign a43190 = ~a43188 & ~a43186;
assign a43192 = ~a43190 & ~a41948;
assign a43194 = a41948 & i766;
assign a43196 = ~a43194 & ~a43192;
assign a43198 = ~a43196 & ~l890;
assign a43200 = ~a43198 & ~a43182;
assign a43202 = ~a43200 & a41962;
assign a43204 = a43202 & ~a40642;
assign a43206 = ~l2216 & l890;
assign a43208 = a41970 & i592;
assign a43210 = a43208 & ~a41974;
assign a43212 = a41974 & i722;
assign a43214 = ~a43212 & ~a43210;
assign a43216 = ~a43214 & ~a41986;
assign a43218 = a41986 & i766;
assign a43220 = ~a43218 & ~a43216;
assign a43222 = ~a43220 & ~l890;
assign a43224 = ~a43222 & ~a43206;
assign a43226 = ~a43224 & a41960;
assign a43228 = a43226 & ~a40992;
assign a43230 = a43228 & a40642;
assign a43232 = ~l2218 & l890;
assign a43234 = a42006 & i592;
assign a43236 = a43234 & ~a42010;
assign a43238 = a42010 & i722;
assign a43240 = ~a43238 & ~a43236;
assign a43242 = ~a43240 & ~a42020;
assign a43244 = a42020 & i766;
assign a43246 = ~a43244 & ~a43242;
assign a43248 = ~a43246 & ~l890;
assign a43250 = ~a43248 & ~a43232;
assign a43252 = ~a43250 & a41960;
assign a43254 = a43252 & a41684;
assign a43256 = ~l2220 & l890;
assign a43258 = a42038 & i592;
assign a43260 = a43258 & ~a42042;
assign a43262 = a42042 & i722;
assign a43264 = ~a43262 & ~a43260;
assign a43266 = ~a43264 & ~a42052;
assign a43268 = a42052 & i766;
assign a43270 = ~a43268 & ~a43266;
assign a43272 = ~a43270 & ~l890;
assign a43274 = ~a43272 & ~a43256;
assign a43276 = ~a43274 & ~l2124;
assign a43278 = a43276 & a41746;
assign a43280 = a43278 & a40642;
assign a43282 = ~l2222 & l890;
assign a43284 = a42074 & i592;
assign a43286 = a43284 & ~a42078;
assign a43288 = a42078 & i722;
assign a43290 = ~a43288 & ~a43286;
assign a43292 = ~a43290 & ~a42086;
assign a43294 = a42086 & i766;
assign a43296 = ~a43294 & ~a43292;
assign a43298 = ~a43296 & ~l890;
assign a43300 = ~a43298 & ~a43282;
assign a43302 = ~a43300 & ~l2124;
assign a43304 = a43302 & a42070;
assign a43306 = a43304 & ~a40642;
assign a43308 = ~l2224 & l890;
assign a43310 = ~a42106 & ~a41304;
assign a43312 = a42106 & i766;
assign a43314 = ~a43312 & ~a43310;
assign a43316 = ~a43314 & ~l890;
assign a43318 = ~a43316 & ~a43308;
assign a43320 = ~a43318 & a42118;
assign a43322 = a43320 & ~a40992;
assign a43324 = a43322 & a40642;
assign a43326 = ~l2226 & l890;
assign a43328 = ~a42128 & ~a41282;
assign a43330 = a42128 & i766;
assign a43332 = ~a43330 & ~a43328;
assign a43334 = ~a43332 & ~l890;
assign a43336 = ~a43334 & ~a43326;
assign a43338 = ~a43336 & a42118;
assign a43340 = a43338 & a40992;
assign a43342 = a43340 & ~a40642;
assign a43344 = ~l2228 & l890;
assign a43346 = ~a42148 & ~a41290;
assign a43348 = a42148 & i766;
assign a43350 = ~a43348 & ~a43346;
assign a43352 = ~a43350 & ~l890;
assign a43354 = ~a43352 & ~a43344;
assign a43356 = ~a43354 & a41880;
assign a43358 = a43356 & a42162;
assign a43360 = ~a43358 & ~a43342;
assign a43362 = a43360 & ~a43324;
assign a43364 = a43362 & ~a43306;
assign a43366 = a43364 & ~a43280;
assign a43368 = a43366 & ~a43254;
assign a43370 = a43368 & ~a43230;
assign a43372 = a43370 & ~a43204;
assign a43374 = a43372 & ~a43180;
assign a43376 = a43374 & ~a43156;
assign a43378 = ~a43376 & ~a41516;
assign a43380 = a43320 & a41684;
assign a43382 = a43340 & a40642;
assign a43384 = ~a43382 & ~a43380;
assign a43386 = a43304 & a40642;
assign a43388 = ~a43386 & a43384;
assign a43390 = a43276 & a41750;
assign a43392 = ~a43390 & a43388;
assign a43394 = a43252 & a40642;
assign a43396 = a43394 & a40992;
assign a43398 = ~a43396 & a43392;
assign a43400 = a43226 & a41684;
assign a43402 = ~a43400 & a43398;
assign a43404 = a43202 & a40642;
assign a43406 = ~a43404 & a43402;
assign a43408 = ~a43176 & a42214;
assign a43410 = ~a43408 & a43406;
assign a43412 = a43154 & a40642;
assign a43414 = ~a43412 & a43410;
assign a43416 = a43356 & ~a40642;
assign a43418 = a43416 & l2124;
assign a43420 = ~a43418 & a43414;
assign a43422 = ~a43420 & a41516;
assign a43424 = ~a43422 & ~a43378;
assign a43426 = a43424 & i764;
assign a43428 = ~a43424 & ~i764;
assign a43430 = ~l2230 & l890;
assign a43432 = ~a41852 & a41564;
assign a43434 = a41852 & i718;
assign a43436 = ~a43434 & ~a43432;
assign a43438 = ~a43436 & ~a41868;
assign a43440 = a41868 & i772;
assign a43442 = ~a43440 & ~a43438;
assign a43444 = ~a43442 & ~l890;
assign a43446 = ~a43444 & ~a43430;
assign a43448 = ~a43446 & a41880;
assign a43450 = a43448 & l2124;
assign a43452 = a43450 & ~a40642;
assign a43454 = ~l2232 & l890;
assign a43456 = a41902 & i634;
assign a43458 = a43456 & ~a41896;
assign a43460 = a41896 & i718;
assign a43462 = ~a43460 & ~a43458;
assign a43464 = ~a43462 & ~a41916;
assign a43466 = a41916 & i772;
assign a43468 = ~a43466 & ~a43464;
assign a43470 = ~a43468 & ~l890;
assign a43472 = ~a43470 & ~a43454;
assign a43474 = ~a43472 & a41928;
assign a43476 = a43474 & a40642;
assign a43478 = ~l2234 & l890;
assign a43480 = a41936 & i634;
assign a43482 = a43480 & ~a41940;
assign a43484 = a41940 & i718;
assign a43486 = ~a43484 & ~a43482;
assign a43488 = ~a43486 & ~a41948;
assign a43490 = a41948 & i772;
assign a43492 = ~a43490 & ~a43488;
assign a43494 = ~a43492 & ~l890;
assign a43496 = ~a43494 & ~a43478;
assign a43498 = ~a43496 & a41962;
assign a43500 = a43498 & ~a40642;
assign a43502 = ~l2236 & l890;
assign a43504 = a41970 & i634;
assign a43506 = a43504 & ~a41974;
assign a43508 = a41974 & i718;
assign a43510 = ~a43508 & ~a43506;
assign a43512 = ~a43510 & ~a41986;
assign a43514 = a41986 & i772;
assign a43516 = ~a43514 & ~a43512;
assign a43518 = ~a43516 & ~l890;
assign a43520 = ~a43518 & ~a43502;
assign a43522 = ~a43520 & a41960;
assign a43524 = a43522 & ~a40992;
assign a43526 = a43524 & a40642;
assign a43528 = ~l2238 & l890;
assign a43530 = a42006 & i634;
assign a43532 = a43530 & ~a42010;
assign a43534 = a42010 & i718;
assign a43536 = ~a43534 & ~a43532;
assign a43538 = ~a43536 & ~a42020;
assign a43540 = a42020 & i772;
assign a43542 = ~a43540 & ~a43538;
assign a43544 = ~a43542 & ~l890;
assign a43546 = ~a43544 & ~a43528;
assign a43548 = ~a43546 & a41960;
assign a43550 = a43548 & a41684;
assign a43552 = ~l2240 & l890;
assign a43554 = a42038 & i634;
assign a43556 = a43554 & ~a42042;
assign a43558 = a42042 & i718;
assign a43560 = ~a43558 & ~a43556;
assign a43562 = ~a43560 & ~a42052;
assign a43564 = a42052 & i772;
assign a43566 = ~a43564 & ~a43562;
assign a43568 = ~a43566 & ~l890;
assign a43570 = ~a43568 & ~a43552;
assign a43572 = ~a43570 & ~l2124;
assign a43574 = a43572 & a41746;
assign a43576 = a43574 & a40642;
assign a43578 = ~l2242 & l890;
assign a43580 = a42074 & i634;
assign a43582 = a43580 & ~a42078;
assign a43584 = a42078 & i718;
assign a43586 = ~a43584 & ~a43582;
assign a43588 = ~a43586 & ~a42086;
assign a43590 = a42086 & i772;
assign a43592 = ~a43590 & ~a43588;
assign a43594 = ~a43592 & ~l890;
assign a43596 = ~a43594 & ~a43578;
assign a43598 = ~a43596 & ~l2124;
assign a43600 = a43598 & a42070;
assign a43602 = a43600 & ~a40642;
assign a43604 = ~l2244 & l890;
assign a43606 = ~a42106 & ~a41258;
assign a43608 = a42106 & i772;
assign a43610 = ~a43608 & ~a43606;
assign a43612 = ~a43610 & ~l890;
assign a43614 = ~a43612 & ~a43604;
assign a43616 = ~a43614 & a42118;
assign a43618 = a43616 & ~a40992;
assign a43620 = a43618 & a40642;
assign a43622 = ~l2246 & l890;
assign a43624 = ~a42128 & ~a41236;
assign a43626 = a42128 & i772;
assign a43628 = ~a43626 & ~a43624;
assign a43630 = ~a43628 & ~l890;
assign a43632 = ~a43630 & ~a43622;
assign a43634 = ~a43632 & a42118;
assign a43636 = a43634 & a40992;
assign a43638 = a43636 & ~a40642;
assign a43640 = ~l2248 & l890;
assign a43642 = ~a42148 & ~a41244;
assign a43644 = a42148 & i772;
assign a43646 = ~a43644 & ~a43642;
assign a43648 = ~a43646 & ~l890;
assign a43650 = ~a43648 & ~a43640;
assign a43652 = ~a43650 & a41880;
assign a43654 = a43652 & a42162;
assign a43656 = ~a43654 & ~a43638;
assign a43658 = a43656 & ~a43620;
assign a43660 = a43658 & ~a43602;
assign a43662 = a43660 & ~a43576;
assign a43664 = a43662 & ~a43550;
assign a43666 = a43664 & ~a43526;
assign a43668 = a43666 & ~a43500;
assign a43670 = a43668 & ~a43476;
assign a43672 = a43670 & ~a43452;
assign a43674 = ~a43672 & ~a41516;
assign a43676 = a43616 & a41684;
assign a43678 = a43636 & a40642;
assign a43680 = ~a43678 & ~a43676;
assign a43682 = a43600 & a40642;
assign a43684 = ~a43682 & a43680;
assign a43686 = a43572 & a41750;
assign a43688 = ~a43686 & a43684;
assign a43690 = a43548 & a40642;
assign a43692 = a43690 & a40992;
assign a43694 = ~a43692 & a43688;
assign a43696 = a43522 & a41684;
assign a43698 = ~a43696 & a43694;
assign a43700 = a43498 & a40642;
assign a43702 = ~a43700 & a43698;
assign a43704 = ~a43472 & a42214;
assign a43706 = ~a43704 & a43702;
assign a43708 = a43450 & a40642;
assign a43710 = ~a43708 & a43706;
assign a43712 = a43652 & ~a40642;
assign a43714 = a43712 & l2124;
assign a43716 = ~a43714 & a43710;
assign a43718 = ~a43716 & a41516;
assign a43720 = ~a43718 & ~a43674;
assign a43722 = a43720 & i770;
assign a43724 = ~a43720 & ~i770;
assign a43726 = ~l2250 & l890;
assign a43728 = ~a40788 & i664;
assign a43730 = ~a43728 & ~i560;
assign a43732 = ~a42128 & ~a41068;
assign a43734 = ~a43732 & a43730;
assign a43736 = ~a43734 & ~l890;
assign a43738 = ~a43736 & ~a43726;
assign a43740 = a43738 & ~l2124;
assign a43742 = ~l2402 & l890;
assign a43744 = ~a40492 & i778;
assign a43746 = ~a43744 & ~i590;
assign a43748 = a40492 & ~i778;
assign a43750 = ~a43748 & ~a43746;
assign a43752 = ~a40510 & i780;
assign a43754 = ~a43752 & ~a43750;
assign a43756 = a40510 & ~i780;
assign a43758 = ~a43756 & ~a43754;
assign a43760 = ~a40528 & i782;
assign a43762 = ~a43760 & ~a43758;
assign a43764 = a40528 & ~i782;
assign a43766 = ~a43764 & ~a43762;
assign a43768 = ~a40546 & i784;
assign a43770 = ~a43768 & ~a43766;
assign a43772 = a40546 & ~i784;
assign a43774 = ~a43772 & ~a43770;
assign a43776 = a43774 & ~i786;
assign a43778 = ~a43776 & a40604;
assign a43780 = ~a43768 & i786;
assign a43782 = a40210 & i622;
assign a43784 = a40238 & ~i622;
assign a43786 = ~a43784 & ~a43782;
assign a43788 = a40328 & i622;
assign a43790 = a40356 & ~i622;
assign a43792 = ~a43790 & ~a43788;
assign a43794 = a43792 & a40404;
assign a43796 = a43794 & a40264;
assign a43798 = a43796 & a40166;
assign a43800 = a43798 & a40672;
assign a43802 = a43800 & a43786;
assign a43804 = a43802 & a39998;
assign a43806 = a43804 & a40692;
assign a43808 = a43806 & i788;
assign a43810 = ~a43808 & ~a43748;
assign a43812 = ~a43810 & ~a43744;
assign a43814 = ~a43812 & ~a43756;
assign a43816 = ~a43814 & ~a43752;
assign a43818 = ~a43816 & ~a43764;
assign a43820 = ~a43818 & ~a43760;
assign a43822 = ~a43820 & ~a43772;
assign a43824 = ~a43822 & a43780;
assign a43826 = ~a43824 & a43778;
assign a43828 = ~a43826 & ~i560;
assign a43830 = ~a41852 & ~a41548;
assign a43832 = ~a43830 & ~a40624;
assign a43834 = ~a43832 & ~a41868;
assign a43836 = ~a43834 & a43828;
assign a43838 = ~a43836 & ~l890;
assign a43840 = ~a43838 & ~a43742;
assign a43842 = a43840 & l2124;
assign a43844 = ~a43842 & ~a43740;
assign a43846 = ~a43844 & a41514;
assign a43848 = ~l2362 & l890;
assign a43850 = a40784 & ~a40716;
assign a43852 = a43850 & a40772;
assign a43854 = ~a43852 & a40788;
assign a43856 = ~a43854 & i664;
assign a43858 = ~a43856 & ~i560;
assign a43860 = ~a42148 & ~a41090;
assign a43862 = ~a43860 & a43858;
assign a43864 = ~a43862 & ~l890;
assign a43866 = ~a43864 & ~a43848;
assign a43868 = a43866 & ~l2124;
assign a43870 = ~l2398 & l890;
assign a43872 = ~a40772 & ~a40716;
assign a43874 = a43872 & i664;
assign a43876 = ~a43874 & ~i560;
assign a43878 = ~a40766 & ~a40664;
assign a43880 = a43878 & i582;
assign a43882 = ~a43880 & ~a40624;
assign a43884 = a41902 & ~a40578;
assign a43886 = a40436 & a40434;
assign a43888 = a43886 & i564;
assign a43890 = ~a43888 & a43884;
assign a43892 = ~a43890 & ~a41896;
assign a43894 = ~a43892 & a43882;
assign a43896 = ~a43894 & ~a41916;
assign a43898 = ~a43896 & a43876;
assign a43900 = ~a43898 & ~l890;
assign a43902 = ~a43900 & ~a43870;
assign a43904 = a43902 & l2124;
assign a43906 = ~a43904 & ~a43868;
assign a43908 = ~a43906 & ~a41514;
assign a43910 = ~a43908 & ~a43846;
assign a43912 = ~a43910 & ~l2120;
assign a43914 = ~l2388 & l890;
assign a43916 = ~a40784 & ~a40748;
assign a43918 = ~a43916 & a40772;
assign a43920 = ~a43918 & i664;
assign a43922 = ~a43920 & ~i560;
assign a43924 = ~a40778 & ~a40742;
assign a43926 = ~a43924 & a40766;
assign a43928 = ~a43926 & i582;
assign a43930 = ~a43928 & ~a40624;
assign a43932 = a42006 & ~a40578;
assign a43934 = a40432 & a40430;
assign a43936 = ~a43934 & ~a40436;
assign a43938 = ~a43936 & i564;
assign a43940 = ~a43938 & a43932;
assign a43942 = ~a43940 & ~a42010;
assign a43944 = ~a43942 & a43930;
assign a43946 = ~a43944 & ~a42020;
assign a43948 = ~a43946 & a43922;
assign a43950 = ~a43948 & ~l890;
assign a43952 = ~a43950 & ~a43914;
assign a43954 = a43952 & ~l2124;
assign a43956 = a43954 & a41514;
assign a43958 = ~l2382 & l890;
assign a43960 = ~a40784 & ~a40716;
assign a43962 = ~a43960 & a43918;
assign a43964 = ~a43962 & i664;
assign a43966 = ~a43964 & ~i560;
assign a43968 = ~a40778 & ~a40664;
assign a43970 = ~a43968 & a43926;
assign a43972 = ~a43970 & i582;
assign a43974 = ~a43972 & ~a40624;
assign a43976 = a42038 & ~a40578;
assign a43978 = a40434 & a40430;
assign a43980 = ~a43978 & a43936;
assign a43982 = ~a43980 & i564;
assign a43984 = ~a43982 & a43976;
assign a43986 = ~a43984 & ~a42042;
assign a43988 = ~a43986 & a43974;
assign a43990 = ~a43988 & ~a42052;
assign a43992 = ~a43990 & a43966;
assign a43994 = ~a43992 & ~l890;
assign a43996 = ~a43994 & ~a43958;
assign a43998 = a43996 & ~l2124;
assign a44000 = a43998 & ~a41514;
assign a44002 = ~a44000 & ~a43956;
assign a44004 = ~a44002 & l2120;
assign a44006 = ~a44004 & ~a43912;
assign a44008 = ~a44006 & a40992;
assign a44010 = ~l2378 & l890;
assign a44012 = a40784 & a40772;
assign a44014 = ~a44012 & i664;
assign a44016 = ~a44014 & ~i560;
assign a44018 = ~a41048 & i582;
assign a44020 = ~a44018 & ~a40624;
assign a44022 = a42074 & ~a40578;
assign a44024 = ~a40582 & i564;
assign a44026 = ~a44024 & a44022;
assign a44028 = ~a44026 & ~a42078;
assign a44030 = ~a44028 & a44020;
assign a44032 = ~a44030 & ~a42086;
assign a44034 = ~a44032 & a44016;
assign a44036 = ~a44034 & ~l890;
assign a44038 = ~a44036 & ~a44010;
assign a44040 = a44038 & ~l2124;
assign a44042 = a44040 & a41514;
assign a44044 = ~l2374 & l890;
assign a44046 = a40784 & ~a40748;
assign a44048 = a44046 & ~a40716;
assign a44050 = ~a44048 & a44012;
assign a44052 = ~a44050 & i664;
assign a44054 = ~a44052 & ~i560;
assign a44056 = ~a42106 & ~a41126;
assign a44058 = ~a44056 & a44054;
assign a44060 = ~a44058 & ~l890;
assign a44062 = ~a44060 & ~a44044;
assign a44064 = a44062 & ~l2124;
assign a44066 = a44064 & ~a41514;
assign a44068 = ~a44066 & ~a44042;
assign a44070 = ~a44068 & ~l2120;
assign a44072 = ~l2394 & l890;
assign a44074 = ~a40772 & i664;
assign a44076 = ~a44074 & ~i560;
assign a44078 = ~a40766 & i582;
assign a44080 = ~a44078 & ~a40624;
assign a44082 = a41936 & ~a40578;
assign a44084 = a40436 & i564;
assign a44086 = ~a44084 & a44082;
assign a44088 = ~a44086 & ~a41940;
assign a44090 = ~a44088 & a44080;
assign a44092 = ~a44090 & ~a41948;
assign a44094 = ~a44092 & a44076;
assign a44096 = ~a44094 & ~l890;
assign a44098 = ~a44096 & ~a44072;
assign a44100 = a44098 & ~l2124;
assign a44102 = a44100 & a41514;
assign a44104 = ~l2392 & l890;
assign a44106 = a43916 & ~a40716;
assign a44108 = ~a44106 & a40772;
assign a44110 = ~a44108 & i664;
assign a44112 = ~a44110 & ~i560;
assign a44114 = a43924 & ~a40664;
assign a44116 = ~a44114 & a40766;
assign a44118 = ~a44116 & i582;
assign a44120 = ~a44118 & ~a40624;
assign a44122 = a41970 & ~a40578;
assign a44124 = a43934 & a40434;
assign a44126 = ~a44124 & ~a40436;
assign a44128 = ~a44126 & i564;
assign a44130 = ~a44128 & a44122;
assign a44132 = ~a44130 & ~a41974;
assign a44134 = ~a44132 & a44120;
assign a44136 = ~a44134 & ~a41986;
assign a44138 = ~a44136 & a44112;
assign a44140 = ~a44138 & ~l890;
assign a44142 = ~a44140 & ~a44104;
assign a44144 = a44142 & ~l2124;
assign a44146 = a44144 & ~a41514;
assign a44148 = ~a44146 & ~a44102;
assign a44150 = ~a44148 & l2120;
assign a44152 = ~a44150 & ~a44070;
assign a44154 = ~a44152 & ~a40992;
assign a44156 = ~a44154 & ~a44008;
assign a44158 = ~a44156 & a40730;
assign a44160 = ~a44148 & a41024;
assign a44162 = a44144 & ~a41024;
assign a44164 = ~a44162 & ~a44160;
assign a44166 = ~a44164 & l2120;
assign a44168 = ~a44166 & ~a44070;
assign a44170 = ~a44168 & a41008;
assign a44172 = ~a44068 & a41024;
assign a44174 = a44064 & ~a41024;
assign a44176 = ~a44174 & ~a44172;
assign a44178 = ~a44176 & ~l2120;
assign a44180 = ~a44178 & ~a44150;
assign a44182 = ~a44180 & ~a41008;
assign a44184 = ~a44182 & ~a44170;
assign a44186 = ~a44184 & ~a40992;
assign a44188 = ~a44186 & ~a44008;
assign a44190 = ~a44188 & a40758;
assign a44192 = ~a44002 & a41024;
assign a44194 = a43998 & ~a41024;
assign a44196 = ~a44194 & ~a44192;
assign a44198 = ~a44196 & l2120;
assign a44200 = ~a44198 & ~a43912;
assign a44202 = ~a44200 & a41008;
assign a44204 = ~a43904 & ~a43740;
assign a44206 = ~a44204 & a41514;
assign a44208 = ~a44206 & ~a43908;
assign a44210 = ~a44208 & a41024;
assign a44212 = ~a43868 & ~a43842;
assign a44214 = ~a44212 & a41514;
assign a44216 = ~a44214 & ~a43908;
assign a44218 = ~a44216 & ~a41024;
assign a44220 = ~a44218 & ~a44210;
assign a44222 = ~a44220 & ~l2120;
assign a44224 = ~a44222 & ~a44004;
assign a44226 = ~a44224 & ~a41008;
assign a44228 = ~a44226 & ~a44202;
assign a44230 = ~a44228 & a40992;
assign a44232 = ~a44230 & ~a44154;
assign a44234 = ~a44232 & ~a40758;
assign a44236 = ~a44234 & ~a44190;
assign a44238 = ~a44236 & ~a40730;
assign a44240 = ~a44238 & ~a44158;
assign a44242 = ~a44240 & a40642;
assign a44244 = a43866 & l2124;
assign a44246 = ~a44244 & ~a44064;
assign a44248 = ~a44246 & a41514;
assign a44250 = ~a43844 & ~a41514;
assign a44252 = ~a44250 & ~a44248;
assign a44254 = ~a44252 & ~l2120;
assign a44256 = a44144 & a41514;
assign a44258 = a43954 & ~a41514;
assign a44260 = ~a44258 & ~a44256;
assign a44262 = ~a44260 & l2120;
assign a44264 = ~a44262 & ~a44254;
assign a44266 = ~a44264 & a40992;
assign a44268 = a43998 & a41514;
assign a44270 = a44040 & ~a41514;
assign a44272 = ~a44270 & ~a44268;
assign a44274 = ~a44272 & ~l2120;
assign a44276 = a43902 & ~l2124;
assign a44278 = a44276 & a41514;
assign a44280 = a44100 & ~a41514;
assign a44282 = ~a44280 & ~a44278;
assign a44284 = ~a44282 & a41024;
assign a44286 = a44100 & ~a41024;
assign a44288 = ~a44286 & ~a44284;
assign a44290 = ~a44288 & l2120;
assign a44292 = ~a44290 & ~a44274;
assign a44294 = ~a44292 & a41008;
assign a44296 = ~a44272 & a41024;
assign a44298 = a44040 & ~a41024;
assign a44300 = ~a44298 & ~a44296;
assign a44302 = ~a44300 & ~l2120;
assign a44304 = ~a44282 & l2120;
assign a44306 = ~a44304 & ~a44302;
assign a44308 = ~a44306 & ~a41008;
assign a44310 = ~a44308 & ~a44294;
assign a44312 = ~a44310 & ~a40992;
assign a44314 = ~a44312 & ~a44266;
assign a44316 = ~a44314 & a40758;
assign a44318 = ~a44260 & a41024;
assign a44320 = a43954 & ~a41024;
assign a44322 = ~a44320 & ~a44318;
assign a44324 = ~a44322 & l2120;
assign a44326 = ~a44324 & ~a44254;
assign a44328 = ~a44326 & a41008;
assign a44330 = ~a44064 & ~a43842;
assign a44332 = ~a44330 & a41514;
assign a44334 = ~a44332 & ~a44250;
assign a44336 = ~a44334 & a41024;
assign a44338 = ~a44244 & ~a43740;
assign a44340 = ~a44338 & a41514;
assign a44342 = ~a44340 & ~a44250;
assign a44344 = ~a44342 & ~a41024;
assign a44346 = ~a44344 & ~a44336;
assign a44348 = ~a44346 & ~l2120;
assign a44350 = ~a44348 & ~a44262;
assign a44352 = ~a44350 & ~a41008;
assign a44354 = ~a44352 & ~a44328;
assign a44356 = ~a44354 & a40992;
assign a44358 = ~a44304 & ~a44274;
assign a44360 = ~a44358 & ~a40992;
assign a44362 = ~a44360 & ~a44356;
assign a44364 = ~a44362 & ~a40758;
assign a44366 = ~a44364 & ~a44316;
assign a44368 = ~a44366 & a40730;
assign a44370 = ~a44360 & ~a44266;
assign a44372 = ~a44370 & ~a40730;
assign a44374 = ~a44372 & ~a44368;
assign a44376 = ~a44374 & ~a40642;
assign a44378 = ~a44376 & ~a44242;
assign a44380 = a44378 & ~i654;
assign a44382 = ~a44380 & ~i654;
assign a44384 = a44382 & i776;
assign a44386 = a44384 & ~a43724;
assign a44388 = a44386 & ~a43722;
assign a44390 = a44388 & ~a43428;
assign a44392 = a44390 & ~a43426;
assign a44394 = a44392 & ~a43130;
assign a44396 = a44394 & ~a43128;
assign a44398 = a44396 & ~a42832;
assign a44400 = a44398 & ~a42830;
assign a44402 = a44400 & ~a42534;
assign a44404 = a44402 & ~a42532;
assign a44406 = a44404 & ~a42236;
assign a44410 = ~l2130 & l890;
assign a44412 = ~a40720 & ~l890;
assign a44414 = ~a44412 & ~a44410;
assign a44416 = a44414 & ~a41024;
assign a44418 = a44416 & ~a40730;
assign a44420 = a44418 & ~a40758;
assign a44422 = a44420 & ~a41008;
assign a44424 = ~a44422 & ~a41878;
assign a44426 = a44422 & i744;
assign a44430 = ~a41008 & ~a40758;
assign a44432 = a44430 & a41024;
assign a44434 = a44432 & a44414;
assign a44436 = a44434 & a40730;
assign a44438 = ~a44436 & ~a41926;
assign a44440 = a44436 & i744;
assign a44444 = a44434 & ~a40730;
assign a44446 = ~a44444 & ~a41958;
assign a44448 = a44444 & i744;
assign a44452 = a44416 & a40730;
assign a44454 = a44452 & a40758;
assign a44456 = a44454 & a41008;
assign a44458 = ~a44456 & ~a41996;
assign a44460 = a44456 & i744;
assign a44464 = a44418 & a40758;
assign a44466 = a44464 & a41008;
assign a44468 = ~a44466 & ~a42030;
assign a44470 = a44466 & i744;
assign a44474 = a44452 & ~a40758;
assign a44476 = a44474 & a41008;
assign a44478 = ~a44476 & ~a42062;
assign a44480 = a44476 & i744;
assign a44484 = a44420 & a41008;
assign a44486 = ~a44484 & ~a42096;
assign a44488 = a44484 & i744;
assign a44492 = a44454 & ~a41008;
assign a44494 = ~a44492 & ~a42116;
assign a44496 = a44492 & i744;
assign a44500 = a44464 & ~a41008;
assign a44502 = ~a44500 & ~a42138;
assign a44504 = a44500 & i744;
assign a44508 = a44474 & ~a41008;
assign a44510 = ~a44508 & ~a42158;
assign a44512 = a44508 & i744;
assign a44516 = ~a44422 & ~a42256;
assign a44518 = a44422 & i750;
assign a44522 = ~a44436 & ~a42282;
assign a44524 = a44436 & i750;
assign a44528 = ~a44444 & ~a42306;
assign a44530 = a44444 & i750;
assign a44534 = ~a44456 & ~a42330;
assign a44536 = a44456 & i750;
assign a44540 = ~a44466 & ~a42356;
assign a44542 = a44466 & i750;
assign a44546 = ~a44476 & ~a42380;
assign a44548 = a44476 & i750;
assign a44552 = ~a44484 & ~a42406;
assign a44554 = a44484 & i750;
assign a44558 = ~a44492 & ~a42424;
assign a44560 = a44492 & i750;
assign a44564 = ~a44500 & ~a42442;
assign a44566 = a44500 & i750;
assign a44570 = ~a44508 & ~a42460;
assign a44572 = a44508 & i750;
assign a44576 = ~a44422 & ~a42554;
assign a44578 = a44422 & i756;
assign a44582 = ~a44436 & ~a42580;
assign a44584 = a44436 & i756;
assign a44588 = ~a44444 & ~a42604;
assign a44590 = a44444 & i756;
assign a44594 = ~a44456 & ~a42628;
assign a44596 = a44456 & i756;
assign a44600 = ~a44466 & ~a42654;
assign a44602 = a44466 & i756;
assign a44606 = ~a44476 & ~a42678;
assign a44608 = a44476 & i756;
assign a44612 = ~a44484 & ~a42704;
assign a44614 = a44484 & i756;
assign a44618 = ~a44492 & ~a42722;
assign a44620 = a44492 & i756;
assign a44624 = ~a44500 & ~a42740;
assign a44626 = a44500 & i756;
assign a44630 = ~a44508 & ~a42758;
assign a44632 = a44508 & i756;
assign a44636 = ~a44422 & ~a42852;
assign a44638 = a44422 & i762;
assign a44642 = ~a44436 & ~a42878;
assign a44644 = a44436 & i762;
assign a44648 = ~a44444 & ~a42902;
assign a44650 = a44444 & i762;
assign a44654 = ~a44456 & ~a42926;
assign a44656 = a44456 & i762;
assign a44660 = ~a44466 & ~a42952;
assign a44662 = a44466 & i762;
assign a44666 = ~a44476 & ~a42976;
assign a44668 = a44476 & i762;
assign a44672 = ~a44484 & ~a43002;
assign a44674 = a44484 & i762;
assign a44678 = ~a44492 & ~a43020;
assign a44680 = a44492 & i762;
assign a44684 = ~a44500 & ~a43038;
assign a44686 = a44500 & i762;
assign a44690 = ~a44508 & ~a43056;
assign a44692 = a44508 & i762;
assign a44696 = ~a44422 & ~a43150;
assign a44698 = a44422 & i768;
assign a44702 = ~a44436 & ~a43176;
assign a44704 = a44436 & i768;
assign a44708 = ~a44444 & ~a43200;
assign a44710 = a44444 & i768;
assign a44714 = ~a44456 & ~a43224;
assign a44716 = a44456 & i768;
assign a44720 = ~a44466 & ~a43250;
assign a44722 = a44466 & i768;
assign a44726 = ~a44476 & ~a43274;
assign a44728 = a44476 & i768;
assign a44732 = ~a44484 & ~a43300;
assign a44734 = a44484 & i768;
assign a44738 = ~a44492 & ~a43318;
assign a44740 = a44492 & i768;
assign a44744 = ~a44500 & ~a43336;
assign a44746 = a44500 & i768;
assign a44750 = ~a44508 & ~a43354;
assign a44752 = a44508 & i768;
assign a44756 = ~a44422 & ~a43446;
assign a44758 = a44422 & i774;
assign a44762 = ~a44436 & ~a43472;
assign a44764 = a44436 & i774;
assign a44768 = ~a44444 & ~a43496;
assign a44770 = a44444 & i774;
assign a44774 = ~a44456 & ~a43520;
assign a44776 = a44456 & i774;
assign a44780 = ~a44466 & ~a43546;
assign a44782 = a44466 & i774;
assign a44786 = ~a44476 & ~a43570;
assign a44788 = a44476 & i774;
assign a44792 = ~a44484 & ~a43596;
assign a44794 = a44484 & i774;
assign a44798 = ~a44492 & ~a43614;
assign a44800 = a44492 & i774;
assign a44804 = ~a44500 & ~a43632;
assign a44806 = a44500 & i774;
assign a44810 = ~a44508 & ~a43650;
assign a44812 = a44508 & i774;
assign a44816 = ~a44500 & ~a43738;
assign a44818 = ~l2252 & l890;
assign a44820 = a41020 & a41004;
assign a44822 = a41004 & ~a40754;
assign a44824 = ~a44822 & a44820;
assign a44826 = ~a44824 & i670;
assign a44828 = ~a44826 & ~i648;
assign a44830 = ~a44828 & ~l890;
assign a44832 = ~a44830 & ~a44818;
assign a44836 = l2256 & ~l2254;
assign a44838 = l2266 & l2264;
assign a44840 = ~a44838 & ~a44836;
assign a44842 = l2270 & l2268;
assign a44844 = ~a44842 & a44840;
assign a44846 = l2272 & l2268;
assign a44848 = l2276 & ~l2254;
assign a44850 = l2274 & l2264;
assign a44852 = ~a44850 & ~a44848;
assign a44854 = a44852 & ~a44846;
assign a44856 = ~a44854 & a41678;
assign a44858 = a44856 & ~a44844;
assign a44860 = a44858 & ~a41742;
assign a44862 = l2284 & l2268;
assign a44864 = l2288 & ~l2254;
assign a44866 = l2286 & l2264;
assign a44868 = ~a44866 & ~a44864;
assign a44870 = a44868 & ~a44862;
assign a44872 = ~a44870 & a41660;
assign a44874 = a44872 & ~a44844;
assign a44876 = a44874 & ~a41742;
assign a44878 = a44876 & a41678;
assign a44880 = a44878 & a44854;
assign a44882 = ~a44854 & ~a41678;
assign a44884 = a44882 & a44876;
assign a44886 = ~a44884 & ~a44880;
assign a44888 = a44886 & ~a44860;
assign a44890 = l2296 & l2268;
assign a44892 = l2300 & ~l2254;
assign a44894 = l2298 & l2264;
assign a44896 = ~a44894 & ~a44892;
assign a44898 = a44896 & ~a44890;
assign a44900 = ~a44898 & a44872;
assign a44902 = a44900 & ~a41806;
assign a44904 = a44844 & a41742;
assign a44906 = a44904 & a44882;
assign a44908 = a44906 & a44872;
assign a44910 = ~a44908 & ~a44902;
assign a44912 = a44910 & a44888;
assign a44914 = a44854 & a44844;
assign a44916 = a44914 & a44898;
assign a44918 = a44916 & ~a41806;
assign a44920 = a44918 & a44870;
assign a44922 = ~a44844 & a41742;
assign a44924 = a44922 & ~a41678;
assign a44926 = ~a44924 & ~a44920;
assign a44928 = a44926 & a44912;
assign a44930 = a44844 & ~a41742;
assign a44932 = a44930 & a44854;
assign a44934 = a44872 & a41678;
assign a44936 = a44934 & a44898;
assign a44938 = a44936 & a44914;
assign a44940 = ~a44938 & ~a44932;
assign a44942 = a44918 & ~a41660;
assign a44944 = a44854 & ~a41678;
assign a44946 = a44944 & a41742;
assign a44948 = ~a44946 & ~a44942;
assign a44950 = a44948 & a44940;
assign a44952 = a44950 & a44928;
assign a44954 = ~a44952 & i674;
assign a44956 = ~l2308 & l890;
assign a44958 = ~a40578 & i560;
assign a44960 = a43826 & ~a40624;
assign a44962 = ~a41616 & ~a40624;
assign a44964 = a44962 & ~a44960;
assign a44966 = ~a41468 & a40578;
assign a44968 = ~a41478 & ~a40578;
assign a44970 = ~a44968 & ~a44966;
assign a44972 = ~a44970 & ~a43826;
assign a44974 = ~a41492 & a40578;
assign a44976 = ~a41468 & ~a40578;
assign a44978 = ~a44976 & ~a44974;
assign a44980 = ~a44978 & a43826;
assign a44982 = ~a44980 & ~a44972;
assign a44984 = a44982 & i610;
assign a44986 = ~a41420 & a40578;
assign a44988 = ~a41428 & ~a40578;
assign a44990 = ~a44988 & ~a44986;
assign a44992 = ~a44990 & ~a43826;
assign a44994 = ~a41442 & a40578;
assign a44996 = ~a41420 & ~a40578;
assign a44998 = ~a44996 & ~a44994;
assign a45000 = ~a44998 & a43826;
assign a45002 = ~a45000 & ~a44992;
assign a45004 = a45002 & i606;
assign a45006 = ~a45004 & ~a44984;
assign a45008 = ~a45002 & ~i606;
assign a45010 = ~a45008 & ~a45006;
assign a45012 = ~a41374 & a40578;
assign a45014 = ~a41382 & ~a40578;
assign a45016 = ~a45014 & ~a45012;
assign a45018 = ~a45016 & ~a43826;
assign a45020 = ~a41396 & a40578;
assign a45022 = ~a41374 & ~a40578;
assign a45024 = ~a45022 & ~a45020;
assign a45026 = ~a45024 & a43826;
assign a45028 = ~a45026 & ~a45018;
assign a45030 = a45028 & i600;
assign a45032 = ~a45030 & ~a45010;
assign a45034 = ~a45028 & ~i600;
assign a45036 = ~a45034 & ~a45032;
assign a45038 = ~a41328 & a40578;
assign a45040 = ~a41336 & ~a40578;
assign a45042 = ~a45040 & ~a45038;
assign a45044 = ~a45042 & ~a43826;
assign a45046 = ~a41350 & a40578;
assign a45048 = ~a41328 & ~a40578;
assign a45050 = ~a45048 & ~a45046;
assign a45052 = ~a45050 & a43826;
assign a45054 = ~a45052 & ~a45044;
assign a45056 = a45054 & i596;
assign a45058 = ~a45056 & ~a45036;
assign a45060 = ~a45054 & ~i596;
assign a45062 = ~a45060 & ~a45058;
assign a45064 = ~a41282 & a40578;
assign a45066 = ~a41290 & ~a40578;
assign a45068 = ~a45066 & ~a45064;
assign a45070 = ~a45068 & ~a43826;
assign a45072 = ~a41304 & a40578;
assign a45074 = ~a41282 & ~a40578;
assign a45076 = ~a45074 & ~a45072;
assign a45078 = ~a45076 & a43826;
assign a45080 = ~a45078 & ~a45070;
assign a45082 = a45080 & i594;
assign a45084 = ~a45082 & ~a45062;
assign a45086 = ~a45080 & ~i594;
assign a45088 = ~a45086 & ~a45084;
assign a45090 = ~a41236 & a40578;
assign a45092 = ~a41244 & ~a40578;
assign a45094 = ~a45092 & ~a45090;
assign a45096 = ~a45094 & ~a43826;
assign a45098 = ~a41258 & a40578;
assign a45100 = ~a41236 & ~a40578;
assign a45102 = ~a45100 & ~a45098;
assign a45104 = ~a45102 & a43826;
assign a45106 = ~a45104 & ~a45096;
assign a45108 = a45106 & i686;
assign a45110 = ~a45108 & ~a45088;
assign a45112 = ~a45106 & ~i686;
assign a45114 = ~a45112 & ~a45110;
assign a45116 = ~a41190 & a40578;
assign a45118 = ~a41198 & ~a40578;
assign a45120 = ~a45118 & ~a45116;
assign a45122 = ~a45120 & ~a43826;
assign a45124 = ~a41212 & a40578;
assign a45126 = ~a41190 & ~a40578;
assign a45128 = ~a45126 & ~a45124;
assign a45130 = ~a45128 & a43826;
assign a45132 = ~a45130 & ~a45122;
assign a45134 = a45132 & i690;
assign a45136 = ~a45134 & ~a45114;
assign a45138 = ~a45132 & ~i690;
assign a45140 = ~a45138 & ~a45136;
assign a45142 = ~a41144 & a40578;
assign a45144 = ~a41152 & ~a40578;
assign a45146 = ~a45144 & ~a45142;
assign a45148 = ~a45146 & ~a43826;
assign a45150 = ~a41166 & a40578;
assign a45152 = ~a41144 & ~a40578;
assign a45154 = ~a45152 & ~a45150;
assign a45156 = ~a45154 & a43826;
assign a45158 = ~a45156 & ~a45148;
assign a45160 = a45158 & i694;
assign a45162 = ~a45158 & ~i694;
assign a45164 = ~a45162 & ~a45160;
assign a45166 = ~a45164 & a45140;
assign a45168 = a45164 & ~a45134;
assign a45170 = ~a44982 & ~i610;
assign a45172 = ~a45170 & ~a45008;
assign a45174 = ~a45172 & ~a45004;
assign a45176 = ~a45174 & ~a45034;
assign a45178 = ~a45176 & ~a45030;
assign a45180 = ~a45178 & ~a45060;
assign a45182 = ~a45180 & ~a45056;
assign a45184 = ~a45182 & ~a45086;
assign a45186 = ~a45184 & ~a45082;
assign a45188 = ~a45186 & ~a45112;
assign a45190 = ~a45188 & ~a45108;
assign a45192 = ~a45190 & ~a45138;
assign a45194 = ~a45192 & a45168;
assign a45196 = ~a45194 & ~a45166;
assign a45198 = a41068 & a40578;
assign a45200 = a41090 & ~a40578;
assign a45202 = ~a45200 & ~a45198;
assign a45204 = ~a45202 & ~a43826;
assign a45206 = a41126 & a40578;
assign a45208 = a41068 & ~a40578;
assign a45210 = ~a45208 & ~a45206;
assign a45212 = ~a45210 & a43826;
assign a45214 = ~a45212 & ~a45204;
assign a45216 = ~a45214 & a45196;
assign a45218 = ~a45216 & ~i560;
assign a45220 = a45218 & ~a44964;
assign a45222 = ~a45220 & ~a44958;
assign a45224 = a45216 & ~i560;
assign a45226 = a45224 & a44964;
assign a45228 = ~a45226 & a45222;
assign a45230 = ~a45228 & ~l890;
assign a45232 = ~a45230 & ~a44956;
assign a45234 = ~l2366 & l890;
assign a45236 = a40578 & i560;
assign a45238 = a45224 & ~a44964;
assign a45240 = ~a45238 & ~a45236;
assign a45242 = ~a45240 & ~l890;
assign a45244 = ~a45242 & ~a45234;
assign a45246 = ~l2368 & l890;
assign a45248 = i792 & i648;
assign a45250 = i830 & ~i648;
assign a45252 = ~a45250 & ~a45248;
assign a45254 = ~a44964 & ~a42134;
assign a45256 = a44964 & ~a42154;
assign a45258 = ~a45256 & ~a45254;
assign a45260 = ~a45258 & ~a45216;
assign a45262 = ~a44964 & ~a42112;
assign a45264 = a44964 & ~a42134;
assign a45266 = ~a45264 & ~a45262;
assign a45268 = ~a45266 & a45216;
assign a45270 = ~a45268 & ~a45260;
assign a45272 = a45270 & a45252;
assign a45274 = i794 & i648;
assign a45276 = i832 & ~i648;
assign a45278 = ~a45276 & ~a45274;
assign a45280 = ~a44964 & ~a42438;
assign a45282 = a44964 & ~a42456;
assign a45284 = ~a45282 & ~a45280;
assign a45286 = ~a45284 & ~a45216;
assign a45288 = ~a44964 & ~a42420;
assign a45290 = a44964 & ~a42438;
assign a45292 = ~a45290 & ~a45288;
assign a45294 = ~a45292 & a45216;
assign a45296 = ~a45294 & ~a45286;
assign a45298 = a45296 & a45278;
assign a45300 = ~a45298 & ~a45272;
assign a45302 = ~a45296 & ~a45278;
assign a45304 = ~a45302 & ~a45300;
assign a45306 = i796 & i648;
assign a45308 = i834 & ~i648;
assign a45310 = ~a45308 & ~a45306;
assign a45312 = ~a44964 & ~a42736;
assign a45314 = a44964 & ~a42754;
assign a45316 = ~a45314 & ~a45312;
assign a45318 = ~a45316 & ~a45216;
assign a45320 = ~a44964 & ~a42718;
assign a45322 = a44964 & ~a42736;
assign a45324 = ~a45322 & ~a45320;
assign a45326 = ~a45324 & a45216;
assign a45328 = ~a45326 & ~a45318;
assign a45330 = a45328 & a45310;
assign a45332 = ~a45330 & ~a45304;
assign a45334 = ~a45328 & ~a45310;
assign a45336 = ~a45334 & ~a45332;
assign a45338 = i798 & i648;
assign a45340 = i836 & ~i648;
assign a45342 = ~a45340 & ~a45338;
assign a45344 = ~a44964 & ~a43034;
assign a45346 = a44964 & ~a43052;
assign a45348 = ~a45346 & ~a45344;
assign a45350 = ~a45348 & ~a45216;
assign a45352 = ~a44964 & ~a43016;
assign a45354 = a44964 & ~a43034;
assign a45356 = ~a45354 & ~a45352;
assign a45358 = ~a45356 & a45216;
assign a45360 = ~a45358 & ~a45350;
assign a45362 = a45360 & a45342;
assign a45364 = ~a45362 & ~a45336;
assign a45366 = ~a45360 & ~a45342;
assign a45368 = ~a45366 & ~a45364;
assign a45370 = i800 & i648;
assign a45372 = i838 & ~i648;
assign a45374 = ~a45372 & ~a45370;
assign a45376 = ~a44964 & ~a43332;
assign a45378 = a44964 & ~a43350;
assign a45380 = ~a45378 & ~a45376;
assign a45382 = ~a45380 & ~a45216;
assign a45384 = ~a44964 & ~a43314;
assign a45386 = a44964 & ~a43332;
assign a45388 = ~a45386 & ~a45384;
assign a45390 = ~a45388 & a45216;
assign a45392 = ~a45390 & ~a45382;
assign a45394 = a45392 & a45374;
assign a45396 = ~a45394 & ~a45368;
assign a45398 = ~a45392 & ~a45374;
assign a45400 = ~a45398 & ~a45396;
assign a45402 = i802 & i648;
assign a45404 = i840 & ~i648;
assign a45406 = ~a45404 & ~a45402;
assign a45408 = ~a44964 & ~a43628;
assign a45410 = a44964 & ~a43646;
assign a45412 = ~a45410 & ~a45408;
assign a45414 = ~a45412 & ~a45216;
assign a45416 = ~a44964 & ~a43610;
assign a45418 = a44964 & ~a43628;
assign a45420 = ~a45418 & ~a45416;
assign a45422 = ~a45420 & a45216;
assign a45424 = ~a45422 & ~a45414;
assign a45426 = a45424 & a45406;
assign a45428 = ~a45426 & ~a45400;
assign a45430 = ~a45424 & ~a45406;
assign a45432 = ~a45430 & ~a45428;
assign a45434 = i804 & i648;
assign a45436 = i842 & ~i648;
assign a45438 = ~a45436 & ~a45434;
assign a45440 = ~a42128 & ~a41190;
assign a45442 = a42128 & i822;
assign a45444 = ~a45442 & ~a45440;
assign a45446 = ~a45444 & ~a44964;
assign a45448 = ~a42148 & ~a41198;
assign a45450 = a42148 & i822;
assign a45452 = ~a45450 & ~a45448;
assign a45454 = ~a45452 & a44964;
assign a45456 = ~a45454 & ~a45446;
assign a45458 = ~a45456 & ~a45216;
assign a45460 = ~a42106 & ~a41212;
assign a45462 = a42106 & i822;
assign a45464 = ~a45462 & ~a45460;
assign a45466 = ~a45464 & ~a44964;
assign a45468 = ~a45444 & a44964;
assign a45470 = ~a45468 & ~a45466;
assign a45472 = ~a45470 & a45216;
assign a45474 = ~a45472 & ~a45458;
assign a45476 = a45474 & a45438;
assign a45478 = ~a45476 & ~a45432;
assign a45480 = ~a45474 & ~a45438;
assign a45482 = ~a45480 & ~a45478;
assign a45484 = i790 & i648;
assign a45486 = i844 & ~i648;
assign a45488 = ~a45486 & ~a45484;
assign a45490 = ~a42128 & ~a41144;
assign a45492 = a42128 & i826;
assign a45494 = ~a45492 & ~a45490;
assign a45496 = ~a45494 & ~a44964;
assign a45498 = ~a42148 & ~a41152;
assign a45500 = a42148 & i826;
assign a45502 = ~a45500 & ~a45498;
assign a45504 = ~a45502 & a44964;
assign a45506 = ~a45504 & ~a45496;
assign a45508 = ~a45506 & ~a45216;
assign a45510 = ~a42106 & ~a41166;
assign a45512 = a42106 & i826;
assign a45514 = ~a45512 & ~a45510;
assign a45516 = ~a45514 & ~a44964;
assign a45518 = ~a45494 & a44964;
assign a45520 = ~a45518 & ~a45516;
assign a45522 = ~a45520 & a45216;
assign a45524 = ~a45522 & ~a45508;
assign a45526 = a45524 & a45488;
assign a45528 = ~a45524 & ~a45488;
assign a45530 = ~a45528 & ~a45526;
assign a45532 = ~a45530 & a45482;
assign a45534 = a45530 & ~a45476;
assign a45536 = ~a45270 & ~a45252;
assign a45538 = ~a45536 & ~a45302;
assign a45540 = ~a45538 & ~a45298;
assign a45542 = ~a45540 & ~a45334;
assign a45544 = ~a45542 & ~a45330;
assign a45546 = ~a45544 & ~a45366;
assign a45548 = ~a45546 & ~a45362;
assign a45550 = ~a45548 & ~a45398;
assign a45552 = ~a45550 & ~a45394;
assign a45554 = ~a45552 & ~a45430;
assign a45556 = ~a45554 & ~a45426;
assign a45558 = ~a45556 & ~a45480;
assign a45560 = ~a45558 & a45534;
assign a45562 = ~a45560 & ~a45532;
assign a45564 = ~a44964 & a43734;
assign a45566 = a44964 & a43862;
assign a45568 = ~a45566 & ~a45564;
assign a45570 = ~a45568 & ~a45216;
assign a45572 = ~a44964 & a44058;
assign a45574 = a44964 & a43734;
assign a45576 = ~a45574 & ~a45572;
assign a45578 = ~a45576 & a45216;
assign a45580 = ~a45578 & ~a45570;
assign a45582 = ~a45580 & a45562;
assign a45584 = ~a45582 & ~l890;
assign a45586 = ~a45584 & ~a45246;
assign a45588 = a45586 & ~a45244;
assign a45590 = a45588 & ~l2370;
assign a45592 = a45590 & a45232;
assign a45594 = ~a45592 & ~a44954;
assign a45598 = ~l2292 & l890;
assign a45600 = ~l890 & i622;
assign a45602 = ~a45600 & ~a45598;
assign a45604 = ~l2294 & l890;
assign a45606 = ~l890 & ~i554;
assign a45610 = a41644 & a41626;
assign a45612 = ~a45586 & ~a41644;
assign a45614 = a45612 & ~a45232;
assign a45616 = a45586 & ~a41644;
assign a45618 = a45616 & a45232;
assign a45620 = ~a45618 & ~a45614;
assign a45624 = ~l2312 & l890;
assign a45626 = ~a41852 & a41550;
assign a45628 = a41852 & i710;
assign a45630 = ~a45628 & ~a45626;
assign a45632 = ~a45630 & a40578;
assign a45634 = a41902 & i642;
assign a45636 = a45634 & ~a41896;
assign a45638 = a41896 & i710;
assign a45640 = ~a45638 & ~a45636;
assign a45642 = ~a45640 & ~a40578;
assign a45644 = ~a45642 & ~a45632;
assign a45646 = ~a45644 & a41612;
assign a45648 = ~a41152 & a40578;
assign a45650 = ~a45630 & ~a40578;
assign a45652 = ~a45650 & ~a45648;
assign a45654 = ~a45652 & a41614;
assign a45656 = ~a45654 & ~a45646;
assign a45658 = ~a45146 & ~a40982;
assign a45660 = ~a45658 & a45656;
assign a45662 = a45660 & ~i790;
assign a45664 = ~a45660 & i790;
assign a45666 = ~a45664 & ~a45662;
assign a45668 = ~a41860 & a40578;
assign a45670 = ~a41910 & ~a40578;
assign a45672 = ~a45670 & ~a45668;
assign a45674 = ~a45672 & a41612;
assign a45676 = ~a41478 & a40578;
assign a45678 = ~a41860 & ~a40578;
assign a45680 = ~a45678 & ~a45676;
assign a45682 = ~a45680 & a41614;
assign a45684 = ~a45682 & ~a45674;
assign a45686 = ~a44970 & ~a40982;
assign a45688 = ~a45686 & a45684;
assign a45690 = ~a45688 & i792;
assign a45692 = ~a42246 & a40578;
assign a45694 = ~a42272 & ~a40578;
assign a45696 = ~a45694 & ~a45692;
assign a45698 = ~a45696 & a41612;
assign a45700 = ~a41428 & a40578;
assign a45702 = ~a42246 & ~a40578;
assign a45704 = ~a45702 & ~a45700;
assign a45706 = ~a45704 & a41614;
assign a45708 = ~a45706 & ~a45698;
assign a45710 = ~a44990 & ~a40982;
assign a45712 = ~a45710 & a45708;
assign a45714 = ~a45712 & i794;
assign a45716 = ~a45714 & ~a45690;
assign a45718 = a45712 & ~i794;
assign a45720 = ~a45718 & ~a45716;
assign a45722 = ~a42544 & a40578;
assign a45724 = ~a42570 & ~a40578;
assign a45726 = ~a45724 & ~a45722;
assign a45728 = ~a45726 & a41612;
assign a45730 = ~a41382 & a40578;
assign a45732 = ~a42544 & ~a40578;
assign a45734 = ~a45732 & ~a45730;
assign a45736 = ~a45734 & a41614;
assign a45738 = ~a45736 & ~a45728;
assign a45740 = ~a45016 & ~a40982;
assign a45742 = ~a45740 & a45738;
assign a45744 = ~a45742 & i796;
assign a45746 = ~a45744 & ~a45720;
assign a45748 = a45742 & ~i796;
assign a45750 = ~a45748 & ~a45746;
assign a45752 = ~a42842 & a40578;
assign a45754 = ~a42868 & ~a40578;
assign a45756 = ~a45754 & ~a45752;
assign a45758 = ~a45756 & a41612;
assign a45760 = ~a41336 & a40578;
assign a45762 = ~a42842 & ~a40578;
assign a45764 = ~a45762 & ~a45760;
assign a45766 = ~a45764 & a41614;
assign a45768 = ~a45766 & ~a45758;
assign a45770 = ~a45042 & ~a40982;
assign a45772 = ~a45770 & a45768;
assign a45774 = ~a45772 & i798;
assign a45776 = ~a45774 & ~a45750;
assign a45778 = a45772 & ~i798;
assign a45780 = ~a45778 & ~a45776;
assign a45782 = ~a43140 & a40578;
assign a45784 = ~a43166 & ~a40578;
assign a45786 = ~a45784 & ~a45782;
assign a45788 = ~a45786 & a41612;
assign a45790 = ~a41290 & a40578;
assign a45792 = ~a43140 & ~a40578;
assign a45794 = ~a45792 & ~a45790;
assign a45796 = ~a45794 & a41614;
assign a45798 = ~a45796 & ~a45788;
assign a45800 = ~a45068 & ~a40982;
assign a45802 = ~a45800 & a45798;
assign a45804 = ~a45802 & i800;
assign a45806 = ~a45804 & ~a45780;
assign a45808 = a45802 & ~i800;
assign a45810 = ~a45808 & ~a45806;
assign a45812 = ~a43436 & a40578;
assign a45814 = ~a43462 & ~a40578;
assign a45816 = ~a45814 & ~a45812;
assign a45818 = ~a45816 & a41612;
assign a45820 = ~a41244 & a40578;
assign a45822 = ~a43436 & ~a40578;
assign a45824 = ~a45822 & ~a45820;
assign a45826 = ~a45824 & a41614;
assign a45828 = ~a45826 & ~a45818;
assign a45830 = ~a45094 & ~a40982;
assign a45832 = ~a45830 & a45828;
assign a45834 = ~a45832 & i802;
assign a45836 = ~a45834 & ~a45810;
assign a45838 = a45832 & ~i802;
assign a45840 = ~a45838 & ~a45836;
assign a45842 = ~a41852 & a41580;
assign a45844 = a41852 & i714;
assign a45846 = ~a45844 & ~a45842;
assign a45848 = ~a45846 & a40578;
assign a45850 = a41902 & i638;
assign a45852 = a45850 & ~a41896;
assign a45854 = a41896 & i714;
assign a45856 = ~a45854 & ~a45852;
assign a45858 = ~a45856 & ~a40578;
assign a45860 = ~a45858 & ~a45848;
assign a45862 = ~a45860 & a41612;
assign a45864 = ~a41198 & a40578;
assign a45866 = ~a45846 & ~a40578;
assign a45868 = ~a45866 & ~a45864;
assign a45870 = ~a45868 & a41614;
assign a45872 = ~a45870 & ~a45862;
assign a45874 = ~a45120 & ~a40982;
assign a45876 = ~a45874 & a45872;
assign a45878 = ~a45876 & i804;
assign a45880 = ~a45878 & ~a45840;
assign a45882 = ~a45880 & a45666;
assign a45884 = a45876 & ~i804;
assign a45886 = ~a45884 & a45882;
assign a45888 = ~a45878 & ~a45666;
assign a45890 = a45688 & ~i792;
assign a45892 = ~a45890 & ~a45718;
assign a45894 = ~a45892 & ~a45714;
assign a45896 = ~a45894 & ~a45748;
assign a45898 = ~a45896 & ~a45744;
assign a45900 = ~a45898 & ~a45778;
assign a45902 = ~a45900 & ~a45774;
assign a45904 = ~a45902 & ~a45808;
assign a45906 = ~a45904 & ~a45804;
assign a45908 = ~a45906 & ~a45838;
assign a45910 = ~a45908 & ~a45834;
assign a45912 = ~a45910 & ~a45884;
assign a45914 = ~a45912 & a45888;
assign a45916 = ~a45914 & ~a45886;
assign a45918 = ~a45916 & ~i560;
assign a45920 = a43832 & a40578;
assign a45922 = a43894 & ~a40578;
assign a45924 = ~a45922 & ~a45920;
assign a45926 = ~a45924 & a41612;
assign a45928 = ~a45202 & ~a40982;
assign a45930 = ~a45928 & ~a45926;
assign a45932 = a41090 & a40578;
assign a45934 = a43832 & ~a40578;
assign a45936 = ~a45934 & ~a45932;
assign a45938 = ~a45936 & a41614;
assign a45940 = ~a45938 & a45930;
assign a45942 = ~a45940 & a45918;
assign a45944 = ~a45942 & ~l890;
assign a45946 = ~a45944 & ~a45624;
assign a45948 = a45946 & a41626;
assign a45950 = ~a41718 & ~a41024;
assign a45952 = a41718 & a41024;
assign a45954 = ~a45952 & ~a45950;
assign a45956 = a41008 & ~l2318;
assign a45958 = ~a45956 & a45954;
assign a45960 = ~a41008 & l2318;
assign a45962 = ~a45960 & a45958;
assign a45964 = a41710 & a40758;
assign a45966 = ~a45964 & a45962;
assign a45968 = ~a41710 & ~a40758;
assign a45970 = ~a45968 & a45966;
assign a45972 = a41626 & a40730;
assign a45974 = ~a45972 & a45970;
assign a45976 = ~a41626 & ~a40730;
assign a45978 = ~a45976 & a45974;
assign a45980 = ~l2320 & l890;
assign a45982 = ~a45652 & a41612;
assign a45984 = ~a45146 & a41614;
assign a45986 = ~a45984 & ~a45982;
assign a45988 = ~a45154 & ~a40982;
assign a45990 = ~a45988 & a45986;
assign a45992 = a45990 & ~i790;
assign a45994 = ~a45990 & i790;
assign a45996 = ~a45994 & ~a45992;
assign a45998 = ~a45868 & a41612;
assign a46000 = ~a45120 & a41614;
assign a46002 = ~a46000 & ~a45998;
assign a46004 = ~a45128 & ~a40982;
assign a46006 = ~a46004 & a46002;
assign a46008 = a46006 & ~i804;
assign a46010 = ~a46008 & a45996;
assign a46012 = ~a46006 & i804;
assign a46014 = ~a45824 & a41612;
assign a46016 = ~a45094 & a41614;
assign a46018 = ~a46016 & ~a46014;
assign a46020 = ~a45102 & ~a40982;
assign a46022 = ~a46020 & a46018;
assign a46024 = a46022 & ~i802;
assign a46026 = ~a46022 & i802;
assign a46028 = ~a45794 & a41612;
assign a46030 = ~a45068 & a41614;
assign a46032 = ~a46030 & ~a46028;
assign a46034 = ~a45076 & ~a40982;
assign a46036 = ~a46034 & a46032;
assign a46038 = a46036 & ~i800;
assign a46040 = ~a46036 & i800;
assign a46042 = ~a45764 & a41612;
assign a46044 = ~a45042 & a41614;
assign a46046 = ~a46044 & ~a46042;
assign a46048 = ~a45050 & ~a40982;
assign a46050 = ~a46048 & a46046;
assign a46052 = a46050 & ~i798;
assign a46054 = ~a46050 & i798;
assign a46056 = ~a45734 & a41612;
assign a46058 = ~a45016 & a41614;
assign a46060 = ~a46058 & ~a46056;
assign a46062 = ~a45024 & ~a40982;
assign a46064 = ~a46062 & a46060;
assign a46066 = a46064 & ~i796;
assign a46068 = ~a46064 & i796;
assign a46070 = ~a45704 & a41612;
assign a46072 = ~a44990 & a41614;
assign a46074 = ~a46072 & ~a46070;
assign a46076 = ~a44998 & ~a40982;
assign a46078 = ~a46076 & a46074;
assign a46080 = a46078 & ~i794;
assign a46082 = ~a46078 & i794;
assign a46084 = ~a45680 & a41612;
assign a46086 = ~a44970 & a41614;
assign a46088 = ~a46086 & ~a46084;
assign a46090 = ~a44978 & ~a40982;
assign a46092 = ~a46090 & a46088;
assign a46094 = ~a46092 & i792;
assign a46096 = ~a46094 & ~a46082;
assign a46098 = ~a46096 & ~a46080;
assign a46100 = ~a46098 & ~a46068;
assign a46102 = ~a46100 & ~a46066;
assign a46104 = ~a46102 & ~a46054;
assign a46106 = ~a46104 & ~a46052;
assign a46108 = ~a46106 & ~a46040;
assign a46110 = ~a46108 & ~a46038;
assign a46112 = ~a46110 & ~a46026;
assign a46114 = ~a46112 & ~a46024;
assign a46116 = ~a46114 & ~a46012;
assign a46118 = ~a46116 & a46010;
assign a46120 = ~a45210 & ~a40982;
assign a46122 = ~a46120 & ~a41612;
assign a46124 = ~a45202 & a41614;
assign a46126 = ~a46124 & a46122;
assign a46128 = ~a46126 & ~a46118;
assign a46130 = a46092 & ~i792;
assign a46132 = ~a46130 & ~a46080;
assign a46134 = ~a46132 & ~a46082;
assign a46136 = ~a46134 & ~a46066;
assign a46138 = ~a46136 & ~a46068;
assign a46140 = ~a46138 & ~a46052;
assign a46142 = ~a46140 & ~a46054;
assign a46144 = ~a46142 & ~a46038;
assign a46146 = ~a46144 & ~a46040;
assign a46148 = ~a46146 & ~a46024;
assign a46150 = ~a46148 & ~a46026;
assign a46152 = ~a46150 & ~a46008;
assign a46154 = ~a46152 & ~a46012;
assign a46156 = a46154 & ~a45996;
assign a46158 = ~a46156 & a46128;
assign a46160 = ~a46158 & ~l890;
assign a46162 = ~a46160 & ~a45980;
assign a46164 = a46162 & ~a45978;
assign a46166 = ~a46164 & ~a40648;
assign a46168 = a46166 & ~a45946;
assign a46170 = a46168 & ~a41626;
assign a46172 = ~a46166 & a41626;
assign a46174 = ~a46172 & ~a46170;
assign a46178 = a41718 & a41710;
assign a46180 = ~l2342 & l890;
assign a46182 = ~a45502 & ~l890;
assign a46184 = ~a46182 & ~a46180;
assign a46186 = ~a46184 & ~l2318;
assign a46188 = a46186 & ~a41626;
assign a46190 = a46188 & a46178;
assign a46192 = a41718 & a41626;
assign a46194 = a46192 & ~l2318;
assign a46196 = a46194 & a41710;
assign a46198 = ~l2344 & l890;
assign a46200 = ~a45630 & ~a41868;
assign a46202 = a41868 & i826;
assign a46204 = ~a46202 & ~a46200;
assign a46206 = ~a46204 & ~l890;
assign a46208 = ~a46206 & ~a46198;
assign a46210 = ~a46208 & a46196;
assign a46212 = ~a46210 & ~a46190;
assign a46214 = a41718 & ~l2318;
assign a46216 = ~l2346 & l890;
assign a46218 = ~a45494 & ~l890;
assign a46220 = ~a46218 & ~a46216;
assign a46222 = ~a46220 & a46214;
assign a46224 = a46222 & ~a41710;
assign a46226 = a46224 & a41626;
assign a46228 = ~a46226 & a46212;
assign a46230 = ~l2348 & l890;
assign a46232 = ~a45514 & ~l890;
assign a46234 = ~a46232 & ~a46230;
assign a46236 = ~a46234 & a46214;
assign a46238 = a46236 & ~a41710;
assign a46240 = a46238 & ~a41626;
assign a46242 = ~a46240 & a46228;
assign a46244 = a46192 & l2318;
assign a46246 = a46244 & a41710;
assign a46248 = ~l2350 & l890;
assign a46250 = a42074 & i642;
assign a46252 = a46250 & ~a42078;
assign a46254 = a42078 & i710;
assign a46256 = ~a46254 & ~a46252;
assign a46258 = ~a46256 & ~a42086;
assign a46260 = a42086 & i826;
assign a46262 = ~a46260 & ~a46258;
assign a46264 = ~a46262 & ~l890;
assign a46266 = ~a46264 & ~a46248;
assign a46268 = ~a46266 & a46246;
assign a46270 = ~a46268 & a46242;
assign a46272 = ~l2352 & l890;
assign a46274 = a42038 & i642;
assign a46276 = a46274 & ~a42042;
assign a46278 = a42042 & i710;
assign a46280 = ~a46278 & ~a46276;
assign a46282 = ~a46280 & ~a42052;
assign a46284 = a42052 & i826;
assign a46286 = ~a46284 & ~a46282;
assign a46288 = ~a46286 & ~l890;
assign a46290 = ~a46288 & ~a46272;
assign a46292 = ~a46290 & a41718;
assign a46294 = a46292 & l2318;
assign a46296 = a46294 & a41720;
assign a46298 = ~a46296 & a46270;
assign a46300 = a41718 & l2318;
assign a46302 = ~l2354 & l890;
assign a46304 = a42006 & i642;
assign a46306 = a46304 & ~a42010;
assign a46308 = a42010 & i710;
assign a46310 = ~a46308 & ~a46306;
assign a46312 = ~a46310 & ~a42020;
assign a46314 = a42020 & i826;
assign a46316 = ~a46314 & ~a46312;
assign a46318 = ~a46316 & ~l890;
assign a46320 = ~a46318 & ~a46302;
assign a46322 = ~a46320 & a46300;
assign a46324 = a46322 & a41712;
assign a46326 = ~a46324 & a46298;
assign a46328 = ~l2356 & l890;
assign a46330 = a41970 & i642;
assign a46332 = a46330 & ~a41974;
assign a46334 = a41974 & i710;
assign a46336 = ~a46334 & ~a46332;
assign a46338 = ~a46336 & ~a41986;
assign a46340 = a41986 & i826;
assign a46342 = ~a46340 & ~a46338;
assign a46344 = ~a46342 & ~l890;
assign a46346 = ~a46344 & ~a46328;
assign a46348 = ~a46346 & a46300;
assign a46350 = a46348 & ~a41626;
assign a46352 = a46350 & ~a41710;
assign a46354 = ~a46352 & a46326;
assign a46356 = ~a41718 & ~l2318;
assign a46358 = ~l2358 & l890;
assign a46360 = a41936 & i642;
assign a46362 = a46360 & ~a41940;
assign a46364 = a41940 & i710;
assign a46366 = ~a46364 & ~a46362;
assign a46368 = ~a46366 & ~a41948;
assign a46370 = a41948 & i826;
assign a46372 = ~a46370 & ~a46368;
assign a46374 = ~a46372 & ~l890;
assign a46376 = ~a46374 & ~a46358;
assign a46378 = ~a46376 & a46356;
assign a46380 = a46378 & a41626;
assign a46382 = ~a46380 & a46354;
assign a46384 = ~l2360 & l890;
assign a46386 = ~a45640 & ~a41916;
assign a46388 = a41916 & i826;
assign a46390 = ~a46388 & ~a46386;
assign a46392 = ~a46390 & ~l890;
assign a46394 = ~a46392 & ~a46384;
assign a46396 = ~a46394 & a46356;
assign a46398 = a46396 & ~a41626;
assign a46400 = ~a46398 & a46382;
assign a46402 = ~a46400 & a46168;
assign a46404 = a46222 & a41720;
assign a46406 = a46196 & ~a46184;
assign a46408 = ~a46406 & ~a46404;
assign a46410 = a46238 & a41626;
assign a46412 = ~a46410 & a46408;
assign a46414 = ~a41710 & ~l2318;
assign a46416 = ~a46266 & a41718;
assign a46418 = a46416 & a46414;
assign a46420 = a46418 & ~a41626;
assign a46422 = ~a46420 & a46412;
assign a46424 = ~a46290 & a46246;
assign a46426 = ~a46424 & a46422;
assign a46428 = a46322 & ~a41626;
assign a46430 = a46428 & a41710;
assign a46432 = ~a46430 & a46426;
assign a46434 = a46348 & a41712;
assign a46436 = ~a46434 & a46432;
assign a46438 = ~a41710 & l2318;
assign a46440 = a46438 & a41718;
assign a46442 = a46440 & ~a46376;
assign a46444 = a46442 & ~a41626;
assign a46446 = ~a46444 & a46436;
assign a46448 = a46396 & a41626;
assign a46450 = ~a46448 & a46446;
assign a46452 = ~a46208 & ~l2318;
assign a46454 = a46452 & ~a41718;
assign a46456 = a46454 & ~a41626;
assign a46458 = ~a46456 & a46450;
assign a46460 = ~a46458 & ~a46166;
assign a46462 = ~a46460 & ~a46402;
assign a46464 = a46452 & a41722;
assign a46466 = ~a46394 & a46196;
assign a46468 = ~a46466 & ~a46464;
assign a46470 = a41718 & a41712;
assign a46472 = a46470 & a46186;
assign a46474 = ~a46472 & a46468;
assign a46476 = a46224 & ~a41626;
assign a46478 = ~a46476 & a46474;
assign a46480 = a46246 & ~a46234;
assign a46482 = ~a46480 & a46478;
assign a46484 = ~a41626 & l2318;
assign a46486 = a46484 & a41710;
assign a46488 = a46486 & a46416;
assign a46490 = ~a46488 & a46482;
assign a46492 = a46294 & a41712;
assign a46494 = ~a46492 & a46490;
assign a46496 = a46428 & ~a41710;
assign a46498 = ~a46496 & a46494;
assign a46500 = a41830 & ~l2318;
assign a46502 = a46500 & ~a46346;
assign a46504 = ~a46502 & a46498;
assign a46506 = a46378 & ~a41626;
assign a46508 = ~a46506 & a46504;
assign a46510 = ~a46508 & a45946;
assign a46512 = ~a46510 & a46462;
assign a46514 = a46512 & ~i806;
assign a46516 = ~a46512 & i806;
assign a46518 = ~a46516 & ~a46514;
assign a46520 = ~a42158 & ~l2318;
assign a46522 = a46520 & ~a41626;
assign a46524 = a46522 & a46178;
assign a46526 = a46196 & ~a41878;
assign a46528 = ~a46526 & ~a46524;
assign a46530 = a46214 & ~a42138;
assign a46532 = a46530 & ~a41710;
assign a46534 = a46532 & a41626;
assign a46536 = ~a46534 & a46528;
assign a46538 = a46214 & ~a42116;
assign a46540 = a46538 & ~a41710;
assign a46542 = a46540 & ~a41626;
assign a46544 = ~a46542 & a46536;
assign a46546 = a46246 & ~a42096;
assign a46548 = ~a46546 & a46544;
assign a46550 = ~a42062 & a41718;
assign a46552 = a46550 & l2318;
assign a46554 = a46552 & a41720;
assign a46556 = ~a46554 & a46548;
assign a46558 = a46300 & ~a42030;
assign a46560 = a46558 & a41712;
assign a46562 = ~a46560 & a46556;
assign a46564 = a46300 & ~a41996;
assign a46566 = a46564 & ~a41626;
assign a46568 = a46566 & ~a41710;
assign a46570 = ~a46568 & a46562;
assign a46572 = a46356 & ~a41958;
assign a46574 = a46572 & a41626;
assign a46576 = ~a46574 & a46570;
assign a46578 = a46356 & ~a41926;
assign a46580 = a46578 & ~a41626;
assign a46582 = ~a46580 & a46576;
assign a46584 = ~a46582 & a46168;
assign a46586 = a46530 & a41720;
assign a46588 = a46196 & ~a42158;
assign a46590 = ~a46588 & ~a46586;
assign a46592 = a46540 & a41626;
assign a46594 = ~a46592 & a46590;
assign a46596 = ~a42096 & a41718;
assign a46598 = a46596 & a46414;
assign a46600 = a46598 & ~a41626;
assign a46602 = ~a46600 & a46594;
assign a46604 = a46246 & ~a42062;
assign a46606 = ~a46604 & a46602;
assign a46608 = a46558 & ~a41626;
assign a46610 = a46608 & a41710;
assign a46612 = ~a46610 & a46606;
assign a46614 = a46564 & a41712;
assign a46616 = ~a46614 & a46612;
assign a46618 = a46440 & ~a41958;
assign a46620 = a46618 & ~a41626;
assign a46622 = ~a46620 & a46616;
assign a46624 = a46578 & a41626;
assign a46626 = ~a46624 & a46622;
assign a46628 = ~a41878 & ~l2318;
assign a46630 = a46628 & ~a41718;
assign a46632 = a46630 & ~a41626;
assign a46634 = ~a46632 & a46626;
assign a46636 = ~a46634 & ~a46166;
assign a46638 = ~a46636 & ~a46584;
assign a46640 = a46628 & a41722;
assign a46642 = a46196 & ~a41926;
assign a46644 = ~a46642 & ~a46640;
assign a46646 = a46520 & a46470;
assign a46648 = ~a46646 & a46644;
assign a46650 = a46532 & ~a41626;
assign a46652 = ~a46650 & a46648;
assign a46654 = a46246 & ~a42116;
assign a46656 = ~a46654 & a46652;
assign a46658 = a46596 & a46486;
assign a46660 = ~a46658 & a46656;
assign a46662 = a46552 & a41712;
assign a46664 = ~a46662 & a46660;
assign a46666 = a46608 & ~a41710;
assign a46668 = ~a46666 & a46664;
assign a46670 = a46500 & ~a41996;
assign a46672 = ~a46670 & a46668;
assign a46674 = a46572 & ~a41626;
assign a46676 = ~a46674 & a46672;
assign a46678 = ~a46676 & a45946;
assign a46680 = ~a46678 & a46638;
assign a46682 = ~a46680 & i808;
assign a46684 = ~a42460 & ~l2318;
assign a46686 = a46684 & ~a41626;
assign a46688 = a46686 & a46178;
assign a46690 = a46196 & ~a42256;
assign a46692 = ~a46690 & ~a46688;
assign a46694 = a46214 & ~a42442;
assign a46696 = a46694 & ~a41710;
assign a46698 = a46696 & a41626;
assign a46700 = ~a46698 & a46692;
assign a46702 = a46214 & ~a42424;
assign a46704 = a46702 & ~a41710;
assign a46706 = a46704 & ~a41626;
assign a46708 = ~a46706 & a46700;
assign a46710 = a46246 & ~a42406;
assign a46712 = ~a46710 & a46708;
assign a46714 = ~a42380 & a41718;
assign a46716 = a46714 & l2318;
assign a46718 = a46716 & a41720;
assign a46720 = ~a46718 & a46712;
assign a46722 = a46300 & ~a42356;
assign a46724 = a46722 & a41712;
assign a46726 = ~a46724 & a46720;
assign a46728 = a46300 & ~a42330;
assign a46730 = a46728 & ~a41626;
assign a46732 = a46730 & ~a41710;
assign a46734 = ~a46732 & a46726;
assign a46736 = a46356 & ~a42306;
assign a46738 = a46736 & a41626;
assign a46740 = ~a46738 & a46734;
assign a46742 = a46356 & ~a42282;
assign a46744 = a46742 & ~a41626;
assign a46746 = ~a46744 & a46740;
assign a46748 = ~a46746 & a46168;
assign a46750 = a46694 & a41720;
assign a46752 = a46196 & ~a42460;
assign a46754 = ~a46752 & ~a46750;
assign a46756 = a46704 & a41626;
assign a46758 = ~a46756 & a46754;
assign a46760 = ~a42406 & a41718;
assign a46762 = a46760 & a46414;
assign a46764 = a46762 & ~a41626;
assign a46766 = ~a46764 & a46758;
assign a46768 = a46246 & ~a42380;
assign a46770 = ~a46768 & a46766;
assign a46772 = a46722 & ~a41626;
assign a46774 = a46772 & a41710;
assign a46776 = ~a46774 & a46770;
assign a46778 = a46728 & a41712;
assign a46780 = ~a46778 & a46776;
assign a46782 = a46440 & ~a42306;
assign a46784 = a46782 & ~a41626;
assign a46786 = ~a46784 & a46780;
assign a46788 = a46742 & a41626;
assign a46790 = ~a46788 & a46786;
assign a46792 = ~a42256 & ~l2318;
assign a46794 = a46792 & ~a41718;
assign a46796 = a46794 & ~a41626;
assign a46798 = ~a46796 & a46790;
assign a46800 = ~a46798 & ~a46166;
assign a46802 = ~a46800 & ~a46748;
assign a46804 = a46792 & a41722;
assign a46806 = a46196 & ~a42282;
assign a46808 = ~a46806 & ~a46804;
assign a46810 = a46684 & a46470;
assign a46812 = ~a46810 & a46808;
assign a46814 = a46696 & ~a41626;
assign a46816 = ~a46814 & a46812;
assign a46818 = a46246 & ~a42424;
assign a46820 = ~a46818 & a46816;
assign a46822 = a46760 & a46486;
assign a46824 = ~a46822 & a46820;
assign a46826 = a46716 & a41712;
assign a46828 = ~a46826 & a46824;
assign a46830 = a46772 & ~a41710;
assign a46832 = ~a46830 & a46828;
assign a46834 = a46500 & ~a42330;
assign a46836 = ~a46834 & a46832;
assign a46838 = a46736 & ~a41626;
assign a46840 = ~a46838 & a46836;
assign a46842 = ~a46840 & a45946;
assign a46844 = ~a46842 & a46802;
assign a46846 = ~a46844 & i810;
assign a46848 = ~a46846 & ~a46682;
assign a46850 = a46844 & ~i810;
assign a46852 = ~a46850 & ~a46848;
assign a46854 = ~a42758 & ~l2318;
assign a46856 = a46854 & ~a41626;
assign a46858 = a46856 & a46178;
assign a46860 = a46196 & ~a42554;
assign a46862 = ~a46860 & ~a46858;
assign a46864 = a46214 & ~a42740;
assign a46866 = a46864 & ~a41710;
assign a46868 = a46866 & a41626;
assign a46870 = ~a46868 & a46862;
assign a46872 = a46214 & ~a42722;
assign a46874 = a46872 & ~a41710;
assign a46876 = a46874 & ~a41626;
assign a46878 = ~a46876 & a46870;
assign a46880 = a46246 & ~a42704;
assign a46882 = ~a46880 & a46878;
assign a46884 = ~a42678 & a41718;
assign a46886 = a46884 & l2318;
assign a46888 = a46886 & a41720;
assign a46890 = ~a46888 & a46882;
assign a46892 = a46300 & ~a42654;
assign a46894 = a46892 & a41712;
assign a46896 = ~a46894 & a46890;
assign a46898 = a46300 & ~a42628;
assign a46900 = a46898 & ~a41626;
assign a46902 = a46900 & ~a41710;
assign a46904 = ~a46902 & a46896;
assign a46906 = a46356 & ~a42604;
assign a46908 = a46906 & a41626;
assign a46910 = ~a46908 & a46904;
assign a46912 = a46356 & ~a42580;
assign a46914 = a46912 & ~a41626;
assign a46916 = ~a46914 & a46910;
assign a46918 = ~a46916 & a46168;
assign a46920 = a46864 & a41720;
assign a46922 = a46196 & ~a42758;
assign a46924 = ~a46922 & ~a46920;
assign a46926 = a46874 & a41626;
assign a46928 = ~a46926 & a46924;
assign a46930 = ~a42704 & a41718;
assign a46932 = a46930 & a46414;
assign a46934 = a46932 & ~a41626;
assign a46936 = ~a46934 & a46928;
assign a46938 = a46246 & ~a42678;
assign a46940 = ~a46938 & a46936;
assign a46942 = a46892 & ~a41626;
assign a46944 = a46942 & a41710;
assign a46946 = ~a46944 & a46940;
assign a46948 = a46898 & a41712;
assign a46950 = ~a46948 & a46946;
assign a46952 = a46440 & ~a42604;
assign a46954 = a46952 & ~a41626;
assign a46956 = ~a46954 & a46950;
assign a46958 = a46912 & a41626;
assign a46960 = ~a46958 & a46956;
assign a46962 = ~a42554 & ~l2318;
assign a46964 = a46962 & ~a41718;
assign a46966 = a46964 & ~a41626;
assign a46968 = ~a46966 & a46960;
assign a46970 = ~a46968 & ~a46166;
assign a46972 = ~a46970 & ~a46918;
assign a46974 = a46962 & a41722;
assign a46976 = a46196 & ~a42580;
assign a46978 = ~a46976 & ~a46974;
assign a46980 = a46854 & a46470;
assign a46982 = ~a46980 & a46978;
assign a46984 = a46866 & ~a41626;
assign a46986 = ~a46984 & a46982;
assign a46988 = a46246 & ~a42722;
assign a46990 = ~a46988 & a46986;
assign a46992 = a46930 & a46486;
assign a46994 = ~a46992 & a46990;
assign a46996 = a46886 & a41712;
assign a46998 = ~a46996 & a46994;
assign a47000 = a46942 & ~a41710;
assign a47002 = ~a47000 & a46998;
assign a47004 = a46500 & ~a42628;
assign a47006 = ~a47004 & a47002;
assign a47008 = a46906 & ~a41626;
assign a47010 = ~a47008 & a47006;
assign a47012 = ~a47010 & a45946;
assign a47014 = ~a47012 & a46972;
assign a47016 = ~a47014 & i812;
assign a47018 = ~a47016 & ~a46852;
assign a47020 = a47014 & ~i812;
assign a47022 = ~a47020 & ~a47018;
assign a47024 = ~a43056 & ~l2318;
assign a47026 = a47024 & ~a41626;
assign a47028 = a47026 & a46178;
assign a47030 = a46196 & ~a42852;
assign a47032 = ~a47030 & ~a47028;
assign a47034 = a46214 & ~a43038;
assign a47036 = a47034 & ~a41710;
assign a47038 = a47036 & a41626;
assign a47040 = ~a47038 & a47032;
assign a47042 = a46214 & ~a43020;
assign a47044 = a47042 & ~a41710;
assign a47046 = a47044 & ~a41626;
assign a47048 = ~a47046 & a47040;
assign a47050 = a46246 & ~a43002;
assign a47052 = ~a47050 & a47048;
assign a47054 = ~a42976 & a41718;
assign a47056 = a47054 & l2318;
assign a47058 = a47056 & a41720;
assign a47060 = ~a47058 & a47052;
assign a47062 = a46300 & ~a42952;
assign a47064 = a47062 & a41712;
assign a47066 = ~a47064 & a47060;
assign a47068 = a46300 & ~a42926;
assign a47070 = a47068 & ~a41626;
assign a47072 = a47070 & ~a41710;
assign a47074 = ~a47072 & a47066;
assign a47076 = a46356 & ~a42902;
assign a47078 = a47076 & a41626;
assign a47080 = ~a47078 & a47074;
assign a47082 = a46356 & ~a42878;
assign a47084 = a47082 & ~a41626;
assign a47086 = ~a47084 & a47080;
assign a47088 = ~a47086 & a46168;
assign a47090 = a47034 & a41720;
assign a47092 = a46196 & ~a43056;
assign a47094 = ~a47092 & ~a47090;
assign a47096 = a47044 & a41626;
assign a47098 = ~a47096 & a47094;
assign a47100 = ~a43002 & a41718;
assign a47102 = a47100 & a46414;
assign a47104 = a47102 & ~a41626;
assign a47106 = ~a47104 & a47098;
assign a47108 = a46246 & ~a42976;
assign a47110 = ~a47108 & a47106;
assign a47112 = a47062 & ~a41626;
assign a47114 = a47112 & a41710;
assign a47116 = ~a47114 & a47110;
assign a47118 = a47068 & a41712;
assign a47120 = ~a47118 & a47116;
assign a47122 = a46440 & ~a42902;
assign a47124 = a47122 & ~a41626;
assign a47126 = ~a47124 & a47120;
assign a47128 = a47082 & a41626;
assign a47130 = ~a47128 & a47126;
assign a47132 = ~a42852 & ~l2318;
assign a47134 = a47132 & ~a41718;
assign a47136 = a47134 & ~a41626;
assign a47138 = ~a47136 & a47130;
assign a47140 = ~a47138 & ~a46166;
assign a47142 = ~a47140 & ~a47088;
assign a47144 = a47132 & a41722;
assign a47146 = a46196 & ~a42878;
assign a47148 = ~a47146 & ~a47144;
assign a47150 = a47024 & a46470;
assign a47152 = ~a47150 & a47148;
assign a47154 = a47036 & ~a41626;
assign a47156 = ~a47154 & a47152;
assign a47158 = a46246 & ~a43020;
assign a47160 = ~a47158 & a47156;
assign a47162 = a47100 & a46486;
assign a47164 = ~a47162 & a47160;
assign a47166 = a47056 & a41712;
assign a47168 = ~a47166 & a47164;
assign a47170 = a47112 & ~a41710;
assign a47172 = ~a47170 & a47168;
assign a47174 = a46500 & ~a42926;
assign a47176 = ~a47174 & a47172;
assign a47178 = a47076 & ~a41626;
assign a47180 = ~a47178 & a47176;
assign a47182 = ~a47180 & a45946;
assign a47184 = ~a47182 & a47142;
assign a47186 = ~a47184 & i814;
assign a47188 = ~a47186 & ~a47022;
assign a47190 = a47184 & ~i814;
assign a47192 = ~a47190 & ~a47188;
assign a47194 = ~a43354 & ~l2318;
assign a47196 = a47194 & ~a41626;
assign a47198 = a47196 & a46178;
assign a47200 = a46196 & ~a43150;
assign a47202 = ~a47200 & ~a47198;
assign a47204 = a46214 & ~a43336;
assign a47206 = a47204 & ~a41710;
assign a47208 = a47206 & a41626;
assign a47210 = ~a47208 & a47202;
assign a47212 = a46214 & ~a43318;
assign a47214 = a47212 & ~a41710;
assign a47216 = a47214 & ~a41626;
assign a47218 = ~a47216 & a47210;
assign a47220 = a46246 & ~a43300;
assign a47222 = ~a47220 & a47218;
assign a47224 = ~a43274 & a41718;
assign a47226 = a47224 & l2318;
assign a47228 = a47226 & a41720;
assign a47230 = ~a47228 & a47222;
assign a47232 = a46300 & ~a43250;
assign a47234 = a47232 & a41712;
assign a47236 = ~a47234 & a47230;
assign a47238 = a46300 & ~a43224;
assign a47240 = a47238 & ~a41626;
assign a47242 = a47240 & ~a41710;
assign a47244 = ~a47242 & a47236;
assign a47246 = a46356 & ~a43200;
assign a47248 = a47246 & a41626;
assign a47250 = ~a47248 & a47244;
assign a47252 = a46356 & ~a43176;
assign a47254 = a47252 & ~a41626;
assign a47256 = ~a47254 & a47250;
assign a47258 = ~a47256 & a46168;
assign a47260 = a47204 & a41720;
assign a47262 = a46196 & ~a43354;
assign a47264 = ~a47262 & ~a47260;
assign a47266 = a47214 & a41626;
assign a47268 = ~a47266 & a47264;
assign a47270 = ~a43300 & a41718;
assign a47272 = a47270 & a46414;
assign a47274 = a47272 & ~a41626;
assign a47276 = ~a47274 & a47268;
assign a47278 = a46246 & ~a43274;
assign a47280 = ~a47278 & a47276;
assign a47282 = a47232 & ~a41626;
assign a47284 = a47282 & a41710;
assign a47286 = ~a47284 & a47280;
assign a47288 = a47238 & a41712;
assign a47290 = ~a47288 & a47286;
assign a47292 = a46440 & ~a43200;
assign a47294 = a47292 & ~a41626;
assign a47296 = ~a47294 & a47290;
assign a47298 = a47252 & a41626;
assign a47300 = ~a47298 & a47296;
assign a47302 = ~a43150 & ~l2318;
assign a47304 = a47302 & ~a41718;
assign a47306 = a47304 & ~a41626;
assign a47308 = ~a47306 & a47300;
assign a47310 = ~a47308 & ~a46166;
assign a47312 = ~a47310 & ~a47258;
assign a47314 = a47302 & a41722;
assign a47316 = a46196 & ~a43176;
assign a47318 = ~a47316 & ~a47314;
assign a47320 = a47194 & a46470;
assign a47322 = ~a47320 & a47318;
assign a47324 = a47206 & ~a41626;
assign a47326 = ~a47324 & a47322;
assign a47328 = a46246 & ~a43318;
assign a47330 = ~a47328 & a47326;
assign a47332 = a47270 & a46486;
assign a47334 = ~a47332 & a47330;
assign a47336 = a47226 & a41712;
assign a47338 = ~a47336 & a47334;
assign a47340 = a47282 & ~a41710;
assign a47342 = ~a47340 & a47338;
assign a47344 = a46500 & ~a43224;
assign a47346 = ~a47344 & a47342;
assign a47348 = a47246 & ~a41626;
assign a47350 = ~a47348 & a47346;
assign a47352 = ~a47350 & a45946;
assign a47354 = ~a47352 & a47312;
assign a47356 = ~a47354 & i816;
assign a47358 = ~a47356 & ~a47192;
assign a47360 = a47354 & ~i816;
assign a47362 = ~a47360 & ~a47358;
assign a47364 = ~a43650 & ~l2318;
assign a47366 = a47364 & ~a41626;
assign a47368 = a47366 & a46178;
assign a47370 = a46196 & ~a43446;
assign a47372 = ~a47370 & ~a47368;
assign a47374 = a46214 & ~a43632;
assign a47376 = a47374 & ~a41710;
assign a47378 = a47376 & a41626;
assign a47380 = ~a47378 & a47372;
assign a47382 = a46214 & ~a43614;
assign a47384 = a47382 & ~a41710;
assign a47386 = a47384 & ~a41626;
assign a47388 = ~a47386 & a47380;
assign a47390 = a46246 & ~a43596;
assign a47392 = ~a47390 & a47388;
assign a47394 = ~a43570 & a41718;
assign a47396 = a47394 & l2318;
assign a47398 = a47396 & a41720;
assign a47400 = ~a47398 & a47392;
assign a47402 = a46300 & ~a43546;
assign a47404 = a47402 & a41712;
assign a47406 = ~a47404 & a47400;
assign a47408 = a46300 & ~a43520;
assign a47410 = a47408 & ~a41626;
assign a47412 = a47410 & ~a41710;
assign a47414 = ~a47412 & a47406;
assign a47416 = a46356 & ~a43496;
assign a47418 = a47416 & a41626;
assign a47420 = ~a47418 & a47414;
assign a47422 = a46356 & ~a43472;
assign a47424 = a47422 & ~a41626;
assign a47426 = ~a47424 & a47420;
assign a47428 = ~a47426 & a46168;
assign a47430 = a47374 & a41720;
assign a47432 = a46196 & ~a43650;
assign a47434 = ~a47432 & ~a47430;
assign a47436 = a47384 & a41626;
assign a47438 = ~a47436 & a47434;
assign a47440 = ~a43596 & a41718;
assign a47442 = a47440 & a46414;
assign a47444 = a47442 & ~a41626;
assign a47446 = ~a47444 & a47438;
assign a47448 = a46246 & ~a43570;
assign a47450 = ~a47448 & a47446;
assign a47452 = a47402 & ~a41626;
assign a47454 = a47452 & a41710;
assign a47456 = ~a47454 & a47450;
assign a47458 = a47408 & a41712;
assign a47460 = ~a47458 & a47456;
assign a47462 = a46440 & ~a43496;
assign a47464 = a47462 & ~a41626;
assign a47466 = ~a47464 & a47460;
assign a47468 = a47422 & a41626;
assign a47470 = ~a47468 & a47466;
assign a47472 = ~a43446 & ~l2318;
assign a47474 = a47472 & ~a41718;
assign a47476 = a47474 & ~a41626;
assign a47478 = ~a47476 & a47470;
assign a47480 = ~a47478 & ~a46166;
assign a47482 = ~a47480 & ~a47428;
assign a47484 = a47472 & a41722;
assign a47486 = a46196 & ~a43472;
assign a47488 = ~a47486 & ~a47484;
assign a47490 = a47364 & a46470;
assign a47492 = ~a47490 & a47488;
assign a47494 = a47376 & ~a41626;
assign a47496 = ~a47494 & a47492;
assign a47498 = a46246 & ~a43614;
assign a47500 = ~a47498 & a47496;
assign a47502 = a47440 & a46486;
assign a47504 = ~a47502 & a47500;
assign a47506 = a47396 & a41712;
assign a47508 = ~a47506 & a47504;
assign a47510 = a47452 & ~a41710;
assign a47512 = ~a47510 & a47508;
assign a47514 = a46500 & ~a43520;
assign a47516 = ~a47514 & a47512;
assign a47518 = a47416 & ~a41626;
assign a47520 = ~a47518 & a47516;
assign a47522 = ~a47520 & a45946;
assign a47524 = ~a47522 & a47482;
assign a47526 = ~a47524 & i818;
assign a47528 = ~a47526 & ~a47362;
assign a47530 = a47524 & ~i818;
assign a47532 = ~a47530 & ~a47528;
assign a47534 = ~l2322 & l890;
assign a47536 = ~a45452 & ~l890;
assign a47538 = ~a47536 & ~a47534;
assign a47540 = ~a47538 & ~l2318;
assign a47542 = a47540 & ~a41626;
assign a47544 = a47542 & a46178;
assign a47546 = ~l2324 & l890;
assign a47548 = ~a45846 & ~a41868;
assign a47550 = a41868 & i822;
assign a47552 = ~a47550 & ~a47548;
assign a47554 = ~a47552 & ~l890;
assign a47556 = ~a47554 & ~a47546;
assign a47558 = ~a47556 & a46196;
assign a47560 = ~a47558 & ~a47544;
assign a47562 = ~l2326 & l890;
assign a47564 = ~a45444 & ~l890;
assign a47566 = ~a47564 & ~a47562;
assign a47568 = ~a47566 & a46214;
assign a47570 = a47568 & ~a41710;
assign a47572 = a47570 & a41626;
assign a47574 = ~a47572 & a47560;
assign a47576 = ~l2328 & l890;
assign a47578 = ~a45464 & ~l890;
assign a47580 = ~a47578 & ~a47576;
assign a47582 = ~a47580 & a46214;
assign a47584 = a47582 & ~a41710;
assign a47586 = a47584 & ~a41626;
assign a47588 = ~a47586 & a47574;
assign a47590 = ~l2330 & l890;
assign a47592 = a42074 & i638;
assign a47594 = a47592 & ~a42078;
assign a47596 = a42078 & i714;
assign a47598 = ~a47596 & ~a47594;
assign a47600 = ~a47598 & ~a42086;
assign a47602 = a42086 & i822;
assign a47604 = ~a47602 & ~a47600;
assign a47606 = ~a47604 & ~l890;
assign a47608 = ~a47606 & ~a47590;
assign a47610 = ~a47608 & a46246;
assign a47612 = ~a47610 & a47588;
assign a47614 = ~l2332 & l890;
assign a47616 = a42038 & i638;
assign a47618 = a47616 & ~a42042;
assign a47620 = a42042 & i714;
assign a47622 = ~a47620 & ~a47618;
assign a47624 = ~a47622 & ~a42052;
assign a47626 = a42052 & i822;
assign a47628 = ~a47626 & ~a47624;
assign a47630 = ~a47628 & ~l890;
assign a47632 = ~a47630 & ~a47614;
assign a47634 = ~a47632 & a41718;
assign a47636 = a47634 & l2318;
assign a47638 = a47636 & a41720;
assign a47640 = ~a47638 & a47612;
assign a47642 = ~l2334 & l890;
assign a47644 = a42006 & i638;
assign a47646 = a47644 & ~a42010;
assign a47648 = a42010 & i714;
assign a47650 = ~a47648 & ~a47646;
assign a47652 = ~a47650 & ~a42020;
assign a47654 = a42020 & i822;
assign a47656 = ~a47654 & ~a47652;
assign a47658 = ~a47656 & ~l890;
assign a47660 = ~a47658 & ~a47642;
assign a47662 = ~a47660 & a46300;
assign a47664 = a47662 & a41712;
assign a47666 = ~a47664 & a47640;
assign a47668 = ~l2336 & l890;
assign a47670 = a41970 & i638;
assign a47672 = a47670 & ~a41974;
assign a47674 = a41974 & i714;
assign a47676 = ~a47674 & ~a47672;
assign a47678 = ~a47676 & ~a41986;
assign a47680 = a41986 & i822;
assign a47682 = ~a47680 & ~a47678;
assign a47684 = ~a47682 & ~l890;
assign a47686 = ~a47684 & ~a47668;
assign a47688 = ~a47686 & a46300;
assign a47690 = a47688 & ~a41626;
assign a47692 = a47690 & ~a41710;
assign a47694 = ~a47692 & a47666;
assign a47696 = ~l2338 & l890;
assign a47698 = a41936 & i638;
assign a47700 = a47698 & ~a41940;
assign a47702 = a41940 & i714;
assign a47704 = ~a47702 & ~a47700;
assign a47706 = ~a47704 & ~a41948;
assign a47708 = a41948 & i822;
assign a47710 = ~a47708 & ~a47706;
assign a47712 = ~a47710 & ~l890;
assign a47714 = ~a47712 & ~a47696;
assign a47716 = ~a47714 & a46356;
assign a47718 = a47716 & a41626;
assign a47720 = ~a47718 & a47694;
assign a47722 = ~l2340 & l890;
assign a47724 = ~a45856 & ~a41916;
assign a47726 = a41916 & i822;
assign a47728 = ~a47726 & ~a47724;
assign a47730 = ~a47728 & ~l890;
assign a47732 = ~a47730 & ~a47722;
assign a47734 = ~a47732 & a46356;
assign a47736 = a47734 & ~a41626;
assign a47738 = ~a47736 & a47720;
assign a47740 = ~a47738 & a46168;
assign a47742 = a47568 & a41720;
assign a47744 = ~a47538 & a46196;
assign a47746 = ~a47744 & ~a47742;
assign a47748 = a47584 & a41626;
assign a47750 = ~a47748 & a47746;
assign a47752 = ~a47608 & a41718;
assign a47754 = a47752 & a46414;
assign a47756 = a47754 & ~a41626;
assign a47758 = ~a47756 & a47750;
assign a47760 = ~a47632 & a46246;
assign a47762 = ~a47760 & a47758;
assign a47764 = a47662 & ~a41626;
assign a47766 = a47764 & a41710;
assign a47768 = ~a47766 & a47762;
assign a47770 = a47688 & a41712;
assign a47772 = ~a47770 & a47768;
assign a47774 = ~a47714 & a46440;
assign a47776 = a47774 & ~a41626;
assign a47778 = ~a47776 & a47772;
assign a47780 = a47734 & a41626;
assign a47782 = ~a47780 & a47778;
assign a47784 = ~a47556 & ~l2318;
assign a47786 = a47784 & ~a41718;
assign a47788 = a47786 & ~a41626;
assign a47790 = ~a47788 & a47782;
assign a47792 = ~a47790 & ~a46166;
assign a47794 = ~a47792 & ~a47740;
assign a47796 = a47784 & a41722;
assign a47798 = ~a47732 & a46196;
assign a47800 = ~a47798 & ~a47796;
assign a47802 = a47540 & a46470;
assign a47804 = ~a47802 & a47800;
assign a47806 = a47570 & ~a41626;
assign a47808 = ~a47806 & a47804;
assign a47810 = ~a47580 & a46246;
assign a47812 = ~a47810 & a47808;
assign a47814 = a47752 & a46486;
assign a47816 = ~a47814 & a47812;
assign a47818 = a47636 & a41712;
assign a47820 = ~a47818 & a47816;
assign a47822 = a47764 & ~a41710;
assign a47824 = ~a47822 & a47820;
assign a47826 = ~a47686 & a46500;
assign a47828 = ~a47826 & a47824;
assign a47830 = a47716 & ~a41626;
assign a47832 = ~a47830 & a47828;
assign a47834 = ~a47832 & a45946;
assign a47836 = ~a47834 & a47794;
assign a47838 = ~a47836 & i820;
assign a47840 = ~a47838 & ~a47532;
assign a47842 = a47836 & ~i820;
assign a47844 = ~a47842 & ~a47840;
assign a47846 = a47844 & a46518;
assign a47848 = a46680 & ~i808;
assign a47850 = ~a47848 & ~a46850;
assign a47852 = ~a47850 & ~a46846;
assign a47854 = ~a47852 & ~a47020;
assign a47856 = ~a47854 & ~a47016;
assign a47858 = ~a47856 & ~a47190;
assign a47860 = ~a47858 & ~a47186;
assign a47862 = ~a47860 & ~a47360;
assign a47864 = ~a47862 & ~a47356;
assign a47866 = ~a47864 & ~a47530;
assign a47868 = ~a47866 & ~a47526;
assign a47870 = ~a47868 & ~a47842;
assign a47872 = ~a47838 & ~a46518;
assign a47874 = a47872 & ~a47870;
assign a47876 = ~a47874 & ~a47846;
assign a47878 = a41722 & ~l2318;
assign a47880 = a47878 & a43738;
assign a47882 = a46196 & a43866;
assign a47884 = ~a47882 & ~a47880;
assign a47886 = a46470 & ~l2318;
assign a47888 = a47886 & a44062;
assign a47890 = ~a47888 & a47884;
assign a47892 = a44038 & a41780;
assign a47894 = ~a47892 & a47890;
assign a47896 = a46246 & a43996;
assign a47898 = ~a47896 & a47894;
assign a47900 = a46484 & a41718;
assign a47902 = a47900 & a43952;
assign a47904 = a47902 & a41710;
assign a47906 = ~a47904 & a47898;
assign a47908 = a46244 & ~a41710;
assign a47910 = a47908 & a44142;
assign a47912 = ~a47910 & a47906;
assign a47914 = a47900 & ~a41710;
assign a47916 = a47914 & a44098;
assign a47918 = ~a47916 & a47912;
assign a47920 = a46500 & a43902;
assign a47922 = ~a47920 & a47918;
assign a47924 = ~a41718 & ~a41626;
assign a47926 = a47924 & ~l2318;
assign a47928 = a47926 & a43840;
assign a47930 = ~a47928 & a47922;
assign a47932 = ~a47930 & ~a46166;
assign a47934 = a47878 & a43866;
assign a47936 = a46196 & a43840;
assign a47938 = ~a47936 & ~a47934;
assign a47940 = a47886 & a43738;
assign a47942 = ~a47940 & a47938;
assign a47944 = a44062 & a41780;
assign a47946 = ~a47944 & a47942;
assign a47948 = a46246 & a44038;
assign a47950 = ~a47948 & a47946;
assign a47952 = a46486 & a43996;
assign a47954 = ~a47952 & a47950;
assign a47956 = a47908 & a43952;
assign a47958 = ~a47956 & a47954;
assign a47960 = a47900 & a44142;
assign a47962 = a47960 & ~a41710;
assign a47964 = ~a47962 & a47958;
assign a47966 = a46500 & a44098;
assign a47968 = ~a47966 & a47964;
assign a47970 = a47926 & a43902;
assign a47972 = ~a47970 & a47968;
assign a47974 = ~a47972 & a46168;
assign a47976 = ~a47974 & ~a47932;
assign a47978 = a47878 & a43840;
assign a47980 = a46196 & a43902;
assign a47982 = ~a47980 & ~a47978;
assign a47984 = a47886 & a43866;
assign a47986 = ~a47984 & a47982;
assign a47988 = a43738 & a41780;
assign a47990 = ~a47988 & a47986;
assign a47992 = a46246 & a44062;
assign a47994 = ~a47992 & a47990;
assign a47996 = a46486 & a44038;
assign a47998 = ~a47996 & a47994;
assign a48000 = a47908 & a43996;
assign a48002 = ~a48000 & a47998;
assign a48004 = a47902 & ~a41710;
assign a48006 = ~a48004 & a48002;
assign a48008 = a46500 & a44142;
assign a48010 = ~a48008 & a48006;
assign a48012 = a47926 & a44098;
assign a48014 = ~a48012 & a48010;
assign a48016 = ~a48014 & a45946;
assign a48018 = ~a48016 & a47976;
assign a48020 = ~a48018 & ~a41644;
assign a48024 = ~a47924 & ~a46196;
assign a48026 = ~a48024 & a45946;
assign a48028 = a46168 & ~a41718;
assign a48030 = ~a46166 & ~a41834;
assign a48032 = ~a48030 & ~a48028;
assign a48036 = ~a46246 & ~a41778;
assign a48038 = a48036 & ~a41830;
assign a48040 = ~a48038 & a45946;
assign a48042 = a46168 & ~a41710;
assign a48044 = ~a46166 & ~a41724;
assign a48046 = ~a48044 & ~a48042;
assign a48050 = ~a46484 & ~a46438;
assign a48052 = a48050 & ~a41830;
assign a48054 = ~a48052 & a45946;
assign a48056 = a46168 & l2318;
assign a48058 = ~a46166 & ~a41788;
assign a48060 = ~a48058 & ~a48056;
assign a48062 = a48060 & ~a48054;
assign a48064 = ~a46582 & a45946;
assign a48066 = ~a46634 & a46168;
assign a48068 = a46538 & a41720;
assign a48070 = a46196 & ~a42138;
assign a48072 = ~a48070 & ~a48068;
assign a48074 = a46598 & a41626;
assign a48076 = ~a48074 & a48072;
assign a48078 = a46550 & a41780;
assign a48080 = ~a48078 & a48076;
assign a48082 = a46246 & ~a42030;
assign a48084 = ~a48082 & a48080;
assign a48086 = a46566 & a41710;
assign a48088 = ~a48086 & a48084;
assign a48090 = a46618 & a41626;
assign a48092 = ~a48090 & a48088;
assign a48094 = a47914 & ~a41926;
assign a48096 = ~a48094 & a48092;
assign a48098 = a46630 & a41626;
assign a48100 = ~a48098 & a48096;
assign a48102 = a46522 & ~a41718;
assign a48104 = ~a48102 & a48100;
assign a48106 = ~a48104 & ~a46166;
assign a48108 = ~a48106 & ~a48066;
assign a48110 = a48108 & ~a48064;
assign a48112 = a48110 & ~i808;
assign a48114 = ~a46746 & a45946;
assign a48116 = ~a46798 & a46168;
assign a48118 = a46702 & a41720;
assign a48120 = a46196 & ~a42442;
assign a48122 = ~a48120 & ~a48118;
assign a48124 = a46762 & a41626;
assign a48126 = ~a48124 & a48122;
assign a48128 = a46714 & a41780;
assign a48130 = ~a48128 & a48126;
assign a48132 = a46246 & ~a42356;
assign a48134 = ~a48132 & a48130;
assign a48136 = a46730 & a41710;
assign a48138 = ~a48136 & a48134;
assign a48140 = a46782 & a41626;
assign a48142 = ~a48140 & a48138;
assign a48144 = a47914 & ~a42282;
assign a48146 = ~a48144 & a48142;
assign a48148 = a46794 & a41626;
assign a48150 = ~a48148 & a48146;
assign a48152 = a46686 & ~a41718;
assign a48154 = ~a48152 & a48150;
assign a48156 = ~a48154 & ~a46166;
assign a48158 = ~a48156 & ~a48116;
assign a48160 = a48158 & ~a48114;
assign a48162 = a48160 & ~i810;
assign a48164 = ~a48162 & ~a48112;
assign a48166 = ~a48160 & i810;
assign a48168 = ~a48166 & ~a48164;
assign a48170 = ~a46916 & a45946;
assign a48172 = ~a46968 & a46168;
assign a48174 = a46872 & a41720;
assign a48176 = a46196 & ~a42740;
assign a48178 = ~a48176 & ~a48174;
assign a48180 = a46932 & a41626;
assign a48182 = ~a48180 & a48178;
assign a48184 = a46884 & a41780;
assign a48186 = ~a48184 & a48182;
assign a48188 = a46246 & ~a42654;
assign a48190 = ~a48188 & a48186;
assign a48192 = a46900 & a41710;
assign a48194 = ~a48192 & a48190;
assign a48196 = a46952 & a41626;
assign a48198 = ~a48196 & a48194;
assign a48200 = a47914 & ~a42580;
assign a48202 = ~a48200 & a48198;
assign a48204 = a46964 & a41626;
assign a48206 = ~a48204 & a48202;
assign a48208 = a46856 & ~a41718;
assign a48210 = ~a48208 & a48206;
assign a48212 = ~a48210 & ~a46166;
assign a48214 = ~a48212 & ~a48172;
assign a48216 = a48214 & ~a48170;
assign a48218 = a48216 & ~i812;
assign a48220 = ~a48218 & ~a48168;
assign a48222 = ~a48216 & i812;
assign a48224 = ~a48222 & ~a48220;
assign a48226 = ~a47086 & a45946;
assign a48228 = ~a47138 & a46168;
assign a48230 = a47042 & a41720;
assign a48232 = a46196 & ~a43038;
assign a48234 = ~a48232 & ~a48230;
assign a48236 = a47102 & a41626;
assign a48238 = ~a48236 & a48234;
assign a48240 = a47054 & a41780;
assign a48242 = ~a48240 & a48238;
assign a48244 = a46246 & ~a42952;
assign a48246 = ~a48244 & a48242;
assign a48248 = a47070 & a41710;
assign a48250 = ~a48248 & a48246;
assign a48252 = a47122 & a41626;
assign a48254 = ~a48252 & a48250;
assign a48256 = a47914 & ~a42878;
assign a48258 = ~a48256 & a48254;
assign a48260 = a47134 & a41626;
assign a48262 = ~a48260 & a48258;
assign a48264 = a47026 & ~a41718;
assign a48266 = ~a48264 & a48262;
assign a48268 = ~a48266 & ~a46166;
assign a48270 = ~a48268 & ~a48228;
assign a48272 = a48270 & ~a48226;
assign a48274 = a48272 & ~i814;
assign a48276 = ~a48274 & ~a48224;
assign a48278 = ~a48272 & i814;
assign a48280 = ~a48278 & ~a48276;
assign a48282 = ~a47256 & a45946;
assign a48284 = ~a47308 & a46168;
assign a48286 = a47212 & a41720;
assign a48288 = a46196 & ~a43336;
assign a48290 = ~a48288 & ~a48286;
assign a48292 = a47272 & a41626;
assign a48294 = ~a48292 & a48290;
assign a48296 = a47224 & a41780;
assign a48298 = ~a48296 & a48294;
assign a48300 = a46246 & ~a43250;
assign a48302 = ~a48300 & a48298;
assign a48304 = a47240 & a41710;
assign a48306 = ~a48304 & a48302;
assign a48308 = a47292 & a41626;
assign a48310 = ~a48308 & a48306;
assign a48312 = a47914 & ~a43176;
assign a48314 = ~a48312 & a48310;
assign a48316 = a47304 & a41626;
assign a48318 = ~a48316 & a48314;
assign a48320 = a47196 & ~a41718;
assign a48322 = ~a48320 & a48318;
assign a48324 = ~a48322 & ~a46166;
assign a48326 = ~a48324 & ~a48284;
assign a48328 = a48326 & ~a48282;
assign a48330 = a48328 & ~i816;
assign a48332 = ~a48330 & ~a48280;
assign a48334 = ~a48328 & i816;
assign a48336 = ~a48334 & ~a48332;
assign a48338 = ~a47426 & a45946;
assign a48340 = ~a47478 & a46168;
assign a48342 = a47382 & a41720;
assign a48344 = a46196 & ~a43632;
assign a48346 = ~a48344 & ~a48342;
assign a48348 = a47442 & a41626;
assign a48350 = ~a48348 & a48346;
assign a48352 = a47394 & a41780;
assign a48354 = ~a48352 & a48350;
assign a48356 = a46246 & ~a43546;
assign a48358 = ~a48356 & a48354;
assign a48360 = a47410 & a41710;
assign a48362 = ~a48360 & a48358;
assign a48364 = a47462 & a41626;
assign a48366 = ~a48364 & a48362;
assign a48368 = a47914 & ~a43472;
assign a48370 = ~a48368 & a48366;
assign a48372 = a47474 & a41626;
assign a48374 = ~a48372 & a48370;
assign a48376 = a47366 & ~a41718;
assign a48378 = ~a48376 & a48374;
assign a48380 = ~a48378 & ~a46166;
assign a48382 = ~a48380 & ~a48340;
assign a48384 = a48382 & ~a48338;
assign a48386 = a48384 & ~i818;
assign a48388 = ~a48386 & ~a48336;
assign a48390 = ~a48384 & i818;
assign a48392 = ~a48390 & ~a48388;
assign a48394 = ~a47738 & a45946;
assign a48396 = ~a47790 & a46168;
assign a48398 = a47582 & a41720;
assign a48400 = ~a47566 & a46196;
assign a48402 = ~a48400 & ~a48398;
assign a48404 = a47754 & a41626;
assign a48406 = ~a48404 & a48402;
assign a48408 = a47634 & a41780;
assign a48410 = ~a48408 & a48406;
assign a48412 = ~a47660 & a46246;
assign a48414 = ~a48412 & a48410;
assign a48416 = a47690 & a41710;
assign a48418 = ~a48416 & a48414;
assign a48420 = a47774 & a41626;
assign a48422 = ~a48420 & a48418;
assign a48424 = a47914 & ~a47732;
assign a48426 = ~a48424 & a48422;
assign a48428 = a47786 & a41626;
assign a48430 = ~a48428 & a48426;
assign a48432 = a47542 & ~a41718;
assign a48434 = ~a48432 & a48430;
assign a48436 = ~a48434 & ~a46166;
assign a48438 = ~a48436 & ~a48396;
assign a48440 = a48438 & ~a48394;
assign a48442 = a48440 & ~i820;
assign a48444 = ~a48442 & ~a48392;
assign a48446 = ~a48440 & i820;
assign a48448 = ~a46400 & a45946;
assign a48450 = ~a46458 & a46168;
assign a48452 = a46236 & a41720;
assign a48454 = ~a46220 & a46196;
assign a48456 = ~a48454 & ~a48452;
assign a48458 = a46418 & a41626;
assign a48460 = ~a48458 & a48456;
assign a48462 = a46292 & a41780;
assign a48464 = ~a48462 & a48460;
assign a48466 = ~a46320 & a46246;
assign a48468 = ~a48466 & a48464;
assign a48470 = a46350 & a41710;
assign a48472 = ~a48470 & a48468;
assign a48474 = a46442 & a41626;
assign a48476 = ~a48474 & a48472;
assign a48478 = a47914 & ~a46394;
assign a48480 = ~a48478 & a48476;
assign a48482 = a46454 & a41626;
assign a48484 = ~a48482 & a48480;
assign a48486 = a46188 & ~a41718;
assign a48488 = ~a48486 & a48484;
assign a48490 = ~a48488 & ~a46166;
assign a48492 = ~a48490 & ~a48450;
assign a48494 = a48492 & ~a48448;
assign a48496 = a48494 & ~i806;
assign a48498 = ~a48494 & i806;
assign a48500 = ~a48498 & ~a48496;
assign a48502 = ~a48500 & ~a48446;
assign a48504 = a48502 & ~a48444;
assign a48506 = ~a48110 & i808;
assign a48508 = ~a48506 & ~a48166;
assign a48510 = ~a48508 & ~a48162;
assign a48512 = ~a48510 & ~a48222;
assign a48514 = ~a48512 & ~a48218;
assign a48516 = ~a48514 & ~a48278;
assign a48518 = ~a48516 & ~a48274;
assign a48520 = ~a48518 & ~a48334;
assign a48522 = ~a48520 & ~a48330;
assign a48524 = ~a48522 & ~a48390;
assign a48526 = ~a48524 & ~a48386;
assign a48528 = ~a48526 & ~a48446;
assign a48530 = ~a48528 & ~a48442;
assign a48532 = a48530 & a48500;
assign a48534 = ~a47972 & a45946;
assign a48536 = a47926 & a43866;
assign a48538 = a46500 & a43840;
assign a48540 = a47914 & a43902;
assign a48542 = a47908 & a44098;
assign a48544 = a47960 & a41710;
assign a48546 = a46246 & a43952;
assign a48548 = a43996 & a41780;
assign a48550 = a47886 & a44038;
assign a48552 = a47878 & a44062;
assign a48554 = a46196 & a43738;
assign a48556 = ~a48554 & ~a48552;
assign a48558 = a48556 & ~a48550;
assign a48560 = a48558 & ~a48548;
assign a48562 = a48560 & ~a48546;
assign a48564 = a48562 & ~a48544;
assign a48566 = a48564 & ~a48542;
assign a48568 = a48566 & ~a48540;
assign a48570 = a48568 & ~a48538;
assign a48572 = a48570 & ~a48536;
assign a48574 = ~a48572 & ~a46166;
assign a48576 = ~a47930 & a46168;
assign a48578 = ~a48576 & ~a48574;
assign a48580 = a48578 & ~a48534;
assign a48582 = ~a48580 & ~a48532;
assign a48586 = ~a47538 & ~a44508;
assign a48588 = a44508 & i824;
assign a48592 = ~a47556 & ~a44422;
assign a48594 = a44422 & i824;
assign a48598 = ~a47566 & ~a44500;
assign a48600 = a44500 & i824;
assign a48604 = ~a47580 & ~a44492;
assign a48606 = a44492 & i824;
assign a48610 = ~a47608 & ~a44484;
assign a48612 = a44484 & i824;
assign a48616 = ~a47632 & ~a44476;
assign a48618 = a44476 & i824;
assign a48622 = ~a47660 & ~a44466;
assign a48624 = a44466 & i824;
assign a48628 = ~a47686 & ~a44456;
assign a48630 = a44456 & i824;
assign a48634 = ~a47714 & ~a44444;
assign a48636 = a44444 & i824;
assign a48640 = ~a47732 & ~a44436;
assign a48642 = a44436 & i824;
assign a48646 = ~a46184 & ~a44508;
assign a48648 = a44508 & i828;
assign a48652 = ~a46208 & ~a44422;
assign a48654 = a44422 & i828;
assign a48658 = ~a46220 & ~a44500;
assign a48660 = a44500 & i828;
assign a48664 = ~a46234 & ~a44492;
assign a48666 = a44492 & i828;
assign a48670 = ~a46266 & ~a44484;
assign a48672 = a44484 & i828;
assign a48676 = ~a46290 & ~a44476;
assign a48678 = a44476 & i828;
assign a48682 = ~a46320 & ~a44466;
assign a48684 = a44466 & i828;
assign a48688 = ~a46346 & ~a44456;
assign a48690 = a44456 & i828;
assign a48694 = ~a46376 & ~a44444;
assign a48696 = a44444 & i828;
assign a48700 = ~a46394 & ~a44436;
assign a48702 = a44436 & i828;
assign a48706 = ~a44508 & ~a43866;
assign a48708 = ~l2364 & l890;
assign a48710 = a41004 & ~a40726;
assign a48712 = a48710 & a41020;
assign a48714 = ~a48712 & a44824;
assign a48716 = ~a48714 & i670;
assign a48718 = a45216 & ~a44964;
assign a48720 = ~a48718 & ~a48716;
assign a48722 = a48720 & ~i648;
assign a48724 = ~a48722 & ~l890;
assign a48726 = ~a48724 & ~a48708;
assign a48730 = ~a44898 & ~a41742;
assign a48732 = ~a44898 & ~a41678;
assign a48734 = ~a44898 & a41806;
assign a48736 = a48734 & ~a41660;
assign a48738 = a44870 & ~a41678;
assign a48740 = a48738 & a44854;
assign a48742 = a48740 & a41742;
assign a48744 = a44932 & a44870;
assign a48746 = a44922 & a41806;
assign a48748 = a48746 & ~a41660;
assign a48750 = a44856 & a41742;
assign a48752 = a48750 & a41806;
assign a48754 = a48752 & ~a41660;
assign a48756 = a44870 & ~a41660;
assign a48758 = a48756 & a41742;
assign a48760 = a48758 & a41806;
assign a48762 = a48760 & a44854;
assign a48764 = ~a48762 & ~a48754;
assign a48766 = a48764 & ~a48748;
assign a48768 = a48766 & ~a48744;
assign a48770 = a48768 & ~a48742;
assign a48772 = a48770 & ~a48736;
assign a48774 = a48772 & ~a48732;
assign a48776 = a48774 & ~a48730;
assign a48778 = a48776 & a44928;
assign a48780 = ~a48778 & i674;
assign a48782 = a45244 & ~l2372;
assign a48784 = a45586 & ~a45232;
assign a48786 = a48784 & ~l2370;
assign a48788 = a48786 & a48782;
assign a48790 = ~a48788 & ~a48780;
assign a48794 = ~a41724 & a41644;
assign a48796 = a45612 & ~a45244;
assign a48798 = ~a45244 & a45232;
assign a48800 = a48782 & ~a45232;
assign a48802 = ~a48800 & ~a48798;
assign a48804 = ~a48802 & a45616;
assign a48806 = ~a48804 & ~a48796;
assign a48810 = i808 & i650;
assign a48812 = i846 & ~i650;
assign a48814 = ~a48812 & ~a48810;
assign a48816 = a48782 & ~l2370;
assign a48818 = a48816 & ~a44506;
assign a48820 = a48818 & ~a45232;
assign a48822 = ~a44514 & ~l2370;
assign a48824 = a48782 & a45232;
assign a48826 = a48824 & a48822;
assign a48828 = ~a48826 & ~a48820;
assign a48830 = ~a44498 & ~l2370;
assign a48832 = a48830 & a48798;
assign a48834 = ~a48832 & a48828;
assign a48836 = ~a45244 & ~a45232;
assign a48838 = a48836 & ~l2370;
assign a48840 = a48838 & ~a44490;
assign a48842 = ~a48840 & a48834;
assign a48844 = a45244 & l2370;
assign a48846 = a48844 & a45232;
assign a48848 = a48846 & ~a44482;
assign a48850 = ~a48848 & a48842;
assign a48852 = a48844 & ~a44472;
assign a48854 = a48852 & ~a45232;
assign a48856 = ~a48854 & a48850;
assign a48858 = a45232 & l2370;
assign a48860 = ~a45244 & ~l2372;
assign a48862 = a48860 & a48858;
assign a48864 = a48862 & ~a44462;
assign a48866 = ~a48864 & a48856;
assign a48868 = a48860 & l2370;
assign a48870 = a48868 & ~a44450;
assign a48872 = a48870 & ~a45232;
assign a48874 = ~a48872 & a48866;
assign a48876 = a45232 & l2372;
assign a48878 = a48876 & ~a44442;
assign a48880 = ~a48878 & a48874;
assign a48882 = ~a45232 & l2372;
assign a48884 = a48882 & ~l2370;
assign a48886 = a48884 & ~a44428;
assign a48888 = ~a48886 & a48880;
assign a48890 = ~a48888 & ~a45586;
assign a48892 = a48830 & a48800;
assign a48894 = a48818 & a45232;
assign a48896 = ~a48894 & ~a48892;
assign a48898 = a48798 & ~l2370;
assign a48900 = a48898 & ~a44490;
assign a48902 = ~a48900 & a48896;
assign a48904 = a48838 & ~a44482;
assign a48906 = ~a48904 & a48902;
assign a48908 = a48852 & a45232;
assign a48910 = ~a48908 & a48906;
assign a48912 = a48844 & ~a45232;
assign a48914 = a48912 & ~a44462;
assign a48916 = ~a48914 & a48910;
assign a48918 = a48870 & a45232;
assign a48920 = ~a48918 & a48916;
assign a48922 = a48836 & l2370;
assign a48924 = a48922 & ~l2372;
assign a48926 = a48924 & ~a44442;
assign a48928 = ~a48926 & a48920;
assign a48930 = a48876 & ~a44428;
assign a48932 = ~a48930 & a48928;
assign a48934 = a48882 & a48822;
assign a48936 = ~a48934 & a48932;
assign a48938 = ~a48936 & a45586;
assign a48940 = ~a48938 & ~a48890;
assign a48942 = a48940 & a48814;
assign a48944 = i810 & i650;
assign a48946 = i848 & ~i650;
assign a48948 = ~a48946 & ~a48944;
assign a48950 = a48816 & ~a44568;
assign a48952 = a48950 & ~a45232;
assign a48954 = ~a44574 & ~l2370;
assign a48956 = a48954 & a48824;
assign a48958 = ~a48956 & ~a48952;
assign a48960 = ~a44562 & ~l2370;
assign a48962 = a48960 & a48798;
assign a48964 = ~a48962 & a48958;
assign a48966 = a48838 & ~a44556;
assign a48968 = ~a48966 & a48964;
assign a48970 = a48846 & ~a44550;
assign a48972 = ~a48970 & a48968;
assign a48974 = a48844 & ~a44544;
assign a48976 = a48974 & ~a45232;
assign a48978 = ~a48976 & a48972;
assign a48980 = a48862 & ~a44538;
assign a48982 = ~a48980 & a48978;
assign a48984 = a48868 & ~a44532;
assign a48986 = a48984 & ~a45232;
assign a48988 = ~a48986 & a48982;
assign a48990 = a48876 & ~a44526;
assign a48992 = ~a48990 & a48988;
assign a48994 = a48884 & ~a44520;
assign a48996 = ~a48994 & a48992;
assign a48998 = ~a48996 & ~a45586;
assign a49000 = a48960 & a48800;
assign a49002 = a48950 & a45232;
assign a49004 = ~a49002 & ~a49000;
assign a49006 = a48898 & ~a44556;
assign a49008 = ~a49006 & a49004;
assign a49010 = a48838 & ~a44550;
assign a49012 = ~a49010 & a49008;
assign a49014 = a48974 & a45232;
assign a49016 = ~a49014 & a49012;
assign a49018 = a48912 & ~a44538;
assign a49020 = ~a49018 & a49016;
assign a49022 = a48984 & a45232;
assign a49024 = ~a49022 & a49020;
assign a49026 = a48924 & ~a44526;
assign a49028 = ~a49026 & a49024;
assign a49030 = a48876 & ~a44520;
assign a49032 = ~a49030 & a49028;
assign a49034 = a48954 & a48882;
assign a49036 = ~a49034 & a49032;
assign a49038 = ~a49036 & a45586;
assign a49040 = ~a49038 & ~a48998;
assign a49042 = a49040 & a48948;
assign a49044 = ~a49042 & ~a48942;
assign a49046 = ~a49040 & ~a48948;
assign a49048 = ~a49046 & ~a49044;
assign a49050 = i812 & i650;
assign a49052 = i850 & ~i650;
assign a49054 = ~a49052 & ~a49050;
assign a49056 = a48816 & ~a44628;
assign a49058 = a49056 & ~a45232;
assign a49060 = ~a44634 & ~l2370;
assign a49062 = a49060 & a48824;
assign a49064 = ~a49062 & ~a49058;
assign a49066 = ~a44622 & ~l2370;
assign a49068 = a49066 & a48798;
assign a49070 = ~a49068 & a49064;
assign a49072 = a48838 & ~a44616;
assign a49074 = ~a49072 & a49070;
assign a49076 = a48846 & ~a44610;
assign a49078 = ~a49076 & a49074;
assign a49080 = a48844 & ~a44604;
assign a49082 = a49080 & ~a45232;
assign a49084 = ~a49082 & a49078;
assign a49086 = a48862 & ~a44598;
assign a49088 = ~a49086 & a49084;
assign a49090 = a48868 & ~a44592;
assign a49092 = a49090 & ~a45232;
assign a49094 = ~a49092 & a49088;
assign a49096 = a48876 & ~a44586;
assign a49098 = ~a49096 & a49094;
assign a49100 = a48884 & ~a44580;
assign a49102 = ~a49100 & a49098;
assign a49104 = ~a49102 & ~a45586;
assign a49106 = a49066 & a48800;
assign a49108 = a49056 & a45232;
assign a49110 = ~a49108 & ~a49106;
assign a49112 = a48898 & ~a44616;
assign a49114 = ~a49112 & a49110;
assign a49116 = a48838 & ~a44610;
assign a49118 = ~a49116 & a49114;
assign a49120 = a49080 & a45232;
assign a49122 = ~a49120 & a49118;
assign a49124 = a48912 & ~a44598;
assign a49126 = ~a49124 & a49122;
assign a49128 = a49090 & a45232;
assign a49130 = ~a49128 & a49126;
assign a49132 = a48924 & ~a44586;
assign a49134 = ~a49132 & a49130;
assign a49136 = a48876 & ~a44580;
assign a49138 = ~a49136 & a49134;
assign a49140 = a49060 & a48882;
assign a49142 = ~a49140 & a49138;
assign a49144 = ~a49142 & a45586;
assign a49146 = ~a49144 & ~a49104;
assign a49148 = a49146 & a49054;
assign a49150 = ~a49148 & ~a49048;
assign a49152 = ~a49146 & ~a49054;
assign a49154 = ~a49152 & ~a49150;
assign a49156 = i814 & i650;
assign a49158 = i852 & ~i650;
assign a49160 = ~a49158 & ~a49156;
assign a49162 = a48816 & ~a44688;
assign a49164 = a49162 & ~a45232;
assign a49166 = ~a44694 & ~l2370;
assign a49168 = a49166 & a48824;
assign a49170 = ~a49168 & ~a49164;
assign a49172 = ~a44682 & ~l2370;
assign a49174 = a49172 & a48798;
assign a49176 = ~a49174 & a49170;
assign a49178 = a48838 & ~a44676;
assign a49180 = ~a49178 & a49176;
assign a49182 = a48846 & ~a44670;
assign a49184 = ~a49182 & a49180;
assign a49186 = a48844 & ~a44664;
assign a49188 = a49186 & ~a45232;
assign a49190 = ~a49188 & a49184;
assign a49192 = a48862 & ~a44658;
assign a49194 = ~a49192 & a49190;
assign a49196 = a48868 & ~a44652;
assign a49198 = a49196 & ~a45232;
assign a49200 = ~a49198 & a49194;
assign a49202 = a48876 & ~a44646;
assign a49204 = ~a49202 & a49200;
assign a49206 = a48884 & ~a44640;
assign a49208 = ~a49206 & a49204;
assign a49210 = ~a49208 & ~a45586;
assign a49212 = a49172 & a48800;
assign a49214 = a49162 & a45232;
assign a49216 = ~a49214 & ~a49212;
assign a49218 = a48898 & ~a44676;
assign a49220 = ~a49218 & a49216;
assign a49222 = a48838 & ~a44670;
assign a49224 = ~a49222 & a49220;
assign a49226 = a49186 & a45232;
assign a49228 = ~a49226 & a49224;
assign a49230 = a48912 & ~a44658;
assign a49232 = ~a49230 & a49228;
assign a49234 = a49196 & a45232;
assign a49236 = ~a49234 & a49232;
assign a49238 = a48924 & ~a44646;
assign a49240 = ~a49238 & a49236;
assign a49242 = a48876 & ~a44640;
assign a49244 = ~a49242 & a49240;
assign a49246 = a49166 & a48882;
assign a49248 = ~a49246 & a49244;
assign a49250 = ~a49248 & a45586;
assign a49252 = ~a49250 & ~a49210;
assign a49254 = a49252 & a49160;
assign a49256 = ~a49254 & ~a49154;
assign a49258 = ~a49252 & ~a49160;
assign a49260 = ~a49258 & ~a49256;
assign a49262 = i816 & i650;
assign a49264 = i854 & ~i650;
assign a49266 = ~a49264 & ~a49262;
assign a49268 = a48816 & ~a44748;
assign a49270 = a49268 & ~a45232;
assign a49272 = ~a44754 & ~l2370;
assign a49274 = a49272 & a48824;
assign a49276 = ~a49274 & ~a49270;
assign a49278 = ~a44742 & ~l2370;
assign a49280 = a49278 & a48798;
assign a49282 = ~a49280 & a49276;
assign a49284 = a48838 & ~a44736;
assign a49286 = ~a49284 & a49282;
assign a49288 = a48846 & ~a44730;
assign a49290 = ~a49288 & a49286;
assign a49292 = a48844 & ~a44724;
assign a49294 = a49292 & ~a45232;
assign a49296 = ~a49294 & a49290;
assign a49298 = a48862 & ~a44718;
assign a49300 = ~a49298 & a49296;
assign a49302 = a48868 & ~a44712;
assign a49304 = a49302 & ~a45232;
assign a49306 = ~a49304 & a49300;
assign a49308 = a48876 & ~a44706;
assign a49310 = ~a49308 & a49306;
assign a49312 = a48884 & ~a44700;
assign a49314 = ~a49312 & a49310;
assign a49316 = ~a49314 & ~a45586;
assign a49318 = a49278 & a48800;
assign a49320 = a49268 & a45232;
assign a49322 = ~a49320 & ~a49318;
assign a49324 = a48898 & ~a44736;
assign a49326 = ~a49324 & a49322;
assign a49328 = a48838 & ~a44730;
assign a49330 = ~a49328 & a49326;
assign a49332 = a49292 & a45232;
assign a49334 = ~a49332 & a49330;
assign a49336 = a48912 & ~a44718;
assign a49338 = ~a49336 & a49334;
assign a49340 = a49302 & a45232;
assign a49342 = ~a49340 & a49338;
assign a49344 = a48924 & ~a44706;
assign a49346 = ~a49344 & a49342;
assign a49348 = a48876 & ~a44700;
assign a49350 = ~a49348 & a49346;
assign a49352 = a49272 & a48882;
assign a49354 = ~a49352 & a49350;
assign a49356 = ~a49354 & a45586;
assign a49358 = ~a49356 & ~a49316;
assign a49360 = a49358 & a49266;
assign a49362 = ~a49360 & ~a49260;
assign a49364 = ~a49358 & ~a49266;
assign a49366 = ~a49364 & ~a49362;
assign a49368 = i818 & i650;
assign a49370 = i856 & ~i650;
assign a49372 = ~a49370 & ~a49368;
assign a49374 = a48816 & ~a44808;
assign a49376 = a49374 & ~a45232;
assign a49378 = ~a44814 & ~l2370;
assign a49380 = a49378 & a48824;
assign a49382 = ~a49380 & ~a49376;
assign a49384 = ~a44802 & ~l2370;
assign a49386 = a49384 & a48798;
assign a49388 = ~a49386 & a49382;
assign a49390 = a48838 & ~a44796;
assign a49392 = ~a49390 & a49388;
assign a49394 = a48846 & ~a44790;
assign a49396 = ~a49394 & a49392;
assign a49398 = a48844 & ~a44784;
assign a49400 = a49398 & ~a45232;
assign a49402 = ~a49400 & a49396;
assign a49404 = a48862 & ~a44778;
assign a49406 = ~a49404 & a49402;
assign a49408 = a48868 & ~a44772;
assign a49410 = a49408 & ~a45232;
assign a49412 = ~a49410 & a49406;
assign a49414 = a48876 & ~a44766;
assign a49416 = ~a49414 & a49412;
assign a49418 = a48884 & ~a44760;
assign a49420 = ~a49418 & a49416;
assign a49422 = ~a49420 & ~a45586;
assign a49424 = a49384 & a48800;
assign a49426 = a49374 & a45232;
assign a49428 = ~a49426 & ~a49424;
assign a49430 = a48898 & ~a44796;
assign a49432 = ~a49430 & a49428;
assign a49434 = a48838 & ~a44790;
assign a49436 = ~a49434 & a49432;
assign a49438 = a49398 & a45232;
assign a49440 = ~a49438 & a49436;
assign a49442 = a48912 & ~a44778;
assign a49444 = ~a49442 & a49440;
assign a49446 = a49408 & a45232;
assign a49448 = ~a49446 & a49444;
assign a49450 = a48924 & ~a44766;
assign a49452 = ~a49450 & a49448;
assign a49454 = a48876 & ~a44760;
assign a49456 = ~a49454 & a49452;
assign a49458 = a49378 & a48882;
assign a49460 = ~a49458 & a49456;
assign a49462 = ~a49460 & a45586;
assign a49464 = ~a49462 & ~a49422;
assign a49466 = a49464 & a49372;
assign a49468 = ~a49466 & ~a49366;
assign a49470 = ~a49464 & ~a49372;
assign a49472 = ~a49470 & ~a49468;
assign a49474 = i820 & i650;
assign a49476 = i858 & ~i650;
assign a49478 = ~a49476 & ~a49474;
assign a49480 = a48816 & ~a48602;
assign a49482 = a49480 & ~a45232;
assign a49484 = ~a48590 & ~l2370;
assign a49486 = a49484 & a48824;
assign a49488 = ~a49486 & ~a49482;
assign a49490 = ~a48608 & ~l2370;
assign a49492 = a49490 & a48798;
assign a49494 = ~a49492 & a49488;
assign a49496 = a48838 & ~a48614;
assign a49498 = ~a49496 & a49494;
assign a49500 = a48846 & ~a48620;
assign a49502 = ~a49500 & a49498;
assign a49504 = a48844 & ~a48626;
assign a49506 = a49504 & ~a45232;
assign a49508 = ~a49506 & a49502;
assign a49510 = a48862 & ~a48632;
assign a49512 = ~a49510 & a49508;
assign a49514 = a48868 & ~a48638;
assign a49516 = a49514 & ~a45232;
assign a49518 = ~a49516 & a49512;
assign a49520 = a48876 & ~a48644;
assign a49522 = ~a49520 & a49518;
assign a49524 = a48884 & ~a48596;
assign a49526 = ~a49524 & a49522;
assign a49528 = ~a49526 & ~a45586;
assign a49530 = a49490 & a48800;
assign a49532 = a49480 & a45232;
assign a49534 = ~a49532 & ~a49530;
assign a49536 = a48898 & ~a48614;
assign a49538 = ~a49536 & a49534;
assign a49540 = a48838 & ~a48620;
assign a49542 = ~a49540 & a49538;
assign a49544 = a49504 & a45232;
assign a49546 = ~a49544 & a49542;
assign a49548 = a48912 & ~a48632;
assign a49550 = ~a49548 & a49546;
assign a49552 = a49514 & a45232;
assign a49554 = ~a49552 & a49550;
assign a49556 = a48924 & ~a48644;
assign a49558 = ~a49556 & a49554;
assign a49560 = a48876 & ~a48596;
assign a49562 = ~a49560 & a49558;
assign a49564 = a49484 & a48882;
assign a49566 = ~a49564 & a49562;
assign a49568 = ~a49566 & a45586;
assign a49570 = ~a49568 & ~a49528;
assign a49572 = a49570 & a49478;
assign a49574 = ~a49572 & ~a49472;
assign a49576 = ~a49570 & ~a49478;
assign a49578 = i806 & i650;
assign a49580 = i860 & ~i650;
assign a49582 = ~a49580 & ~a49578;
assign a49584 = a48816 & ~a48662;
assign a49586 = a49584 & ~a45232;
assign a49588 = ~a48650 & ~l2370;
assign a49590 = a49588 & a48824;
assign a49592 = ~a49590 & ~a49586;
assign a49594 = ~a48668 & ~l2370;
assign a49596 = a49594 & a48798;
assign a49598 = ~a49596 & a49592;
assign a49600 = a48838 & ~a48674;
assign a49602 = ~a49600 & a49598;
assign a49604 = a48846 & ~a48680;
assign a49606 = ~a49604 & a49602;
assign a49608 = a48844 & ~a48686;
assign a49610 = a49608 & ~a45232;
assign a49612 = ~a49610 & a49606;
assign a49614 = a48862 & ~a48692;
assign a49616 = ~a49614 & a49612;
assign a49618 = a48868 & ~a48698;
assign a49620 = a49618 & ~a45232;
assign a49622 = ~a49620 & a49616;
assign a49624 = a48876 & ~a48704;
assign a49626 = ~a49624 & a49622;
assign a49628 = a48884 & ~a48656;
assign a49630 = ~a49628 & a49626;
assign a49632 = ~a49630 & ~a45586;
assign a49634 = a49594 & a48800;
assign a49636 = a49584 & a45232;
assign a49638 = ~a49636 & ~a49634;
assign a49640 = a48898 & ~a48674;
assign a49642 = ~a49640 & a49638;
assign a49644 = a48838 & ~a48680;
assign a49646 = ~a49644 & a49642;
assign a49648 = a49608 & a45232;
assign a49650 = ~a49648 & a49646;
assign a49652 = a48912 & ~a48692;
assign a49654 = ~a49652 & a49650;
assign a49656 = a49618 & a45232;
assign a49658 = ~a49656 & a49654;
assign a49660 = a48924 & ~a48704;
assign a49662 = ~a49660 & a49658;
assign a49664 = a48876 & ~a48656;
assign a49666 = ~a49664 & a49662;
assign a49668 = a49588 & a48882;
assign a49670 = ~a49668 & a49666;
assign a49672 = ~a49670 & a45586;
assign a49674 = ~a49672 & ~a49632;
assign a49676 = a49674 & a49582;
assign a49678 = ~a49674 & ~a49582;
assign a49680 = ~a49678 & ~a49676;
assign a49682 = ~a49680 & ~a49576;
assign a49684 = a49682 & ~a49574;
assign a49686 = ~a48940 & ~a48814;
assign a49688 = ~a49686 & ~a49046;
assign a49690 = ~a49688 & ~a49042;
assign a49692 = ~a49690 & ~a49152;
assign a49694 = ~a49692 & ~a49148;
assign a49696 = ~a49694 & ~a49258;
assign a49698 = ~a49696 & ~a49254;
assign a49700 = ~a49698 & ~a49364;
assign a49702 = ~a49700 & ~a49360;
assign a49704 = ~a49702 & ~a49470;
assign a49706 = ~a49704 & ~a49466;
assign a49708 = ~a49706 & ~a49576;
assign a49710 = ~a49708 & ~a49572;
assign a49712 = a49710 & a49680;
assign a49714 = a48800 & ~l2370;
assign a49716 = a49714 & a44834;
assign a49718 = a48824 & ~l2370;
assign a49720 = a49718 & a48728;
assign a49722 = ~a49720 & ~a49716;
assign a49724 = ~a44492 & ~a44062;
assign a49726 = ~l2376 & l890;
assign a49728 = a44822 & ~a40726;
assign a49730 = ~a49728 & a44820;
assign a49732 = ~a49730 & i670;
assign a49734 = ~a49732 & ~i648;
assign a49736 = ~a49734 & ~l890;
assign a49738 = ~a49736 & ~a49726;
assign a49742 = a49740 & a48898;
assign a49744 = ~a49742 & a49722;
assign a49746 = ~a44484 & ~a44038;
assign a49748 = ~l2380 & l890;
assign a49750 = ~a44820 & i670;
assign a49752 = ~a49750 & ~i648;
assign a49754 = ~a49752 & ~l890;
assign a49756 = ~a49754 & ~a49748;
assign a49760 = a49758 & a48838;
assign a49762 = ~a49760 & a49744;
assign a49764 = ~a44476 & ~a43996;
assign a49766 = ~l2384 & l890;
assign a49768 = ~a41004 & ~a40754;
assign a49770 = ~a49768 & a41020;
assign a49772 = ~a41004 & ~a40726;
assign a49774 = ~a49772 & a49770;
assign a49776 = ~a49774 & i670;
assign a49778 = ~a49776 & ~i648;
assign a49780 = ~a49778 & ~l890;
assign a49782 = ~a49780 & ~a49766;
assign a49786 = a49784 & a48846;
assign a49788 = ~a49786 & a49762;
assign a49790 = ~l2386 & l890;
assign a49792 = ~a49770 & i670;
assign a49794 = a49792 & ~l890;
assign a49796 = ~a49794 & ~a49790;
assign a49798 = a49796 & ~a41644;
assign a49800 = ~a44466 & ~a43952;
assign a49804 = a49802 & a48912;
assign a49806 = ~a49804 & a49788;
assign a49808 = ~l2390 & l890;
assign a49810 = a49768 & ~a40726;
assign a49812 = ~a49810 & a41020;
assign a49814 = ~a49812 & i670;
assign a49816 = a49814 & ~l890;
assign a49818 = ~a49816 & ~a49808;
assign a49820 = a49818 & ~a41644;
assign a49822 = ~a44456 & ~a44142;
assign a49826 = a49824 & a48862;
assign a49828 = ~a49826 & a49806;
assign a49830 = ~a44444 & ~a44098;
assign a49832 = ~l2396 & l890;
assign a49834 = ~a41020 & i670;
assign a49836 = ~a49834 & ~i648;
assign a49838 = ~a49836 & ~l890;
assign a49840 = ~a49838 & ~a49832;
assign a49844 = a49842 & a48924;
assign a49846 = ~a49844 & a49828;
assign a49848 = ~a44436 & ~a43902;
assign a49850 = ~l2400 & l890;
assign a49852 = ~a41020 & ~a40726;
assign a49854 = a49852 & i670;
assign a49856 = ~a49854 & ~i648;
assign a49858 = ~a49856 & ~l890;
assign a49860 = ~a49858 & ~a49850;
assign a49864 = a49862 & a48876;
assign a49866 = ~a49864 & a49846;
assign a49868 = ~a44422 & ~a43840;
assign a49870 = ~l2404 & l890;
assign a49872 = a45216 & a44964;
assign a49874 = ~a49872 & ~i648;
assign a49876 = ~a49874 & ~l890;
assign a49878 = ~a49876 & ~a49870;
assign a49882 = a49880 & a48884;
assign a49884 = ~a49882 & a49866;
assign a49886 = ~a49884 & ~a45586;
assign a49888 = a49740 & a49714;
assign a49890 = a49718 & a44834;
assign a49892 = ~a49890 & ~a49888;
assign a49894 = a49758 & a48898;
assign a49896 = ~a49894 & a49892;
assign a49898 = a49784 & a48838;
assign a49900 = ~a49898 & a49896;
assign a49902 = a49802 & a48846;
assign a49904 = ~a49902 & a49900;
assign a49906 = a49824 & a48912;
assign a49908 = ~a49906 & a49904;
assign a49910 = a49842 & a48862;
assign a49912 = ~a49910 & a49908;
assign a49914 = a49862 & a48924;
assign a49916 = ~a49914 & a49912;
assign a49918 = a49880 & a48876;
assign a49920 = ~a49918 & a49916;
assign a49922 = a48884 & a48728;
assign a49924 = ~a49922 & a49920;
assign a49926 = ~a49924 & a45586;
assign a49928 = ~a49926 & ~a49886;
assign a49930 = ~a49928 & ~a49712;
assign a49934 = ~a41788 & a41644;
assign a49936 = a45612 & l2370;
assign a49938 = ~a48858 & ~a48838;
assign a49940 = a49938 & ~a48844;
assign a49942 = ~a49940 & a45616;
assign a49944 = ~a49942 & ~a49936;
assign a49946 = a49944 & ~a49934;
assign a49948 = ~a41834 & a41644;
assign a49950 = a45612 & l2372;
assign a49952 = ~a48922 & ~a48876;
assign a49954 = ~a49952 & a45616;
assign a49956 = ~a49954 & ~a49950;
assign a49958 = a49956 & ~a49948;
assign a49960 = ~a44942 & a44888;
assign a49962 = a48750 & a44844;
assign a49964 = a49962 & a44870;
assign a49966 = ~a49964 & ~a44920;
assign a49968 = a49966 & ~a44902;
assign a49970 = a49968 & a49960;
assign a49972 = a44930 & a44870;
assign a49974 = a44946 & ~a41660;
assign a49976 = a48758 & ~a41678;
assign a49978 = a44924 & ~a41660;
assign a49980 = ~a49978 & ~a49976;
assign a49982 = a49980 & ~a49974;
assign a49984 = a49982 & ~a49972;
assign a49986 = a49984 & a44940;
assign a49988 = a49986 & a49970;
assign a49990 = ~a49988 & i674;
assign a49992 = a48838 & a45586;
assign a49994 = ~a49992 & ~a49990;
assign a49998 = a45586 & a45232;
assign a50000 = a49998 & a48844;
assign a50002 = a44856 & ~a41660;
assign a50004 = a50002 & a44904;
assign a50006 = ~a50004 & ~a44908;
assign a50008 = a50006 & a49960;
assign a50010 = a44936 & a41742;
assign a50012 = a50010 & a44844;
assign a50014 = ~a50012 & a49968;
assign a50016 = a50014 & ~a44930;
assign a50018 = a50016 & a50008;
assign a50020 = ~a50018 & i674;
assign a50022 = ~a50020 & ~i650;
assign a50026 = a48844 & a48784;
assign a50028 = a50014 & ~a44942;
assign a50030 = a50028 & a50006;
assign a50032 = a44930 & ~a41678;
assign a50034 = ~a50032 & ~a44884;
assign a50036 = a50034 & a50030;
assign a50038 = a44930 & ~a41660;
assign a50040 = a44922 & a44854;
assign a50042 = a50040 & a44870;
assign a50044 = a48740 & ~a41742;
assign a50046 = a48756 & a41678;
assign a50048 = a50046 & ~a41742;
assign a50050 = a50002 & ~a41742;
assign a50052 = ~a50050 & ~a50048;
assign a50054 = a50052 & ~a50044;
assign a50056 = a50054 & ~a50042;
assign a50058 = a50056 & ~a50038;
assign a50060 = a50058 & a50036;
assign a50062 = ~a50060 & i674;
assign a50064 = ~a50062 & ~i650;
assign a50068 = a44944 & ~a41742;
assign a50070 = ~a50040 & ~a44880;
assign a50072 = a50070 & ~a50068;
assign a50074 = a50072 & a50036;
assign a50076 = ~a50074 & i674;
assign a50078 = a45588 & l2370;
assign a50080 = a50078 & ~l2372;
assign a50082 = a50080 & a45232;
assign a50086 = a44922 & a44870;
assign a50088 = a50068 & ~a41660;
assign a50090 = a50032 & ~a41660;
assign a50092 = ~a44844 & ~a41660;
assign a50094 = a50092 & a48738;
assign a50096 = a44870 & a44858;
assign a50098 = ~a50096 & ~a50094;
assign a50100 = a50098 & ~a50090;
assign a50102 = a50100 & ~a50088;
assign a50104 = a50102 & ~a50086;
assign a50106 = a50104 & a50070;
assign a50108 = a50106 & a50030;
assign a50110 = ~a50108 & i674;
assign a50112 = a50080 & ~a45232;
assign a50116 = a48876 & a45586;
assign a50118 = ~a44854 & ~a41806;
assign a50120 = ~a50012 & ~a48754;
assign a50122 = a50120 & ~a50040;
assign a50124 = a50122 & ~a44908;
assign a50126 = a50124 & ~a48746;
assign a50128 = a50126 & ~a50118;
assign a50130 = a50128 & a49970;
assign a50132 = ~a50130 & i674;
assign a50134 = ~a50132 & ~i650;
assign a50138 = a48786 & l2372;
assign a50140 = a50010 & a41806;
assign a50142 = ~a50140 & ~a48752;
assign a50144 = a50142 & ~a48746;
assign a50146 = a50092 & a41742;
assign a50148 = a48756 & ~a41806;
assign a50150 = a48734 & a44870;
assign a50152 = ~a50150 & ~a50148;
assign a50154 = a50152 & ~a50146;
assign a50156 = a50154 & a50144;
assign a50158 = a50156 & a50008;
assign a50160 = ~a50158 & i674;
assign a50162 = ~a50160 & ~i650;
assign a50166 = a50144 & ~a48734;
assign a50168 = a50166 & a44912;
assign a50170 = ~a50168 & i674;
assign a50172 = a49998 & a48816;
assign a50174 = ~a50172 & ~i650;
assign a50178 = l2418 & i864;
assign a50180 = l2422 & ~i864;
assign a50182 = ~a50180 & ~a50178;
assign a50184 = l2406 & i864;
assign a50186 = l2424 & ~i864;
assign a50188 = ~a50186 & ~a50184;
assign a50190 = l2414 & i864;
assign a50192 = l2426 & ~i864;
assign a50194 = ~a50192 & ~a50190;
assign a50196 = l2410 & i864;
assign a50198 = l2428 & ~i864;
assign a50200 = ~a50198 & ~a50196;
assign a50202 = ~a33512 & l2430;
assign a50204 = a35382 & ~a35314;
assign a50206 = ~a35382 & a35314;
assign a50208 = ~a50206 & ~a50204;
assign a50210 = a50208 & ~a35248;
assign a50212 = ~a50208 & a35248;
assign a50214 = ~a50212 & ~a50210;
assign a50216 = a50214 & ~a35182;
assign a50218 = ~a50214 & a35182;
assign a50220 = ~a50218 & ~a50216;
assign a50222 = a50220 & ~a35116;
assign a50224 = ~a50220 & a35116;
assign a50226 = ~a50224 & ~a50222;
assign a50228 = a50226 & ~a35050;
assign a50230 = ~a50226 & a35050;
assign a50232 = ~a50230 & ~a50228;
assign a50234 = a50232 & ~a34984;
assign a50236 = ~a50232 & a34984;
assign a50238 = ~a50236 & ~a50234;
assign a50240 = a50238 & ~a31036;
assign a50242 = ~a50238 & a31036;
assign a50244 = ~a50242 & ~a50240;
assign a50246 = ~a50244 & a33512;
assign a50248 = ~a50246 & ~a50202;
assign a50250 = ~a34964 & l2432;
assign a50252 = ~a50244 & a34964;
assign a50254 = ~a50252 & ~a50250;
assign a50256 = ~a34956 & l2434;
assign a50258 = ~a50244 & a34956;
assign a50260 = ~a50258 & ~a50256;
assign a50262 = ~a34948 & l2436;
assign a50264 = ~a50244 & a34948;
assign a50266 = ~a50264 & ~a50262;
assign a50268 = ~a34940 & l2438;
assign a50270 = ~a50244 & a34940;
assign a50272 = ~a50270 & ~a50268;
assign a50274 = ~a34930 & l2440;
assign a50276 = ~a50244 & a34930;
assign a50278 = ~a50276 & ~a50274;
assign a50280 = ~a34922 & l2442;
assign a50282 = ~a50244 & a34922;
assign a50284 = ~a50282 & ~a50280;
assign a50286 = ~l2444 & l890;
assign a50288 = i866 & ~i14;
assign a50290 = i868 & ~i14;
assign a50292 = ~a50290 & ~a11208;
assign a50294 = ~a50292 & ~a50288;
assign a50296 = a50292 & a50288;
assign a50298 = ~a50296 & ~a50294;
assign a50300 = a50298 & ~a4826;
assign a50302 = ~a50298 & a4826;
assign a50304 = ~a50302 & ~a50300;
assign a50306 = a50304 & ~a4684;
assign a50308 = ~a50304 & a4684;
assign a50310 = ~a50308 & ~a50306;
assign a50312 = a50310 & ~a4524;
assign a50314 = ~a50310 & a4524;
assign a50316 = ~a50314 & ~a50312;
assign a50318 = a50316 & ~a4364;
assign a50320 = ~a50316 & a4364;
assign a50322 = ~a50320 & ~a50318;
assign a50324 = a50322 & ~a4218;
assign a50326 = ~a50322 & a4218;
assign a50328 = ~a50326 & ~a50324;
assign a50330 = a50328 & ~a4104;
assign a50332 = ~a50328 & a4104;
assign a50334 = ~a50332 & ~a50330;
assign a50336 = ~a50334 & a2722;
assign a50338 = a50336 & ~l890;
assign a50340 = ~a50338 & ~a50286;
assign a50342 = ~a50340 & ~a31028;
assign a50344 = ~a50244 & a31028;
assign a50348 = ~l2446 & l890;
assign a50350 = i870 & ~i12;
assign a50352 = ~a50350 & a2658;
assign a50354 = i872 & ~i12;
assign a50356 = ~a50354 & ~a4528;
assign a50358 = i874 & ~i12;
assign a50360 = ~a50358 & ~a4688;
assign a50362 = i876 & ~i12;
assign a50364 = ~a50362 & ~i12;
assign a50366 = i878 & ~i12;
assign a50368 = ~a50366 & ~a4830;
assign a50370 = ~a50368 & ~a50364;
assign a50372 = a50368 & a50364;
assign a50374 = ~a50372 & ~a50370;
assign a50376 = a50374 & ~a50360;
assign a50378 = ~a50374 & a50360;
assign a50380 = ~a50378 & ~a50376;
assign a50382 = a50380 & ~a50356;
assign a50384 = ~a50380 & a50356;
assign a50386 = ~a50384 & ~a50382;
assign a50388 = a50386 & a2568;
assign a50390 = ~a50386 & ~a2568;
assign a50392 = ~a50390 & ~a50388;
assign a50394 = a50392 & a2662;
assign a50396 = ~a50392 & ~a2662;
assign a50398 = ~a50396 & ~a50394;
assign a50400 = a50398 & a50352;
assign a50402 = ~a50398 & ~a50352;
assign a50404 = ~a50402 & ~a50400;
assign a50406 = ~a50404 & ~a2700;
assign a50408 = ~a50334 & a4086;
assign a50410 = ~a50408 & ~a50406;
assign a50412 = ~a50410 & ~l890;
assign a50414 = ~a50412 & ~a50348;
assign a50416 = ~a50414 & ~a19884;
assign a50418 = ~a50244 & a19884;
assign a50422 = ~a34914 & l2448;
assign a50424 = ~a50244 & a34914;
assign a50426 = ~a50424 & ~a50422;
assign a50428 = ~l2450 & l890;
assign a50430 = ~i642 & i638;
assign a50432 = i642 & ~i638;
assign a50434 = ~a50432 & ~a50430;
assign a50436 = a50434 & i634;
assign a50438 = ~a50434 & ~i634;
assign a50440 = ~a50438 & ~a50436;
assign a50442 = a50440 & i592;
assign a50444 = ~a50440 & ~i592;
assign a50446 = ~a50444 & ~a50442;
assign a50448 = a50446 & i598;
assign a50450 = ~a50446 & ~i598;
assign a50452 = ~a50450 & ~a50448;
assign a50454 = a50452 & i602;
assign a50456 = ~a50452 & ~i602;
assign a50458 = ~a50456 & ~a50454;
assign a50460 = a50458 & i604;
assign a50462 = ~a50458 & ~i604;
assign a50464 = ~a50462 & ~a50460;
assign a50466 = a50464 & a38260;
assign a50468 = ~a50464 & ~a38260;
assign a50470 = ~a50468 & ~a50466;
assign a50472 = ~a50470 & a41902;
assign a50474 = a50472 & ~a41896;
assign a50476 = i714 & ~i710;
assign a50478 = ~i714 & i710;
assign a50480 = ~a50478 & ~a50476;
assign a50482 = a50480 & i718;
assign a50484 = ~a50480 & ~i718;
assign a50486 = ~a50484 & ~a50482;
assign a50488 = a50486 & i722;
assign a50490 = ~a50486 & ~i722;
assign a50492 = ~a50490 & ~a50488;
assign a50494 = a50492 & i726;
assign a50496 = ~a50492 & ~i726;
assign a50498 = ~a50496 & ~a50494;
assign a50500 = a50498 & i730;
assign a50502 = ~a50498 & ~i730;
assign a50504 = ~a50502 & ~a50500;
assign a50506 = a50504 & i734;
assign a50508 = ~a50504 & ~i734;
assign a50510 = ~a50508 & ~a50506;
assign a50512 = a50510 & i738;
assign a50514 = ~a50510 & ~i738;
assign a50516 = ~a50514 & ~a50512;
assign a50518 = ~a50516 & a41896;
assign a50520 = ~a50518 & ~a50474;
assign a50522 = ~a50520 & ~a41916;
assign a50524 = ~i826 & i822;
assign a50526 = i826 & ~i822;
assign a50528 = ~a50526 & ~a50524;
assign a50530 = a50528 & i772;
assign a50532 = ~a50528 & ~i772;
assign a50534 = ~a50532 & ~a50530;
assign a50536 = a50534 & i766;
assign a50538 = ~a50534 & ~i766;
assign a50540 = ~a50538 & ~a50536;
assign a50542 = a50540 & i760;
assign a50544 = ~a50540 & ~i760;
assign a50546 = ~a50544 & ~a50542;
assign a50548 = a50546 & i754;
assign a50550 = ~a50546 & ~i754;
assign a50552 = ~a50550 & ~a50548;
assign a50554 = a50552 & i748;
assign a50556 = ~a50552 & ~i748;
assign a50558 = ~a50556 & ~a50554;
assign a50560 = a50558 & i742;
assign a50562 = ~a50558 & ~i742;
assign a50564 = ~a50562 & ~a50560;
assign a50566 = ~a50564 & a41916;
assign a50568 = ~a50566 & ~a50522;
assign a50570 = ~a50568 & ~l890;
assign a50572 = ~a50570 & ~a50428;
assign a50574 = ~a50572 & ~a44436;
assign a50576 = ~i828 & i824;
assign a50578 = i828 & ~i824;
assign a50580 = ~a50578 & ~a50576;
assign a50582 = a50580 & i774;
assign a50584 = ~a50580 & ~i774;
assign a50586 = ~a50584 & ~a50582;
assign a50588 = a50586 & i768;
assign a50590 = ~a50586 & ~i768;
assign a50592 = ~a50590 & ~a50588;
assign a50594 = a50592 & i762;
assign a50596 = ~a50592 & ~i762;
assign a50598 = ~a50596 & ~a50594;
assign a50600 = a50598 & i756;
assign a50602 = ~a50598 & ~i756;
assign a50604 = ~a50602 & ~a50600;
assign a50606 = a50604 & i750;
assign a50608 = ~a50604 & ~i750;
assign a50610 = ~a50608 & ~a50606;
assign a50612 = a50610 & i744;
assign a50614 = ~a50610 & ~i744;
assign a50616 = ~a50614 & ~a50612;
assign a50618 = ~a50616 & a44436;
assign a50622 = ~l2452 & l890;
assign a50624 = ~a50470 & a41936;
assign a50626 = a50624 & ~a41940;
assign a50628 = ~a50516 & a41940;
assign a50630 = ~a50628 & ~a50626;
assign a50632 = ~a50630 & ~a41948;
assign a50634 = ~a50564 & a41948;
assign a50636 = ~a50634 & ~a50632;
assign a50638 = ~a50636 & ~l890;
assign a50640 = ~a50638 & ~a50622;
assign a50642 = ~a50640 & ~a44444;
assign a50644 = ~a50616 & a44444;
assign a50648 = ~l2454 & l890;
assign a50650 = ~a50470 & a41970;
assign a50652 = a50650 & ~a41974;
assign a50654 = ~a50516 & a41974;
assign a50656 = ~a50654 & ~a50652;
assign a50658 = ~a50656 & ~a41986;
assign a50660 = ~a50564 & a41986;
assign a50662 = ~a50660 & ~a50658;
assign a50664 = ~a50662 & ~l890;
assign a50666 = ~a50664 & ~a50648;
assign a50668 = ~a50666 & ~a44456;
assign a50670 = ~a50616 & a44456;
assign a50674 = ~l2456 & l890;
assign a50676 = ~a50470 & a42006;
assign a50678 = a50676 & ~a42010;
assign a50680 = ~a50516 & a42010;
assign a50682 = ~a50680 & ~a50678;
assign a50684 = ~a50682 & ~a42020;
assign a50686 = ~a50564 & a42020;
assign a50688 = ~a50686 & ~a50684;
assign a50690 = ~a50688 & ~l890;
assign a50692 = ~a50690 & ~a50674;
assign a50694 = ~a50692 & ~a44466;
assign a50696 = ~a50616 & a44466;
assign a50700 = ~l2458 & l890;
assign a50702 = ~a50470 & a42038;
assign a50704 = a50702 & ~a42042;
assign a50706 = ~a50516 & a42042;
assign a50708 = ~a50706 & ~a50704;
assign a50710 = ~a50708 & ~a42052;
assign a50712 = ~a50564 & a42052;
assign a50714 = ~a50712 & ~a50710;
assign a50716 = ~a50714 & ~l890;
assign a50718 = ~a50716 & ~a50700;
assign a50720 = ~a50718 & ~a44476;
assign a50722 = ~a50616 & a44476;
assign a50726 = ~l2460 & l890;
assign a50728 = ~a50470 & a42074;
assign a50730 = a50728 & ~a42078;
assign a50732 = ~a50516 & a42078;
assign a50734 = ~a50732 & ~a50730;
assign a50736 = ~a50734 & ~a42086;
assign a50738 = ~a50564 & a42086;
assign a50740 = ~a50738 & ~a50736;
assign a50742 = ~a50740 & ~l890;
assign a50744 = ~a50742 & ~a50726;
assign a50746 = ~a50744 & ~a44484;
assign a50748 = ~a50616 & a44484;
assign a50752 = ~l2462 & l890;
assign a50754 = ~a50470 & a41112;
assign a50756 = a50754 & ~a41108;
assign a50758 = ~a50516 & a41108;
assign a50760 = ~a50758 & ~a50756;
assign a50762 = ~a50760 & ~a42106;
assign a50764 = ~a50564 & a42106;
assign a50766 = ~a50764 & ~a50762;
assign a50768 = ~a50766 & ~l890;
assign a50770 = ~a50768 & ~a50752;
assign a50772 = ~a50770 & ~a44492;
assign a50774 = ~a50616 & a44492;
assign a50778 = ~l2464 & l890;
assign a50780 = ~a50470 & a40444;
assign a50782 = a50780 & ~a41064;
assign a50784 = ~a50516 & a41064;
assign a50786 = ~a50784 & ~a50782;
assign a50788 = ~a50786 & ~a42128;
assign a50790 = ~a50564 & a42128;
assign a50792 = ~a50790 & ~a50788;
assign a50794 = ~a50792 & ~l890;
assign a50796 = ~a50794 & ~a50778;
assign a50798 = ~a50796 & ~a44500;
assign a50800 = ~a50616 & a44500;
assign a50804 = ~l2466 & l890;
assign a50806 = ~a50470 & a40454;
assign a50808 = a50806 & ~a41086;
assign a50810 = ~a50516 & a41086;
assign a50812 = ~a50810 & ~a50808;
assign a50814 = ~a50812 & ~a42148;
assign a50816 = ~a50564 & a42148;
assign a50818 = ~a50816 & ~a50814;
assign a50820 = ~a50818 & ~l890;
assign a50822 = ~a50820 & ~a50804;
assign a50824 = ~a50822 & ~a44508;
assign a50826 = ~a50616 & a44508;
assign a50830 = ~l2468 & l890;
assign a50832 = ~a50470 & a41546;
assign a50834 = a50832 & ~a41852;
assign a50836 = ~a50516 & a41852;
assign a50838 = ~a50836 & ~a50834;
assign a50840 = ~a50838 & ~a41868;
assign a50842 = ~a50564 & a41868;
assign a50844 = ~a50842 & ~a50840;
assign a50846 = ~a50844 & ~l890;
assign a50848 = ~a50846 & ~a50830;
assign a50850 = ~a50848 & ~a44422;
assign a50852 = ~a50616 & a44422;
assign a50856 = a15496 & a15330;
assign a50858 = a15164 & a14994;
assign a50860 = a14826 & a14656;
assign a50862 = a50860 & a50858;
assign a50864 = a50862 & a50856;
assign a50866 = a50864 & ~a15662;
assign a50868 = a50866 & a16170;
assign a50870 = a50860 & ~a14994;
assign a50872 = a50870 & a16178;
assign a50874 = ~a50872 & ~a50868;
assign a50876 = a50864 & a15662;
assign a50878 = a50876 & ~a15832;
assign a50880 = a50878 & a16168;
assign a50882 = a50876 & ~a16000;
assign a50884 = a50882 & a15832;
assign a50886 = a50884 & a16166;
assign a50888 = ~a50886 & ~a50880;
assign a50890 = a50860 & a14994;
assign a50892 = a50890 & ~a15164;
assign a50894 = a50892 & a16176;
assign a50896 = a50862 & ~a15330;
assign a50898 = a50896 & a16174;
assign a50900 = a15330 & a15164;
assign a50902 = a50890 & ~a15496;
assign a50904 = a50902 & a16172;
assign a50906 = a50904 & a50900;
assign a50908 = ~a50906 & ~a50898;
assign a50910 = a50908 & ~a50868;
assign a50912 = a50910 & ~a50894;
assign a50914 = a16000 & a15832;
assign a50916 = a50914 & a15662;
assign a50918 = a50916 & a50856;
assign a50920 = a50918 & a15164;
assign a50922 = a50920 & a14994;
assign a50924 = a50922 & a14826;
assign a50926 = a50924 & ~a16166;
assign a50928 = a50926 & a14656;
assign a50930 = a16182 & ~a14656;
assign a50932 = a16180 & ~a14826;
assign a50934 = a50932 & a14656;
assign a50936 = ~a50934 & ~a50872;
assign a50938 = a50936 & ~a50930;
assign a50940 = a50938 & ~a50928;
assign a50942 = a50940 & a50912;
assign a50944 = a50942 & a50888;
assign a50946 = a50944 & l2470;
assign a50948 = ~a50930 & ~a50898;
assign a50950 = a50948 & ~a50886;
assign a50952 = a50950 & ~a50946;
assign a50954 = a50952 & a50874;
assign a50956 = a50944 & l2472;
assign a50958 = ~a50956 & a50888;
assign a50960 = a50944 & l2474;
assign a50962 = ~a50960 & a50912;
assign a50964 = a50944 & l2476;
assign a50966 = ~a50934 & ~a50906;
assign a50968 = a50966 & ~a50964;
assign a50970 = a50968 & a50874;
assign a50974 = ~l2484 & l2482;
assign a50976 = l2484 & l2482;
assign a50978 = a50976 & ~l2486;
assign a50980 = l2484 & ~l2482;
assign a50982 = ~a50980 & ~a50978;
assign a50984 = a50982 & ~a50974;
assign a50988 = ~a50978 & l2484;
assign a50992 = ~a50976 & ~l2486;
assign a50994 = ~a50992 & ~a50976;
assign a50996 = ~a50994 & ~l924;
assign a50998 = ~l2488 & ~l1186;
assign a51002 = ~a19394 & a18838;
assign a51004 = a19394 & ~a18838;
assign a51006 = ~a51004 & ~a51002;
assign a51008 = a51006 & ~a19318;
assign a51010 = ~a51006 & a19318;
assign a51012 = ~a51010 & ~a51008;
assign a51014 = a51012 & ~a19236;
assign a51016 = ~a51012 & a19236;
assign a51018 = ~a51016 & ~a51014;
assign a51020 = a51018 & ~a19154;
assign a51022 = ~a51018 & a19154;
assign a51024 = ~a51022 & ~a51020;
assign a51026 = a51024 & ~a19072;
assign a51028 = ~a51024 & a19072;
assign a51030 = ~a51028 & ~a51026;
assign a51032 = a51030 & ~a18990;
assign a51034 = ~a51030 & a18990;
assign a51036 = ~a51034 & ~a51032;
assign a51038 = a51036 & ~a18916;
assign a51040 = ~a51036 & a18916;
assign a51042 = ~a51040 & ~a51038;
assign a51044 = a18834 & l2430;
assign a51046 = a18650 & l2432;
assign a51048 = a18638 & l2434;
assign a51050 = a51048 & l880;
assign a51052 = l2436 & ~l880;
assign a51054 = a51052 & a18638;
assign a51056 = a2530 & l2438;
assign a51058 = a51056 & l880;
assign a51060 = a18618 & l2440;
assign a51062 = a2526 & ~l1006;
assign a51064 = a51062 & l2442;
assign a51066 = a18608 & ~l880;
assign a51068 = a51066 & ~a50340;
assign a51070 = a18670 & a18598;
assign a51072 = a51070 & ~a50414;
assign a51074 = a18586 & ~l1002;
assign a51076 = a51074 & l2448;
assign a51078 = ~a51076 & ~a51072;
assign a51080 = a51078 & ~a51068;
assign a51082 = a51080 & ~a51064;
assign a51084 = a51082 & ~a51060;
assign a51086 = a51084 & ~a51058;
assign a51088 = a51086 & ~a51054;
assign a51090 = a51088 & ~a51050;
assign a51092 = a51090 & ~a51046;
assign a51094 = a51092 & ~a51044;
assign a51096 = a51094 & ~a51042;
assign a51098 = ~a51094 & a51042;
assign a51100 = ~a51098 & ~a51096;
assign p0 = ~a51100;

assert property (~p0);

endmodule
